// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire clknet_leaf_0_i_clk;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net74;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net75;
 wire net90;
 wire net91;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net108;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdx[5] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_mapdy[5] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.texu[5] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.spi_registers.got_new_floor ;
 wire \rbzero.spi_registers.got_new_leak ;
 wire \rbzero.spi_registers.got_new_mapd ;
 wire \rbzero.spi_registers.got_new_other ;
 wire \rbzero.spi_registers.got_new_sky ;
 wire \rbzero.spi_registers.got_new_vinf ;
 wire \rbzero.spi_registers.got_new_vshift ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.new_floor[0] ;
 wire \rbzero.spi_registers.new_floor[1] ;
 wire \rbzero.spi_registers.new_floor[2] ;
 wire \rbzero.spi_registers.new_floor[3] ;
 wire \rbzero.spi_registers.new_floor[4] ;
 wire \rbzero.spi_registers.new_floor[5] ;
 wire \rbzero.spi_registers.new_leak[0] ;
 wire \rbzero.spi_registers.new_leak[1] ;
 wire \rbzero.spi_registers.new_leak[2] ;
 wire \rbzero.spi_registers.new_leak[3] ;
 wire \rbzero.spi_registers.new_leak[4] ;
 wire \rbzero.spi_registers.new_leak[5] ;
 wire \rbzero.spi_registers.new_mapd[0] ;
 wire \rbzero.spi_registers.new_mapd[10] ;
 wire \rbzero.spi_registers.new_mapd[11] ;
 wire \rbzero.spi_registers.new_mapd[12] ;
 wire \rbzero.spi_registers.new_mapd[13] ;
 wire \rbzero.spi_registers.new_mapd[14] ;
 wire \rbzero.spi_registers.new_mapd[15] ;
 wire \rbzero.spi_registers.new_mapd[1] ;
 wire \rbzero.spi_registers.new_mapd[2] ;
 wire \rbzero.spi_registers.new_mapd[3] ;
 wire \rbzero.spi_registers.new_mapd[4] ;
 wire \rbzero.spi_registers.new_mapd[5] ;
 wire \rbzero.spi_registers.new_mapd[6] ;
 wire \rbzero.spi_registers.new_mapd[7] ;
 wire \rbzero.spi_registers.new_mapd[8] ;
 wire \rbzero.spi_registers.new_mapd[9] ;
 wire \rbzero.spi_registers.new_other[0] ;
 wire \rbzero.spi_registers.new_other[10] ;
 wire \rbzero.spi_registers.new_other[1] ;
 wire \rbzero.spi_registers.new_other[2] ;
 wire \rbzero.spi_registers.new_other[3] ;
 wire \rbzero.spi_registers.new_other[4] ;
 wire \rbzero.spi_registers.new_other[6] ;
 wire \rbzero.spi_registers.new_other[7] ;
 wire \rbzero.spi_registers.new_other[8] ;
 wire \rbzero.spi_registers.new_other[9] ;
 wire \rbzero.spi_registers.new_sky[0] ;
 wire \rbzero.spi_registers.new_sky[1] ;
 wire \rbzero.spi_registers.new_sky[2] ;
 wire \rbzero.spi_registers.new_sky[3] ;
 wire \rbzero.spi_registers.new_sky[4] ;
 wire \rbzero.spi_registers.new_sky[5] ;
 wire \rbzero.spi_registers.new_vinf ;
 wire \rbzero.spi_registers.new_vshift[0] ;
 wire \rbzero.spi_registers.new_vshift[1] ;
 wire \rbzero.spi_registers.new_vshift[2] ;
 wire \rbzero.spi_registers.new_vshift[3] ;
 wire \rbzero.spi_registers.new_vshift[4] ;
 wire \rbzero.spi_registers.new_vshift[5] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.side ;
 wire \rbzero.wall_tracer.state[0] ;
 wire \rbzero.wall_tracer.state[10] ;
 wire \rbzero.wall_tracer.state[11] ;
 wire \rbzero.wall_tracer.state[12] ;
 wire \rbzero.wall_tracer.state[13] ;
 wire \rbzero.wall_tracer.state[14] ;
 wire \rbzero.wall_tracer.state[1] ;
 wire \rbzero.wall_tracer.state[2] ;
 wire \rbzero.wall_tracer.state[3] ;
 wire \rbzero.wall_tracer.state[4] ;
 wire \rbzero.wall_tracer.state[5] ;
 wire \rbzero.wall_tracer.state[6] ;
 wire \rbzero.wall_tracer.state[7] ;
 wire \rbzero.wall_tracer.state[8] ;
 wire \rbzero.wall_tracer.state[9] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.texu[0] ;
 wire \rbzero.wall_tracer.texu[1] ;
 wire \rbzero.wall_tracer.texu[2] ;
 wire \rbzero.wall_tracer.texu[3] ;
 wire \rbzero.wall_tracer.texu[4] ;
 wire \rbzero.wall_tracer.texu[5] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \rbzero.wall_tracer.wall[0] ;
 wire \rbzero.wall_tracer.wall[1] ;
 wire net92;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net125;
 wire net72;
 wire net73;
 wire net124;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_0__04486_;
 wire clknet_1_0__leaf__04486_;
 wire clknet_1_1__leaf__04486_;
 wire clknet_0__02755_;
 wire clknet_1_0__leaf__02755_;
 wire clknet_1_1__leaf__02755_;
 wire clknet_0__02754_;
 wire clknet_1_0__leaf__02754_;
 wire clknet_1_1__leaf__02754_;
 wire clknet_0__02743_;
 wire clknet_1_0__leaf__02743_;
 wire clknet_1_1__leaf__02743_;
 wire clknet_0__02753_;
 wire clknet_1_0__leaf__02753_;
 wire clknet_1_1__leaf__02753_;
 wire clknet_0__02752_;
 wire clknet_1_0__leaf__02752_;
 wire clknet_1_1__leaf__02752_;
 wire clknet_0__02751_;
 wire clknet_1_0__leaf__02751_;
 wire clknet_1_1__leaf__02751_;
 wire clknet_0__02750_;
 wire clknet_1_0__leaf__02750_;
 wire clknet_1_1__leaf__02750_;
 wire clknet_0__02749_;
 wire clknet_1_0__leaf__02749_;
 wire clknet_1_1__leaf__02749_;
 wire clknet_0__02748_;
 wire clknet_1_0__leaf__02748_;
 wire clknet_1_1__leaf__02748_;
 wire clknet_0__02747_;
 wire clknet_1_0__leaf__02747_;
 wire clknet_1_1__leaf__02747_;
 wire clknet_0__02746_;
 wire clknet_1_0__leaf__02746_;
 wire clknet_1_1__leaf__02746_;
 wire clknet_0__02745_;
 wire clknet_1_0__leaf__02745_;
 wire clknet_1_1__leaf__02745_;
 wire clknet_0__02744_;
 wire clknet_1_0__leaf__02744_;
 wire clknet_1_1__leaf__02744_;
 wire clknet_0__02732_;
 wire clknet_1_0__leaf__02732_;
 wire clknet_1_1__leaf__02732_;
 wire clknet_0__02742_;
 wire clknet_1_0__leaf__02742_;
 wire clknet_1_1__leaf__02742_;
 wire clknet_0__02741_;
 wire clknet_1_0__leaf__02741_;
 wire clknet_1_1__leaf__02741_;
 wire clknet_0__02740_;
 wire clknet_1_0__leaf__02740_;
 wire clknet_1_1__leaf__02740_;
 wire clknet_0__02739_;
 wire clknet_1_0__leaf__02739_;
 wire clknet_1_1__leaf__02739_;
 wire clknet_0__02738_;
 wire clknet_1_0__leaf__02738_;
 wire clknet_1_1__leaf__02738_;
 wire clknet_0__02737_;
 wire clknet_1_0__leaf__02737_;
 wire clknet_1_1__leaf__02737_;
 wire clknet_0__02736_;
 wire clknet_1_0__leaf__02736_;
 wire clknet_1_1__leaf__02736_;
 wire clknet_0__02735_;
 wire clknet_1_0__leaf__02735_;
 wire clknet_1_1__leaf__02735_;
 wire clknet_0__02734_;
 wire clknet_1_0__leaf__02734_;
 wire clknet_1_1__leaf__02734_;
 wire clknet_0__02733_;
 wire clknet_1_0__leaf__02733_;
 wire clknet_1_1__leaf__02733_;
 wire clknet_0__02440_;
 wire clknet_1_0__leaf__02440_;
 wire clknet_1_1__leaf__02440_;
 wire clknet_0__02731_;
 wire clknet_1_0__leaf__02731_;
 wire clknet_1_1__leaf__02731_;
 wire clknet_0__02730_;
 wire clknet_1_0__leaf__02730_;
 wire clknet_1_1__leaf__02730_;
 wire clknet_0__02729_;
 wire clknet_1_0__leaf__02729_;
 wire clknet_1_1__leaf__02729_;
 wire clknet_0__02728_;
 wire clknet_1_0__leaf__02728_;
 wire clknet_1_1__leaf__02728_;
 wire clknet_0__02727_;
 wire clknet_1_0__leaf__02727_;
 wire clknet_1_1__leaf__02727_;
 wire clknet_0__02726_;
 wire clknet_1_0__leaf__02726_;
 wire clknet_1_1__leaf__02726_;
 wire clknet_0__02725_;
 wire clknet_1_0__leaf__02725_;
 wire clknet_1_1__leaf__02725_;
 wire clknet_0__02724_;
 wire clknet_1_0__leaf__02724_;
 wire clknet_1_1__leaf__02724_;
 wire clknet_0__02723_;
 wire clknet_1_0__leaf__02723_;
 wire clknet_1_1__leaf__02723_;
 wire clknet_0__02441_;
 wire clknet_1_0__leaf__02441_;
 wire clknet_1_1__leaf__02441_;
 wire clknet_0__02433_;
 wire clknet_1_0__leaf__02433_;
 wire clknet_1_1__leaf__02433_;
 wire clknet_0__02439_;
 wire clknet_1_0__leaf__02439_;
 wire clknet_1_1__leaf__02439_;
 wire clknet_0__02438_;
 wire clknet_1_0__leaf__02438_;
 wire clknet_1_1__leaf__02438_;
 wire clknet_0__02437_;
 wire clknet_1_0__leaf__02437_;
 wire clknet_1_1__leaf__02437_;
 wire clknet_0__02436_;
 wire clknet_1_0__leaf__02436_;
 wire clknet_1_1__leaf__02436_;
 wire clknet_0__02435_;
 wire clknet_1_0__leaf__02435_;
 wire clknet_1_1__leaf__02435_;
 wire clknet_0__02434_;
 wire clknet_1_0__leaf__02434_;
 wire clknet_1_1__leaf__02434_;
 wire net71;

 sky130_fd_sc_hd__buf_2 _09717_ (.A(\gpout0.hpos[0] ),
    .X(_02899_));
 sky130_fd_sc_hd__buf_4 _09718_ (.A(\gpout0.hpos[7] ),
    .X(_02900_));
 sky130_fd_sc_hd__clkbuf_4 _09719_ (.A(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__clkbuf_4 _09720_ (.A(\gpout0.hpos[8] ),
    .X(_02902_));
 sky130_fd_sc_hd__inv_2 _09721_ (.A(\gpout0.hpos[9] ),
    .Y(_02903_));
 sky130_fd_sc_hd__nor2_1 _09722_ (.A(_02902_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__and2_1 _09723_ (.A(_02901_),
    .B(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__xor2_4 _09724_ (.A(net46),
    .B(net45),
    .X(_02906_));
 sky130_fd_sc_hd__buf_6 _09725_ (.A(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__and3_2 _09726_ (.A(_02899_),
    .B(_02905_),
    .C(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__buf_4 _09727_ (.A(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__clkbuf_4 _09728_ (.A(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _09729_ (.A0(\rbzero.tex_r1[63] ),
    .A1(net47),
    .S(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__clkbuf_1 _09730_ (.A(_02911_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _09731_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[63] ),
    .S(_02910_),
    .X(_02912_));
 sky130_fd_sc_hd__clkbuf_1 _09732_ (.A(_02912_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _09733_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_02910_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_1 _09734_ (.A(_02913_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _09735_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(_02910_),
    .X(_02914_));
 sky130_fd_sc_hd__clkbuf_1 _09736_ (.A(_02914_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _09737_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_02910_),
    .X(_02915_));
 sky130_fd_sc_hd__clkbuf_1 _09738_ (.A(_02915_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _09739_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_02910_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_1 _09740_ (.A(_02916_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _09741_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_02910_),
    .X(_02917_));
 sky130_fd_sc_hd__clkbuf_1 _09742_ (.A(_02917_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _09743_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(_02910_),
    .X(_02918_));
 sky130_fd_sc_hd__clkbuf_1 _09744_ (.A(_02918_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _09745_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_02910_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_1 _09746_ (.A(_02919_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(_02910_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _09748_ (.A(_02920_),
    .X(_01394_));
 sky130_fd_sc_hd__clkbuf_4 _09749_ (.A(_02909_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _09750_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__clkbuf_1 _09751_ (.A(_02922_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _09752_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(_02921_),
    .X(_02923_));
 sky130_fd_sc_hd__clkbuf_1 _09753_ (.A(_02923_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _09754_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_02921_),
    .X(_02924_));
 sky130_fd_sc_hd__clkbuf_1 _09755_ (.A(_02924_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _09756_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_02921_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_1 _09757_ (.A(_02925_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _09758_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_02921_),
    .X(_02926_));
 sky130_fd_sc_hd__clkbuf_1 _09759_ (.A(_02926_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _09760_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(_02921_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _09761_ (.A(_02927_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _09762_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_02921_),
    .X(_02928_));
 sky130_fd_sc_hd__clkbuf_1 _09763_ (.A(_02928_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(_02921_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_1 _09765_ (.A(_02929_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _09766_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_02921_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_1 _09767_ (.A(_02930_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _09768_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(_02921_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _09769_ (.A(_02931_),
    .X(_01384_));
 sky130_fd_sc_hd__clkbuf_4 _09770_ (.A(_02909_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _09771_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_1 _09772_ (.A(_02933_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _09773_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(_02932_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _09774_ (.A(_02934_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _09775_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_02932_),
    .X(_02935_));
 sky130_fd_sc_hd__clkbuf_1 _09776_ (.A(_02935_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _09777_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(_02932_),
    .X(_02936_));
 sky130_fd_sc_hd__clkbuf_1 _09778_ (.A(_02936_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _09779_ (.A0(\rbzero.tex_r1[39] ),
    .A1(net71),
    .S(_02932_),
    .X(_02937_));
 sky130_fd_sc_hd__clkbuf_1 _09780_ (.A(_02937_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _09781_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(_02932_),
    .X(_02938_));
 sky130_fd_sc_hd__clkbuf_1 _09782_ (.A(_02938_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _09783_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_02932_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_1 _09784_ (.A(_02939_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_02932_),
    .X(_02940_));
 sky130_fd_sc_hd__clkbuf_1 _09786_ (.A(_02940_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_02932_),
    .X(_02941_));
 sky130_fd_sc_hd__clkbuf_1 _09788_ (.A(_02941_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(_02932_),
    .X(_02942_));
 sky130_fd_sc_hd__clkbuf_1 _09790_ (.A(_02942_),
    .X(_01374_));
 sky130_fd_sc_hd__clkbuf_4 _09791_ (.A(_02909_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _09792_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _09793_ (.A(_02944_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _09794_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(_02943_),
    .X(_02945_));
 sky130_fd_sc_hd__clkbuf_1 _09795_ (.A(_02945_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _09796_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_02943_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _09797_ (.A(_02946_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _09798_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(_02943_),
    .X(_02947_));
 sky130_fd_sc_hd__clkbuf_1 _09799_ (.A(_02947_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _09800_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_02943_),
    .X(_02948_));
 sky130_fd_sc_hd__clkbuf_1 _09801_ (.A(_02948_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _09802_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(_02943_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _09803_ (.A(_02949_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_02943_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _09805_ (.A(_02950_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(_02943_),
    .X(_02951_));
 sky130_fd_sc_hd__clkbuf_1 _09807_ (.A(_02951_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _09808_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_02943_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_1 _09809_ (.A(_02952_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _09810_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(_02943_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _09811_ (.A(_02953_),
    .X(_01364_));
 sky130_fd_sc_hd__clkbuf_4 _09812_ (.A(_02909_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _09813_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__clkbuf_1 _09814_ (.A(_02955_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _09815_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(_02954_),
    .X(_02956_));
 sky130_fd_sc_hd__clkbuf_1 _09816_ (.A(_02956_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_02954_),
    .X(_02957_));
 sky130_fd_sc_hd__clkbuf_1 _09818_ (.A(_02957_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _09819_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(_02954_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_1 _09820_ (.A(_02958_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_02954_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_1 _09822_ (.A(_02959_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _09823_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(_02954_),
    .X(_02960_));
 sky130_fd_sc_hd__clkbuf_1 _09824_ (.A(_02960_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_02954_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_1 _09826_ (.A(_02961_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(_02954_),
    .X(_02962_));
 sky130_fd_sc_hd__clkbuf_1 _09828_ (.A(_02962_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _09829_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_02954_),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_1 _09830_ (.A(_02963_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _09831_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(_02954_),
    .X(_02964_));
 sky130_fd_sc_hd__clkbuf_1 _09832_ (.A(_02964_),
    .X(_01354_));
 sky130_fd_sc_hd__clkbuf_4 _09833_ (.A(_02909_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _09834_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__clkbuf_1 _09835_ (.A(_02966_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _09836_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_02965_),
    .X(_02967_));
 sky130_fd_sc_hd__clkbuf_1 _09837_ (.A(_02967_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _09838_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_02965_),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_1 _09839_ (.A(_02968_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _09840_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(_02965_),
    .X(_02969_));
 sky130_fd_sc_hd__clkbuf_1 _09841_ (.A(_02969_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _09842_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_02965_),
    .X(_02970_));
 sky130_fd_sc_hd__clkbuf_1 _09843_ (.A(_02970_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _09844_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_02965_),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_1 _09845_ (.A(_02971_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _09846_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_02965_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _09847_ (.A(_02972_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _09848_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(_02965_),
    .X(_02973_));
 sky130_fd_sc_hd__clkbuf_1 _09849_ (.A(_02973_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _09850_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_02965_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _09851_ (.A(_02974_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _09852_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(_02965_),
    .X(_02975_));
 sky130_fd_sc_hd__clkbuf_1 _09853_ (.A(_02975_),
    .X(_01344_));
 sky130_fd_sc_hd__clkbuf_4 _09854_ (.A(_02909_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _09855_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__clkbuf_1 _09856_ (.A(_02977_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _09857_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_02976_),
    .X(_02978_));
 sky130_fd_sc_hd__clkbuf_1 _09858_ (.A(_02978_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _09859_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_02976_),
    .X(_02979_));
 sky130_fd_sc_hd__clkbuf_1 _09860_ (.A(_02979_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _09861_ (.A0(\rbzero.tex_r1[0] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(_02976_),
    .X(_02980_));
 sky130_fd_sc_hd__clkbuf_1 _09862_ (.A(_02980_),
    .X(_01340_));
 sky130_fd_sc_hd__clkinv_8 _09863_ (.A(_02906_),
    .Y(_02981_));
 sky130_fd_sc_hd__or3b_2 _09864_ (.A(_02981_),
    .B(_02899_),
    .C_N(_02905_),
    .X(_02982_));
 sky130_fd_sc_hd__buf_4 _09865_ (.A(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__clkbuf_4 _09866_ (.A(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _09867_ (.A0(net47),
    .A1(\rbzero.tex_r0[63] ),
    .S(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__clkbuf_1 _09868_ (.A(_02985_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _09869_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_02984_),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_1 _09870_ (.A(_02986_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _09871_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_02984_),
    .X(_02987_));
 sky130_fd_sc_hd__clkbuf_1 _09872_ (.A(_02987_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _09873_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_02984_),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_1 _09874_ (.A(_02988_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _09875_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(_02984_),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_1 _09876_ (.A(_02989_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _09877_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_02984_),
    .X(_02990_));
 sky130_fd_sc_hd__clkbuf_1 _09878_ (.A(_02990_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(_02984_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _09880_ (.A(_02991_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _09881_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_02984_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _09882_ (.A(_02992_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(_02984_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_1 _09884_ (.A(_02993_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _09885_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_02984_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_1 _09886_ (.A(_02994_),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_4 _09887_ (.A(_02983_),
    .X(_02995_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_1 _09889_ (.A(_02996_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _09890_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_02995_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_1 _09891_ (.A(_02997_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _09892_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_02995_),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_1 _09893_ (.A(_02998_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_02995_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _09895_ (.A(_02999_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _09896_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(_02995_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_1 _09897_ (.A(_03000_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _09898_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_02995_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_1 _09899_ (.A(_03001_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _09900_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(_02995_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_1 _09901_ (.A(_03002_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _09902_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_02995_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_1 _09903_ (.A(_03003_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _09904_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_02995_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_1 _09905_ (.A(_03004_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _09906_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_02995_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_1 _09907_ (.A(_03005_),
    .X(_01320_));
 sky130_fd_sc_hd__clkbuf_4 _09908_ (.A(_02983_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _09909_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _09910_ (.A(_03007_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _09911_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_03006_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _09912_ (.A(_03008_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _09913_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(_03006_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _09914_ (.A(_03009_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _09915_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_03006_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_1 _09916_ (.A(_03010_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _09917_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(_03006_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_1 _09918_ (.A(_03011_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _09919_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_03006_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _09920_ (.A(_03012_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _09921_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(_03006_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _09922_ (.A(_03013_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _09923_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_03006_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_1 _09924_ (.A(_03014_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _09925_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(_03006_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_1 _09926_ (.A(_03015_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _09927_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_03006_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_1 _09928_ (.A(_03016_),
    .X(_01310_));
 sky130_fd_sc_hd__clkbuf_4 _09929_ (.A(_02983_),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _09930_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _09931_ (.A(_03018_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _09932_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_03017_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _09933_ (.A(_03019_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _09934_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(_03017_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_1 _09935_ (.A(_03020_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _09936_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_03017_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_1 _09937_ (.A(_03021_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _09938_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(_03017_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_1 _09939_ (.A(_03022_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _09940_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_03017_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_1 _09941_ (.A(_03023_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _09942_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_03017_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _09943_ (.A(_03024_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _09944_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_03017_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_1 _09945_ (.A(_03025_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _09946_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(_03017_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_1 _09947_ (.A(_03026_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _09948_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_03017_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_1 _09949_ (.A(_03027_),
    .X(_01300_));
 sky130_fd_sc_hd__clkbuf_4 _09950_ (.A(_02983_),
    .X(_03028_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _09952_ (.A(_03029_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_03028_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _09954_ (.A(_03030_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _09955_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(_03028_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _09956_ (.A(_03031_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_03028_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _09958_ (.A(_03032_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(_03028_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _09960_ (.A(_03033_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_03028_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _09962_ (.A(_03034_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(_03028_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _09964_ (.A(_03035_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_03028_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_1 _09966_ (.A(_03036_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(_03028_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_1 _09968_ (.A(_03037_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_03028_),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_1 _09970_ (.A(_03038_),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_4 _09971_ (.A(_02983_),
    .X(_03039_));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _09973_ (.A(_03040_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_03039_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _09975_ (.A(_03041_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _09976_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(_03039_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _09977_ (.A(_03042_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _09978_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_03039_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _09979_ (.A(_03043_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _09980_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_03039_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_1 _09981_ (.A(_03044_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _09982_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_03039_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _09983_ (.A(_03045_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _09984_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(_03039_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _09985_ (.A(_03046_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _09986_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_03039_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_1 _09987_ (.A(_03047_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _09988_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(_03039_),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _09989_ (.A(_03048_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _09990_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_03039_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _09991_ (.A(_03049_),
    .X(_01280_));
 sky130_fd_sc_hd__clkbuf_4 _09992_ (.A(_02983_),
    .X(_03050_));
 sky130_fd_sc_hd__mux2_1 _09993_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _09994_ (.A(_03051_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _09995_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_03050_),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _09996_ (.A(_03052_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _09997_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_03050_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _09998_ (.A(_03053_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_03050_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _10000_ (.A(_03054_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(\rbzero.tex_g1[63] ),
    .A1(net48),
    .S(_02976_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _10002_ (.A(_03055_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _10003_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[63] ),
    .S(_02976_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _10004_ (.A(_03056_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_02976_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _10006_ (.A(_03057_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(_02976_),
    .X(_03058_));
 sky130_fd_sc_hd__clkbuf_1 _10008_ (.A(_03058_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_02976_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_1 _10010_ (.A(_03059_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_02976_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_1 _10012_ (.A(_03060_),
    .X(_01270_));
 sky130_fd_sc_hd__clkbuf_4 _10013_ (.A(_02909_),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_1 _10014_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_1 _10015_ (.A(_03062_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _10016_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(_03061_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _10017_ (.A(_03063_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _10018_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_03061_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _10019_ (.A(_03064_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _10020_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(_03061_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _10021_ (.A(_03065_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _10022_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_03061_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _10023_ (.A(_03066_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(_03061_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _10025_ (.A(_03067_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_03061_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _10027_ (.A(_03068_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _10028_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(_03061_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _10029_ (.A(_03069_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _10030_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_03061_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _10031_ (.A(_03070_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _10032_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_03061_),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_1 _10033_ (.A(_03071_),
    .X(_01260_));
 sky130_fd_sc_hd__buf_4 _10034_ (.A(_02908_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_4 _10035_ (.A(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_1 _10036_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_1 _10037_ (.A(_03074_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _10038_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(_03073_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_1 _10039_ (.A(_03075_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _10040_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_03073_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _10041_ (.A(_03076_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _10042_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(_03073_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_1 _10043_ (.A(_03077_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _10044_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_03073_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _10045_ (.A(_03078_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(_03073_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _10047_ (.A(_03079_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_03073_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _10049_ (.A(_03080_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _10050_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_03073_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _10051_ (.A(_03081_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _10052_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_03073_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _10053_ (.A(_03082_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _10054_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(_03073_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _10055_ (.A(_03083_),
    .X(_01250_));
 sky130_fd_sc_hd__clkbuf_4 _10056_ (.A(_03072_),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _10058_ (.A(_03085_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _10059_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(_03084_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _10060_ (.A(_03086_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _10061_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_03084_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _10062_ (.A(_03087_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _10063_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(_03084_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_1 _10064_ (.A(_03088_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _10065_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_03084_),
    .X(_03089_));
 sky130_fd_sc_hd__clkbuf_1 _10066_ (.A(_03089_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _10067_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(_03084_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _10068_ (.A(_03090_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _10069_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_03084_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _10070_ (.A(_03091_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _10071_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(_03084_),
    .X(_03092_));
 sky130_fd_sc_hd__clkbuf_1 _10072_ (.A(_03092_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _10073_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_03084_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _10074_ (.A(_03093_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(_03084_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_1 _10076_ (.A(_03094_),
    .X(_01240_));
 sky130_fd_sc_hd__clkbuf_4 _10077_ (.A(_03072_),
    .X(_03095_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _10079_ (.A(_03096_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _10080_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(_03095_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _10081_ (.A(_03097_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_03095_),
    .X(_03098_));
 sky130_fd_sc_hd__clkbuf_1 _10083_ (.A(_03098_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _10084_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(_03095_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _10085_ (.A(_03099_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _10086_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_03095_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _10087_ (.A(_03100_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _10088_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(_03095_),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_1 _10089_ (.A(_03101_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_03095_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _10091_ (.A(_03102_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(_03095_),
    .X(_03103_));
 sky130_fd_sc_hd__clkbuf_1 _10093_ (.A(_03103_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _10094_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_03095_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _10095_ (.A(_03104_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _10096_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(_03095_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _10097_ (.A(_03105_),
    .X(_01230_));
 sky130_fd_sc_hd__clkbuf_4 _10098_ (.A(_03072_),
    .X(_03106_));
 sky130_fd_sc_hd__mux2_1 _10099_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__clkbuf_1 _10100_ (.A(_03107_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _10101_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(_03106_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _10102_ (.A(_03108_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _10103_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_03106_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _10104_ (.A(_03109_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _10105_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(_03106_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _10106_ (.A(_03110_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _10107_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_03106_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _10108_ (.A(_03111_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(_03106_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _10110_ (.A(_03112_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _10111_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_03106_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_1 _10112_ (.A(_03113_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _10113_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(_03106_),
    .X(_03114_));
 sky130_fd_sc_hd__clkbuf_1 _10114_ (.A(_03114_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_03106_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _10116_ (.A(_03115_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(_03106_),
    .X(_03116_));
 sky130_fd_sc_hd__clkbuf_1 _10118_ (.A(_03116_),
    .X(_01220_));
 sky130_fd_sc_hd__buf_4 _10119_ (.A(_03072_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _10120_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _10121_ (.A(_03118_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _10122_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(_03117_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _10123_ (.A(_03119_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_03117_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _10125_ (.A(_03120_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(_03117_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_1 _10127_ (.A(_03121_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _10128_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_03117_),
    .X(_03122_));
 sky130_fd_sc_hd__clkbuf_1 _10129_ (.A(_03122_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(_03117_),
    .X(_03123_));
 sky130_fd_sc_hd__clkbuf_1 _10131_ (.A(_03123_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _10132_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_03117_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_1 _10133_ (.A(_03124_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(\rbzero.tex_g1[0] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_03117_),
    .X(_03125_));
 sky130_fd_sc_hd__clkbuf_1 _10135_ (.A(_03125_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(net48),
    .A1(\rbzero.tex_g0[63] ),
    .S(_03050_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _10137_ (.A(_03126_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_03050_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_1 _10139_ (.A(_03127_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _10140_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(_03050_),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _10141_ (.A(_03128_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_03050_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _10143_ (.A(_03129_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _10144_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_03050_),
    .X(_03130_));
 sky130_fd_sc_hd__clkbuf_1 _10145_ (.A(_03130_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _10146_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_03050_),
    .X(_03131_));
 sky130_fd_sc_hd__clkbuf_1 _10147_ (.A(_03131_),
    .X(_01206_));
 sky130_fd_sc_hd__clkbuf_4 _10148_ (.A(_02983_),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_1 _10149_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__clkbuf_1 _10150_ (.A(_03133_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_03132_),
    .X(_03134_));
 sky130_fd_sc_hd__clkbuf_1 _10152_ (.A(_03134_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(_03132_),
    .X(_03135_));
 sky130_fd_sc_hd__clkbuf_1 _10154_ (.A(_03135_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _10155_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_03132_),
    .X(_03136_));
 sky130_fd_sc_hd__clkbuf_1 _10156_ (.A(_03136_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _10157_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(_03132_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_1 _10158_ (.A(_03137_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _10159_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_03132_),
    .X(_03138_));
 sky130_fd_sc_hd__clkbuf_1 _10160_ (.A(_03138_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(_03132_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_1 _10162_ (.A(_03139_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _10163_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_03132_),
    .X(_03140_));
 sky130_fd_sc_hd__clkbuf_1 _10164_ (.A(_03140_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _10165_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(_03132_),
    .X(_03141_));
 sky130_fd_sc_hd__clkbuf_1 _10166_ (.A(_03141_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _10167_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_03132_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_1 _10168_ (.A(_03142_),
    .X(_01196_));
 sky130_fd_sc_hd__buf_4 _10169_ (.A(_02982_),
    .X(_03143_));
 sky130_fd_sc_hd__clkbuf_4 _10170_ (.A(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_1 _10171_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__clkbuf_1 _10172_ (.A(_03145_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_03144_),
    .X(_03146_));
 sky130_fd_sc_hd__clkbuf_1 _10174_ (.A(_03146_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _10175_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(_03144_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_1 _10176_ (.A(_03147_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _10177_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_03144_),
    .X(_03148_));
 sky130_fd_sc_hd__clkbuf_1 _10178_ (.A(_03148_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _10179_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(_03144_),
    .X(_03149_));
 sky130_fd_sc_hd__clkbuf_1 _10180_ (.A(_03149_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _10181_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_03144_),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_1 _10182_ (.A(_03150_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _10183_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_03144_),
    .X(_03151_));
 sky130_fd_sc_hd__clkbuf_1 _10184_ (.A(_03151_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _10185_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_03144_),
    .X(_03152_));
 sky130_fd_sc_hd__clkbuf_1 _10186_ (.A(_03152_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _10187_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(_03144_),
    .X(_03153_));
 sky130_fd_sc_hd__clkbuf_1 _10188_ (.A(_03153_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _10189_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_03144_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_1 _10190_ (.A(_03154_),
    .X(_01186_));
 sky130_fd_sc_hd__clkbuf_4 _10191_ (.A(_03143_),
    .X(_03155_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__clkbuf_1 _10193_ (.A(_03156_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_03155_),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_1 _10195_ (.A(_03157_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(_03155_),
    .X(_03158_));
 sky130_fd_sc_hd__clkbuf_1 _10197_ (.A(_03158_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_03155_),
    .X(_03159_));
 sky130_fd_sc_hd__clkbuf_1 _10199_ (.A(_03159_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(_03155_),
    .X(_03160_));
 sky130_fd_sc_hd__clkbuf_1 _10201_ (.A(_03160_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_03155_),
    .X(_03161_));
 sky130_fd_sc_hd__clkbuf_1 _10203_ (.A(_03161_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(_03155_),
    .X(_03162_));
 sky130_fd_sc_hd__clkbuf_1 _10205_ (.A(_03162_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_03155_),
    .X(_03163_));
 sky130_fd_sc_hd__clkbuf_1 _10207_ (.A(_03163_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(_03155_),
    .X(_03164_));
 sky130_fd_sc_hd__clkbuf_1 _10209_ (.A(_03164_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_03155_),
    .X(_03165_));
 sky130_fd_sc_hd__clkbuf_1 _10211_ (.A(_03165_),
    .X(_01176_));
 sky130_fd_sc_hd__clkbuf_4 _10212_ (.A(_03143_),
    .X(_03166_));
 sky130_fd_sc_hd__mux2_1 _10213_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__clkbuf_1 _10214_ (.A(_03167_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_03166_),
    .X(_03168_));
 sky130_fd_sc_hd__clkbuf_1 _10216_ (.A(_03168_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(_03166_),
    .X(_03169_));
 sky130_fd_sc_hd__clkbuf_1 _10218_ (.A(_03169_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _10219_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_03166_),
    .X(_03170_));
 sky130_fd_sc_hd__clkbuf_1 _10220_ (.A(_03170_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _10221_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(_03166_),
    .X(_03171_));
 sky130_fd_sc_hd__clkbuf_1 _10222_ (.A(_03171_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _10223_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_03166_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_1 _10224_ (.A(_03172_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _10225_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(_03166_),
    .X(_03173_));
 sky130_fd_sc_hd__clkbuf_1 _10226_ (.A(_03173_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _10227_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_03166_),
    .X(_03174_));
 sky130_fd_sc_hd__clkbuf_1 _10228_ (.A(_03174_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _10229_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(_03166_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_1 _10230_ (.A(_03175_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _10231_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_03166_),
    .X(_03176_));
 sky130_fd_sc_hd__clkbuf_1 _10232_ (.A(_03176_),
    .X(_01166_));
 sky130_fd_sc_hd__clkbuf_4 _10233_ (.A(_03143_),
    .X(_03177_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__clkbuf_1 _10235_ (.A(_03178_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_03177_),
    .X(_03179_));
 sky130_fd_sc_hd__clkbuf_1 _10237_ (.A(_03179_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(_03177_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_1 _10239_ (.A(_03180_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_03177_),
    .X(_03181_));
 sky130_fd_sc_hd__clkbuf_1 _10241_ (.A(_03181_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(_03177_),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_1 _10243_ (.A(_03182_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _10244_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_03177_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_1 _10245_ (.A(_03183_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _10246_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_03177_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_1 _10247_ (.A(_03184_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_03177_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_1 _10249_ (.A(_03185_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(_03177_),
    .X(_03186_));
 sky130_fd_sc_hd__clkbuf_1 _10251_ (.A(_03186_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _10252_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_03177_),
    .X(_03187_));
 sky130_fd_sc_hd__clkbuf_1 _10253_ (.A(_03187_),
    .X(_01156_));
 sky130_fd_sc_hd__buf_4 _10254_ (.A(_03143_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _10255_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__clkbuf_1 _10256_ (.A(_03189_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_03188_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_1 _10258_ (.A(_03190_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _10259_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(_03188_),
    .X(_03191_));
 sky130_fd_sc_hd__clkbuf_1 _10260_ (.A(_03191_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_03188_),
    .X(_03192_));
 sky130_fd_sc_hd__clkbuf_1 _10262_ (.A(_03192_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _10263_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(_03188_),
    .X(_03193_));
 sky130_fd_sc_hd__clkbuf_1 _10264_ (.A(_03193_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_03188_),
    .X(_03194_));
 sky130_fd_sc_hd__clkbuf_1 _10266_ (.A(_03194_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _10267_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_03188_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _10268_ (.A(_03195_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_03188_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _10270_ (.A(_03196_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(\rbzero.tex_b1[63] ),
    .A1(net49),
    .S(_03117_),
    .X(_03197_));
 sky130_fd_sc_hd__clkbuf_1 _10272_ (.A(_03197_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _10273_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[63] ),
    .S(_03117_),
    .X(_03198_));
 sky130_fd_sc_hd__clkbuf_1 _10274_ (.A(_03198_),
    .X(_01146_));
 sky130_fd_sc_hd__clkbuf_4 _10275_ (.A(_03072_),
    .X(_03199_));
 sky130_fd_sc_hd__mux2_1 _10276_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_1 _10277_ (.A(_03200_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(_03199_),
    .X(_03201_));
 sky130_fd_sc_hd__clkbuf_1 _10279_ (.A(_03201_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _10280_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_03199_),
    .X(_03202_));
 sky130_fd_sc_hd__clkbuf_1 _10281_ (.A(_03202_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _10282_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(_03199_),
    .X(_03203_));
 sky130_fd_sc_hd__clkbuf_1 _10283_ (.A(_03203_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_03199_),
    .X(_03204_));
 sky130_fd_sc_hd__clkbuf_1 _10285_ (.A(_03204_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(_03199_),
    .X(_03205_));
 sky130_fd_sc_hd__clkbuf_1 _10287_ (.A(_03205_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_03199_),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_1 _10289_ (.A(_03206_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(_03199_),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_1 _10291_ (.A(_03207_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _10292_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_03199_),
    .X(_03208_));
 sky130_fd_sc_hd__clkbuf_1 _10293_ (.A(_03208_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _10294_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(_03199_),
    .X(_03209_));
 sky130_fd_sc_hd__clkbuf_1 _10295_ (.A(_03209_),
    .X(_01136_));
 sky130_fd_sc_hd__clkbuf_4 _10296_ (.A(_03072_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _10297_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__clkbuf_1 _10298_ (.A(_03211_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _10299_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(_03210_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_1 _10300_ (.A(_03212_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _10301_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_03210_),
    .X(_03213_));
 sky130_fd_sc_hd__clkbuf_1 _10302_ (.A(_03213_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _10303_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(_03210_),
    .X(_03214_));
 sky130_fd_sc_hd__clkbuf_1 _10304_ (.A(_03214_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _10305_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_03210_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_1 _10306_ (.A(_03215_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _10307_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(_03210_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_1 _10308_ (.A(_03216_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _10309_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_03210_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_1 _10310_ (.A(_03217_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _10311_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(_03210_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_1 _10312_ (.A(_03218_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _10313_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_03210_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_1 _10314_ (.A(_03219_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _10315_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(_03210_),
    .X(_03220_));
 sky130_fd_sc_hd__clkbuf_1 _10316_ (.A(_03220_),
    .X(_01126_));
 sky130_fd_sc_hd__clkbuf_4 _10317_ (.A(_03072_),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__clkbuf_1 _10319_ (.A(_03222_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(_03221_),
    .X(_03223_));
 sky130_fd_sc_hd__clkbuf_1 _10321_ (.A(_03223_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_03221_),
    .X(_03224_));
 sky130_fd_sc_hd__clkbuf_1 _10323_ (.A(_03224_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(_03221_),
    .X(_03225_));
 sky130_fd_sc_hd__clkbuf_1 _10325_ (.A(_03225_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _10326_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_03221_),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_1 _10327_ (.A(_03226_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _10328_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(_03221_),
    .X(_03227_));
 sky130_fd_sc_hd__clkbuf_1 _10329_ (.A(_03227_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _10330_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_03221_),
    .X(_03228_));
 sky130_fd_sc_hd__clkbuf_1 _10331_ (.A(_03228_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _10332_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(_03221_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_1 _10333_ (.A(_03229_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _10334_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_03221_),
    .X(_03230_));
 sky130_fd_sc_hd__clkbuf_1 _10335_ (.A(_03230_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(_03221_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_1 _10337_ (.A(_03231_),
    .X(_01116_));
 sky130_fd_sc_hd__clkbuf_4 _10338_ (.A(_03072_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _10339_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__clkbuf_1 _10340_ (.A(_03233_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _10341_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(_03232_),
    .X(_03234_));
 sky130_fd_sc_hd__clkbuf_1 _10342_ (.A(_03234_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _10343_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_03232_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_1 _10344_ (.A(_03235_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _10345_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_03232_),
    .X(_03236_));
 sky130_fd_sc_hd__clkbuf_1 _10346_ (.A(_03236_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _10347_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_03232_),
    .X(_03237_));
 sky130_fd_sc_hd__clkbuf_1 _10348_ (.A(_03237_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _10349_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(_03232_),
    .X(_03238_));
 sky130_fd_sc_hd__clkbuf_1 _10350_ (.A(_03238_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _10351_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_03232_),
    .X(_03239_));
 sky130_fd_sc_hd__clkbuf_1 _10352_ (.A(_03239_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(_03232_),
    .X(_03240_));
 sky130_fd_sc_hd__clkbuf_1 _10354_ (.A(_03240_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _10355_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_03232_),
    .X(_03241_));
 sky130_fd_sc_hd__clkbuf_1 _10356_ (.A(_03241_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _10357_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_03232_),
    .X(_03242_));
 sky130_fd_sc_hd__clkbuf_1 _10358_ (.A(_03242_),
    .X(_01106_));
 sky130_fd_sc_hd__clkbuf_4 _10359_ (.A(_03072_),
    .X(_03243_));
 sky130_fd_sc_hd__mux2_1 _10360_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__clkbuf_1 _10361_ (.A(_03244_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _10362_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(_03243_),
    .X(_03245_));
 sky130_fd_sc_hd__clkbuf_1 _10363_ (.A(_03245_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _10364_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_03243_),
    .X(_03246_));
 sky130_fd_sc_hd__clkbuf_1 _10365_ (.A(_03246_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _10366_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(_03243_),
    .X(_03247_));
 sky130_fd_sc_hd__clkbuf_1 _10367_ (.A(_03247_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _10368_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_03243_),
    .X(_03248_));
 sky130_fd_sc_hd__clkbuf_1 _10369_ (.A(_03248_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _10370_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(_03243_),
    .X(_03249_));
 sky130_fd_sc_hd__clkbuf_1 _10371_ (.A(_03249_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _10372_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_03243_),
    .X(_03250_));
 sky130_fd_sc_hd__clkbuf_1 _10373_ (.A(_03250_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _10374_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_03243_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_1 _10375_ (.A(_03251_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _10376_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_03243_),
    .X(_03252_));
 sky130_fd_sc_hd__clkbuf_1 _10377_ (.A(_03252_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _10378_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(_03243_),
    .X(_03253_));
 sky130_fd_sc_hd__clkbuf_1 _10379_ (.A(_03253_),
    .X(_01096_));
 sky130_fd_sc_hd__clkbuf_4 _10380_ (.A(_02908_),
    .X(_03254_));
 sky130_fd_sc_hd__mux2_1 _10381_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__clkbuf_1 _10382_ (.A(_03255_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _10383_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(_03254_),
    .X(_03256_));
 sky130_fd_sc_hd__clkbuf_1 _10384_ (.A(_03256_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _10385_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_03254_),
    .X(_03257_));
 sky130_fd_sc_hd__clkbuf_1 _10386_ (.A(_03257_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _10387_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_03254_),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_1 _10388_ (.A(_03258_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _10389_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_03254_),
    .X(_03259_));
 sky130_fd_sc_hd__clkbuf_1 _10390_ (.A(_03259_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _10391_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(_03254_),
    .X(_03260_));
 sky130_fd_sc_hd__clkbuf_1 _10392_ (.A(_03260_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _10393_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_03254_),
    .X(_03261_));
 sky130_fd_sc_hd__clkbuf_1 _10394_ (.A(_03261_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _10395_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_03254_),
    .X(_03262_));
 sky130_fd_sc_hd__clkbuf_1 _10396_ (.A(_03262_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _10397_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_03254_),
    .X(_03263_));
 sky130_fd_sc_hd__clkbuf_1 _10398_ (.A(_03263_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _10399_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_03254_),
    .X(_03264_));
 sky130_fd_sc_hd__clkbuf_1 _10400_ (.A(_03264_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _10401_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_02909_),
    .X(_03265_));
 sky130_fd_sc_hd__clkbuf_1 _10402_ (.A(_03265_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _10403_ (.A0(\rbzero.tex_b1[0] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_02909_),
    .X(_03266_));
 sky130_fd_sc_hd__clkbuf_1 _10404_ (.A(_03266_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _10405_ (.A0(net49),
    .A1(\rbzero.tex_b0[63] ),
    .S(_03188_),
    .X(_03267_));
 sky130_fd_sc_hd__clkbuf_1 _10406_ (.A(_03267_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _10407_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_03188_),
    .X(_03268_));
 sky130_fd_sc_hd__clkbuf_1 _10408_ (.A(_03268_),
    .X(_00913_));
 sky130_fd_sc_hd__clkbuf_4 _10409_ (.A(_03143_),
    .X(_03269_));
 sky130_fd_sc_hd__mux2_1 _10410_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__clkbuf_1 _10411_ (.A(_03270_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _10412_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_03269_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_1 _10413_ (.A(_03271_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(_03269_),
    .X(_03272_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_03272_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _10416_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_03269_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_1 _10417_ (.A(_03273_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(_03269_),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_1 _10419_ (.A(_03274_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_03269_),
    .X(_03275_));
 sky130_fd_sc_hd__clkbuf_1 _10421_ (.A(_03275_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(_03269_),
    .X(_03276_));
 sky130_fd_sc_hd__clkbuf_1 _10423_ (.A(_03276_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_03269_),
    .X(_03277_));
 sky130_fd_sc_hd__clkbuf_1 _10425_ (.A(_03277_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(_03269_),
    .X(_03278_));
 sky130_fd_sc_hd__clkbuf_1 _10427_ (.A(_03278_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_03269_),
    .X(_03279_));
 sky130_fd_sc_hd__clkbuf_1 _10429_ (.A(_03279_),
    .X(_00903_));
 sky130_fd_sc_hd__clkbuf_4 _10430_ (.A(_03143_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _10431_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__clkbuf_1 _10432_ (.A(_03281_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _10433_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_03280_),
    .X(_03282_));
 sky130_fd_sc_hd__clkbuf_1 _10434_ (.A(_03282_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(_03280_),
    .X(_03283_));
 sky130_fd_sc_hd__clkbuf_1 _10436_ (.A(_03283_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_03280_),
    .X(_03284_));
 sky130_fd_sc_hd__clkbuf_1 _10438_ (.A(_03284_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(_03280_),
    .X(_03285_));
 sky130_fd_sc_hd__clkbuf_1 _10440_ (.A(_03285_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_03280_),
    .X(_03286_));
 sky130_fd_sc_hd__clkbuf_1 _10442_ (.A(_03286_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_03280_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_1 _10444_ (.A(_03287_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _10445_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_03280_),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_1 _10446_ (.A(_03288_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _10447_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_03280_),
    .X(_03289_));
 sky130_fd_sc_hd__clkbuf_1 _10448_ (.A(_03289_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _10449_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_03280_),
    .X(_03290_));
 sky130_fd_sc_hd__clkbuf_1 _10450_ (.A(_03290_),
    .X(_00893_));
 sky130_fd_sc_hd__clkbuf_4 _10451_ (.A(_03143_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _10452_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__clkbuf_1 _10453_ (.A(_03292_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _10454_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_03291_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_1 _10455_ (.A(_03293_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(_03291_),
    .X(_03294_));
 sky130_fd_sc_hd__clkbuf_1 _10457_ (.A(_03294_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _10458_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_03291_),
    .X(_03295_));
 sky130_fd_sc_hd__clkbuf_1 _10459_ (.A(_03295_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(_03291_),
    .X(_03296_));
 sky130_fd_sc_hd__clkbuf_1 _10461_ (.A(_03296_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_03291_),
    .X(_03297_));
 sky130_fd_sc_hd__clkbuf_1 _10463_ (.A(_03297_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_03291_),
    .X(_03298_));
 sky130_fd_sc_hd__clkbuf_1 _10465_ (.A(_03298_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _10466_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_03291_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_1 _10467_ (.A(_03299_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(_03291_),
    .X(_03300_));
 sky130_fd_sc_hd__clkbuf_1 _10469_ (.A(_03300_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_03291_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_1 _10471_ (.A(_03301_),
    .X(_00883_));
 sky130_fd_sc_hd__clkbuf_4 _10472_ (.A(_03143_),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_1 _10473_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _10474_ (.A(_03303_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_03302_),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_1 _10476_ (.A(_03304_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(_03302_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_1 _10478_ (.A(_03305_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_03302_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _10480_ (.A(_03306_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(_03302_),
    .X(_03307_));
 sky130_fd_sc_hd__clkbuf_1 _10482_ (.A(_03307_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_03302_),
    .X(_03308_));
 sky130_fd_sc_hd__clkbuf_1 _10484_ (.A(_03308_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(_03302_),
    .X(_03309_));
 sky130_fd_sc_hd__clkbuf_1 _10486_ (.A(_03309_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_03302_),
    .X(_03310_));
 sky130_fd_sc_hd__clkbuf_1 _10488_ (.A(_03310_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(_03302_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_1 _10490_ (.A(_03311_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_03302_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_1 _10492_ (.A(_03312_),
    .X(_00873_));
 sky130_fd_sc_hd__clkbuf_4 _10493_ (.A(_03143_),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_1 _10495_ (.A(_03314_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_03313_),
    .X(_03315_));
 sky130_fd_sc_hd__clkbuf_1 _10497_ (.A(_03315_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(_03313_),
    .X(_03316_));
 sky130_fd_sc_hd__clkbuf_1 _10499_ (.A(_03316_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_03313_),
    .X(_03317_));
 sky130_fd_sc_hd__clkbuf_1 _10501_ (.A(_03317_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _10502_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(_03313_),
    .X(_03318_));
 sky130_fd_sc_hd__clkbuf_1 _10503_ (.A(_03318_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _10504_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_03313_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_1 _10505_ (.A(_03319_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(_03313_),
    .X(_03320_));
 sky130_fd_sc_hd__clkbuf_1 _10507_ (.A(_03320_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_03313_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_1 _10509_ (.A(_03321_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_03313_),
    .X(_03322_));
 sky130_fd_sc_hd__clkbuf_1 _10511_ (.A(_03322_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _10512_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_03313_),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_1 _10513_ (.A(_03323_),
    .X(_00863_));
 sky130_fd_sc_hd__clkbuf_4 _10514_ (.A(_02982_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _10516_ (.A(_03325_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_03324_),
    .X(_03326_));
 sky130_fd_sc_hd__clkbuf_1 _10518_ (.A(_03326_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(_03324_),
    .X(_03327_));
 sky130_fd_sc_hd__clkbuf_1 _10520_ (.A(_03327_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_03324_),
    .X(_03328_));
 sky130_fd_sc_hd__clkbuf_1 _10522_ (.A(_03328_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _10523_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(_03324_),
    .X(_03329_));
 sky130_fd_sc_hd__clkbuf_1 _10524_ (.A(_03329_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_03324_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_1 _10526_ (.A(_03330_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _10527_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(_03324_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _10528_ (.A(_03331_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_03324_),
    .X(_03332_));
 sky130_fd_sc_hd__clkbuf_1 _10530_ (.A(_03332_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(_03324_),
    .X(_03333_));
 sky130_fd_sc_hd__clkbuf_1 _10532_ (.A(_03333_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _10533_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_03324_),
    .X(_03334_));
 sky130_fd_sc_hd__clkbuf_1 _10534_ (.A(_03334_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_02983_),
    .X(_03335_));
 sky130_fd_sc_hd__clkbuf_1 _10536_ (.A(_03335_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_02983_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_1 _10538_ (.A(_03336_),
    .X(_00851_));
 sky130_fd_sc_hd__inv_6 _10539_ (.A(\rbzero.vga_sync.vsync ),
    .Y(net72));
 sky130_fd_sc_hd__buf_4 _10540_ (.A(_02981_),
    .X(_03337_));
 sky130_fd_sc_hd__buf_6 _10541_ (.A(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__buf_6 _10542_ (.A(_03338_),
    .X(net61));
 sky130_fd_sc_hd__nand2_4 _10543_ (.A(net72),
    .B(_02907_),
    .Y(_03339_));
 sky130_fd_sc_hd__buf_4 _10544_ (.A(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__clkinv_4 _10545_ (.A(\rbzero.wall_tracer.state[1] ),
    .Y(_03341_));
 sky130_fd_sc_hd__inv_2 _10546_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .Y(_03342_));
 sky130_fd_sc_hd__clkbuf_4 _10547_ (.A(\rbzero.map_rom.f3 ),
    .X(_03343_));
 sky130_fd_sc_hd__inv_2 _10548_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .Y(_03344_));
 sky130_fd_sc_hd__clkbuf_4 _10549_ (.A(\rbzero.map_rom.b6 ),
    .X(_03345_));
 sky130_fd_sc_hd__inv_2 _10550_ (.A(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__inv_2 _10551_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .Y(_03347_));
 sky130_fd_sc_hd__a2bb2o_1 _10552_ (.A1_N(\rbzero.debug_overlay.playerY[2] ),
    .A2_N(_03346_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__a221o_1 _10553_ (.A1(_03342_),
    .A2(_03343_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_03344_),
    .C1(_03348_),
    .X(_03349_));
 sky130_fd_sc_hd__inv_2 _10554_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .Y(_03350_));
 sky130_fd_sc_hd__inv_2 _10555_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .Y(_03351_));
 sky130_fd_sc_hd__clkinv_2 _10556_ (.A(\rbzero.map_rom.d6 ),
    .Y(_03352_));
 sky130_fd_sc_hd__clkbuf_4 _10557_ (.A(\rbzero.map_rom.f2 ),
    .X(_03353_));
 sky130_fd_sc_hd__inv_2 _10558_ (.A(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__a2bb2o_1 _10559_ (.A1_N(\rbzero.debug_overlay.playerY[0] ),
    .A2_N(_03352_),
    .B1(_03354_),
    .B2(\rbzero.debug_overlay.playerX[2] ),
    .X(_03355_));
 sky130_fd_sc_hd__a221o_1 _10560_ (.A1(_03350_),
    .A2(\rbzero.map_rom.i_col[4] ),
    .B1(_03351_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .C1(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__inv_2 _10561_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .Y(_03357_));
 sky130_fd_sc_hd__clkbuf_4 _10562_ (.A(\rbzero.map_rom.c6 ),
    .X(_03358_));
 sky130_fd_sc_hd__inv_2 _10563_ (.A(\rbzero.map_rom.i_row[4] ),
    .Y(_03359_));
 sky130_fd_sc_hd__inv_2 _10564_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .Y(_03360_));
 sky130_fd_sc_hd__a22o_1 _10565_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_03359_),
    .B1(\rbzero.wall_tracer.mapY[5] ),
    .B2(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__clkinv_2 _10566_ (.A(_03343_),
    .Y(_03362_));
 sky130_fd_sc_hd__inv_2 _10567_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .Y(_03363_));
 sky130_fd_sc_hd__clkinv_2 _10568_ (.A(\rbzero.map_rom.i_col[4] ),
    .Y(_03364_));
 sky130_fd_sc_hd__a22o_1 _10569_ (.A1(_03363_),
    .A2(_03353_),
    .B1(_03364_),
    .B2(\rbzero.debug_overlay.playerX[4] ),
    .X(_03365_));
 sky130_fd_sc_hd__a221o_1 _10570_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03362_),
    .B1(_03346_),
    .B2(\rbzero.debug_overlay.playerY[2] ),
    .C1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__a211o_1 _10571_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03361_),
    .C1(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__or3_1 _10572_ (.A(_03349_),
    .B(_03356_),
    .C(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_4 _10573_ (.A(\rbzero.map_rom.f1 ),
    .X(_03369_));
 sky130_fd_sc_hd__nand2_1 _10574_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__or2_1 _10575_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_03369_),
    .X(_03371_));
 sky130_fd_sc_hd__a21o_1 _10576_ (.A1(_03370_),
    .A2(_03371_),
    .B1(\rbzero.wall_tracer.mapY[7] ),
    .X(_03372_));
 sky130_fd_sc_hd__inv_2 _10577_ (.A(\rbzero.map_rom.f4 ),
    .Y(_03373_));
 sky130_fd_sc_hd__inv_2 _10578_ (.A(_03358_),
    .Y(_03374_));
 sky130_fd_sc_hd__clkinv_2 _10579_ (.A(\rbzero.map_rom.a6 ),
    .Y(_03375_));
 sky130_fd_sc_hd__a22o_1 _10580_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_03352_),
    .B1(_03375_),
    .B2(\rbzero.debug_overlay.playerY[3] ),
    .X(_03376_));
 sky130_fd_sc_hd__a221o_1 _10581_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\rbzero.debug_overlay.playerY[1] ),
    .C1(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__inv_2 _10582_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .Y(_03378_));
 sky130_fd_sc_hd__a211oi_1 _10583_ (.A1(_03378_),
    .A2(\rbzero.wall_tracer.mapX[5] ),
    .B1(\rbzero.wall_tracer.mapX[7] ),
    .C1(\rbzero.wall_tracer.mapX[6] ),
    .Y(_03379_));
 sky130_fd_sc_hd__o221ai_1 _10584_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03373_),
    .B1(\rbzero.wall_tracer.mapX[5] ),
    .B2(_03378_),
    .C1(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__or4_1 _10585_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(\rbzero.wall_tracer.mapY[9] ),
    .C(\rbzero.wall_tracer.mapY[8] ),
    .D(\rbzero.wall_tracer.mapY[10] ),
    .X(_03381_));
 sky130_fd_sc_hd__or4_1 _10586_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(\rbzero.wall_tracer.mapX[8] ),
    .C(\rbzero.wall_tracer.mapX[10] ),
    .D(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__or4_1 _10587_ (.A(_03372_),
    .B(_03377_),
    .C(_03380_),
    .D(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__or4_1 _10588_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(\rbzero.wall_tracer.visualWallDist[6] ),
    .C(\rbzero.wall_tracer.visualWallDist[5] ),
    .D(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_03384_));
 sky130_fd_sc_hd__or4_1 _10589_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(\rbzero.wall_tracer.visualWallDist[2] ),
    .C(\rbzero.wall_tracer.visualWallDist[1] ),
    .D(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_03385_));
 sky130_fd_sc_hd__or4_1 _10590_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(\rbzero.wall_tracer.visualWallDist[-2] ),
    .C(\rbzero.wall_tracer.visualWallDist[-3] ),
    .D(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__or4_1 _10591_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(\rbzero.wall_tracer.visualWallDist[8] ),
    .C(_03384_),
    .D(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__inv_2 _10592_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .Y(_03388_));
 sky130_fd_sc_hd__o211a_1 _10593_ (.A1(_03368_),
    .A2(_03383_),
    .B1(_03387_),
    .C1(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_4 _10594_ (.A(\rbzero.map_rom.d6 ),
    .X(_03390_));
 sky130_fd_sc_hd__nand2_1 _10595_ (.A(_03390_),
    .B(_03358_),
    .Y(_03391_));
 sky130_fd_sc_hd__or2_1 _10596_ (.A(_03390_),
    .B(_03358_),
    .X(_03392_));
 sky130_fd_sc_hd__nand2_1 _10597_ (.A(_03391_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__a22o_1 _10598_ (.A1(_03373_),
    .A2(_03352_),
    .B1(_03393_),
    .B2(_03343_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_4 _10599_ (.A(\rbzero.map_rom.f4 ),
    .X(_03395_));
 sky130_fd_sc_hd__and3_1 _10600_ (.A(\rbzero.map_rom.f2 ),
    .B(\rbzero.map_rom.f1 ),
    .C(\rbzero.map_rom.i_col[4] ),
    .X(_03396_));
 sky130_fd_sc_hd__nor4_1 _10601_ (.A(_03346_),
    .B(_03375_),
    .C(_03359_),
    .D(_03391_),
    .Y(_03397_));
 sky130_fd_sc_hd__a31o_1 _10602_ (.A1(_03395_),
    .A2(_03343_),
    .A3(_03396_),
    .B1(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__or2_1 _10603_ (.A(\rbzero.map_rom.f2 ),
    .B(\rbzero.map_rom.b6 ),
    .X(_03399_));
 sky130_fd_sc_hd__xnor2_1 _10604_ (.A(_03343_),
    .B(_03358_),
    .Y(_03400_));
 sky130_fd_sc_hd__o21ai_1 _10605_ (.A1(_03373_),
    .A2(_03352_),
    .B1(_03399_),
    .Y(_03401_));
 sky130_fd_sc_hd__a2111o_1 _10606_ (.A1(_03373_),
    .A2(_03352_),
    .B1(\rbzero.map_rom.a6 ),
    .C1(_03401_),
    .D1(\rbzero.map_rom.f1 ),
    .X(_03402_));
 sky130_fd_sc_hd__a211o_1 _10607_ (.A1(_03353_),
    .A2(_03345_),
    .B1(_03400_),
    .C1(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__or4_1 _10608_ (.A(_03345_),
    .B(\rbzero.map_rom.a6 ),
    .C(\rbzero.map_rom.i_row[4] ),
    .D(_03392_),
    .X(_03404_));
 sky130_fd_sc_hd__o311a_1 _10609_ (.A1(_03395_),
    .A2(_03390_),
    .A3(_03399_),
    .B1(_03403_),
    .C1(_03404_),
    .X(_03405_));
 sky130_fd_sc_hd__or2_1 _10610_ (.A(_03395_),
    .B(_03343_),
    .X(_03406_));
 sky130_fd_sc_hd__or4_1 _10611_ (.A(_03353_),
    .B(_03369_),
    .C(\rbzero.map_rom.i_col[4] ),
    .D(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__nand3b_1 _10612_ (.A_N(_03398_),
    .B(_03405_),
    .C(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__a31o_1 _10613_ (.A1(_03353_),
    .A2(_03345_),
    .A3(_03394_),
    .B1(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__or4_1 _10614_ (.A(\rbzero.map_rom.i_col[4] ),
    .B(_03390_),
    .C(_03375_),
    .D(\rbzero.map_rom.i_row[4] ),
    .X(_03410_));
 sky130_fd_sc_hd__nand2_1 _10615_ (.A(_03369_),
    .B(_03358_),
    .Y(_03411_));
 sky130_fd_sc_hd__or4_1 _10616_ (.A(_03406_),
    .B(_03399_),
    .C(_03410_),
    .D(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__inv_2 _10617_ (.A(_03369_),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_1 _10618_ (.A(_03343_),
    .B(_03390_),
    .Y(_03414_));
 sky130_fd_sc_hd__a221o_1 _10619_ (.A1(_03413_),
    .A2(_03374_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(_03353_),
    .C1(_03414_),
    .X(_03415_));
 sky130_fd_sc_hd__a22o_1 _10620_ (.A1(_03395_),
    .A2(_03345_),
    .B1(_03375_),
    .B2(_03354_),
    .X(_03416_));
 sky130_fd_sc_hd__o21ai_1 _10621_ (.A1(_03395_),
    .A2(_03345_),
    .B1(_03411_),
    .Y(_03417_));
 sky130_fd_sc_hd__or3_1 _10622_ (.A(_03415_),
    .B(_03416_),
    .C(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__nand2_1 _10623_ (.A(_03412_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__inv_2 _10624_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .Y(_03420_));
 sky130_fd_sc_hd__or4_1 _10625_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(\rbzero.map_overlay.i_mapdx[2] ),
    .C(\rbzero.map_overlay.i_mapdx[1] ),
    .D(\rbzero.map_overlay.i_mapdx[0] ),
    .X(_03421_));
 sky130_fd_sc_hd__a21o_1 _10626_ (.A1(_03420_),
    .A2(_03421_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .X(_03422_));
 sky130_fd_sc_hd__o2bb2a_1 _10627_ (.A1_N(\rbzero.map_overlay.i_mapdx[3] ),
    .A2_N(_03413_),
    .B1(_03373_),
    .B2(\rbzero.map_overlay.i_mapdx[0] ),
    .X(_03423_));
 sky130_fd_sc_hd__xnor2_1 _10628_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_03353_),
    .Y(_03424_));
 sky130_fd_sc_hd__inv_2 _10629_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .Y(_03425_));
 sky130_fd_sc_hd__xnor2_1 _10630_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .B(_03343_),
    .Y(_03426_));
 sky130_fd_sc_hd__o221a_1 _10631_ (.A1(_03425_),
    .A2(_03395_),
    .B1(_03364_),
    .B2(\rbzero.map_overlay.i_mapdx[4] ),
    .C1(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__o2111a_1 _10632_ (.A1(\rbzero.map_overlay.i_mapdx[3] ),
    .A2(_03413_),
    .B1(_03423_),
    .C1(_03424_),
    .D1(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__and2_1 _10633_ (.A(_03422_),
    .B(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__inv_2 _10634_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .Y(_03430_));
 sky130_fd_sc_hd__xor2_1 _10635_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .B(_03369_),
    .X(_03431_));
 sky130_fd_sc_hd__a221o_1 _10636_ (.A1(_03430_),
    .A2(_03343_),
    .B1(_03352_),
    .B2(\rbzero.map_overlay.i_othery[0] ),
    .C1(_03431_),
    .X(_03432_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(\rbzero.map_overlay.i_othery[2] ),
    .B(_03345_),
    .Y(_03433_));
 sky130_fd_sc_hd__or2_1 _10638_ (.A(\rbzero.map_overlay.i_othery[2] ),
    .B(_03345_),
    .X(_03434_));
 sky130_fd_sc_hd__xor2_1 _10639_ (.A(\rbzero.map_overlay.i_othery[3] ),
    .B(\rbzero.map_rom.a6 ),
    .X(_03435_));
 sky130_fd_sc_hd__xor2_1 _10640_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .B(\rbzero.map_rom.i_row[4] ),
    .X(_03436_));
 sky130_fd_sc_hd__inv_2 _10641_ (.A(\rbzero.map_overlay.i_othery[0] ),
    .Y(_03437_));
 sky130_fd_sc_hd__xor2_1 _10642_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(_03358_),
    .X(_03438_));
 sky130_fd_sc_hd__a221o_1 _10643_ (.A1(\rbzero.map_overlay.i_otherx[4] ),
    .A2(_03364_),
    .B1(_03390_),
    .B2(_03437_),
    .C1(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__xor2_1 _10644_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .B(\rbzero.map_rom.f2 ),
    .X(_03440_));
 sky130_fd_sc_hd__inv_2 _10645_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .Y(_03441_));
 sky130_fd_sc_hd__xor2_1 _10646_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(_03395_),
    .X(_03442_));
 sky130_fd_sc_hd__a221o_1 _10647_ (.A1(\rbzero.map_overlay.i_otherx[1] ),
    .A2(_03362_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .B2(_03441_),
    .C1(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__or4_1 _10648_ (.A(_03436_),
    .B(_03439_),
    .C(_03440_),
    .D(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__a211o_1 _10649_ (.A1(_03433_),
    .A2(_03434_),
    .B1(_03435_),
    .C1(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__inv_2 _10650_ (.A(\rbzero.map_overlay.i_mapdy[1] ),
    .Y(_03446_));
 sky130_fd_sc_hd__inv_2 _10651_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .Y(_03447_));
 sky130_fd_sc_hd__xnor2_1 _10652_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(\rbzero.map_rom.b6 ),
    .Y(_03448_));
 sky130_fd_sc_hd__o221a_1 _10653_ (.A1(_03446_),
    .A2(_03358_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(_03447_),
    .C1(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__o221a_1 _10654_ (.A1(\rbzero.map_overlay.i_mapdy[1] ),
    .A2(_03374_),
    .B1(_03359_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__inv_2 _10655_ (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .Y(_03451_));
 sky130_fd_sc_hd__xnor2_1 _10656_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(_03390_),
    .Y(_03452_));
 sky130_fd_sc_hd__o221a_1 _10657_ (.A1(\rbzero.map_overlay.i_mapdy[3] ),
    .A2(_03375_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_03451_),
    .C1(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__and3_1 _10658_ (.A(_03404_),
    .B(_03450_),
    .C(_03453_),
    .X(_03454_));
 sky130_fd_sc_hd__o21ba_1 _10659_ (.A1(_03432_),
    .A2(_03445_),
    .B1_N(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__or4b_1 _10660_ (.A(_03409_),
    .B(_03419_),
    .C(_03429_),
    .D_N(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__nand2_2 _10661_ (.A(_03389_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__or2_4 _10662_ (.A(_03341_),
    .B(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__nor2_2 _10663_ (.A(_03340_),
    .B(_03458_),
    .Y(_00016_));
 sky130_fd_sc_hd__clkbuf_4 _10664_ (.A(_02902_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_4 _10665_ (.A(\gpout0.hpos[5] ),
    .X(_03460_));
 sky130_fd_sc_hd__buf_2 _10666_ (.A(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__inv_2 _10667_ (.A(\gpout0.hpos[3] ),
    .Y(_03462_));
 sky130_fd_sc_hd__inv_2 _10668_ (.A(\gpout0.hpos[4] ),
    .Y(_03463_));
 sky130_fd_sc_hd__buf_4 _10669_ (.A(_03463_),
    .X(_03464_));
 sky130_fd_sc_hd__nor2_1 _10670_ (.A(_03462_),
    .B(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__buf_4 _10671_ (.A(\gpout0.hpos[6] ),
    .X(_03466_));
 sky130_fd_sc_hd__or2_2 _10672_ (.A(_02900_),
    .B(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__o31a_1 _10673_ (.A1(_03461_),
    .A2(_02901_),
    .A3(_03465_),
    .B1(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_4 _10674_ (.A(\gpout0.hpos[9] ),
    .X(_03469_));
 sky130_fd_sc_hd__o21ai_1 _10675_ (.A1(_02902_),
    .A2(_03468_),
    .B1(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__a21o_1 _10676_ (.A1(_03459_),
    .A2(_03468_),
    .B1(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__nor2_1 _10677_ (.A(_03461_),
    .B(_03465_),
    .Y(_03472_));
 sky130_fd_sc_hd__inv_2 _10678_ (.A(\gpout0.hpos[6] ),
    .Y(_03473_));
 sky130_fd_sc_hd__buf_4 _10679_ (.A(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__or3_1 _10680_ (.A(_02901_),
    .B(_03474_),
    .C(_02902_),
    .X(_03475_));
 sky130_fd_sc_hd__and3_1 _10681_ (.A(\gpout0.hpos[3] ),
    .B(\gpout0.hpos[4] ),
    .C(\gpout0.hpos[5] ),
    .X(_03476_));
 sky130_fd_sc_hd__or4_1 _10682_ (.A(_03471_),
    .B(_03472_),
    .C(_03475_),
    .D(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__buf_6 _10683_ (.A(_03477_),
    .X(net69));
 sky130_fd_sc_hd__nand2_2 _10684_ (.A(_02904_),
    .B(_03468_),
    .Y(net68));
 sky130_fd_sc_hd__inv_2 _10685_ (.A(\rbzero.wall_tracer.state[11] ),
    .Y(_03478_));
 sky130_fd_sc_hd__nor2_1 _10686_ (.A(_03478_),
    .B(_03340_),
    .Y(_00000_));
 sky130_fd_sc_hd__clkbuf_4 _10687_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_03479_));
 sky130_fd_sc_hd__buf_2 _10688_ (.A(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__inv_2 _10689_ (.A(\rbzero.wall_tracer.state[8] ),
    .Y(_03481_));
 sky130_fd_sc_hd__inv_2 _10690_ (.A(\rbzero.wall_tracer.state[0] ),
    .Y(_03482_));
 sky130_fd_sc_hd__nor2_2 _10691_ (.A(\rbzero.vga_sync.vsync ),
    .B(_02981_),
    .Y(_03483_));
 sky130_fd_sc_hd__buf_6 _10692_ (.A(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__buf_6 _10693_ (.A(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__a41o_1 _10694_ (.A1(_03480_),
    .A2(_03481_),
    .A3(_03482_),
    .A4(_03485_),
    .B1(_00000_),
    .X(_00012_));
 sky130_fd_sc_hd__buf_4 _10695_ (.A(_03340_),
    .X(_03486_));
 sky130_fd_sc_hd__nor2_1 _10696_ (.A(_03482_),
    .B(_03486_),
    .Y(_00005_));
 sky130_fd_sc_hd__buf_2 _10697_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_03487_));
 sky130_fd_sc_hd__clkbuf_4 _10698_ (.A(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_4 _10699_ (.A(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__a311o_1 _10700_ (.A1(_03489_),
    .A2(_03481_),
    .A3(_03478_),
    .B1(_03486_),
    .C1(\rbzero.wall_tracer.state[0] ),
    .X(_00011_));
 sky130_fd_sc_hd__clkbuf_4 _10701_ (.A(\rbzero.wall_tracer.state[13] ),
    .X(_03490_));
 sky130_fd_sc_hd__buf_4 _10702_ (.A(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_4 _10703_ (.A(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__buf_4 _10704_ (.A(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__and2_1 _10705_ (.A(\rbzero.wall_tracer.state[1] ),
    .B(_03457_),
    .X(_03494_));
 sky130_fd_sc_hd__buf_2 _10706_ (.A(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_4 _10707_ (.A(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__buf_6 _10708_ (.A(_03484_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_4 _10709_ (.A(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__o21a_1 _10710_ (.A1(_03493_),
    .A2(_03496_),
    .B1(_03498_),
    .X(_00015_));
 sky130_fd_sc_hd__inv_2 _10711_ (.A(\gpout0.hpos[1] ),
    .Y(_03499_));
 sky130_fd_sc_hd__inv_2 _10712_ (.A(\gpout0.hpos[0] ),
    .Y(_03500_));
 sky130_fd_sc_hd__nor2_1 _10713_ (.A(_03499_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__nand2_1 _10714_ (.A(\gpout0.hpos[2] ),
    .B(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__nor2_1 _10715_ (.A(_03462_),
    .B(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__o21a_1 _10716_ (.A1(_02900_),
    .A2(\gpout0.hpos[8] ),
    .B1(\gpout0.hpos[9] ),
    .X(_03504_));
 sky130_fd_sc_hd__nor2_1 _10717_ (.A(_03464_),
    .B(_03461_),
    .Y(_03505_));
 sky130_fd_sc_hd__and4b_4 _10718_ (.A_N(_03467_),
    .B(_03503_),
    .C(_03504_),
    .D(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__nand2_1 _10719_ (.A(\rbzero.wall_tracer.state[14] ),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__and2_1 _10720_ (.A(_03484_),
    .B(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__clkinv_4 _10721_ (.A(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__buf_4 _10722_ (.A(_03509_),
    .X(_00013_));
 sky130_fd_sc_hd__and2b_1 _10723_ (.A_N(_03506_),
    .B(\rbzero.wall_tracer.state[14] ),
    .X(_03510_));
 sky130_fd_sc_hd__o21a_1 _10724_ (.A1(\rbzero.wall_tracer.state[10] ),
    .A2(_03510_),
    .B1(_03498_),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _10725_ (.A(\gpout0.hpos[4] ),
    .B(_03503_),
    .X(_03511_));
 sky130_fd_sc_hd__o21a_1 _10726_ (.A1(\gpout0.hpos[5] ),
    .A2(_03511_),
    .B1(\gpout0.hpos[6] ),
    .X(_03512_));
 sky130_fd_sc_hd__and2_1 _10727_ (.A(\gpout0.hpos[7] ),
    .B(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__a21oi_2 _10728_ (.A1(\gpout0.hpos[8] ),
    .A2(_03513_),
    .B1(\gpout0.hpos[9] ),
    .Y(_03514_));
 sky130_fd_sc_hd__buf_4 _10729_ (.A(\gpout0.vpos[7] ),
    .X(_03515_));
 sky130_fd_sc_hd__or4b_1 _10730_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.vpos[8] ),
    .C(_03515_),
    .D_N(net2),
    .X(_03516_));
 sky130_fd_sc_hd__clkbuf_4 _10731_ (.A(\gpout0.vpos[3] ),
    .X(_03517_));
 sky130_fd_sc_hd__or3_2 _10732_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(\gpout0.vpos[0] ),
    .X(_03518_));
 sky130_fd_sc_hd__or2_2 _10733_ (.A(\gpout0.vpos[5] ),
    .B(\gpout0.vpos[4] ),
    .X(_03519_));
 sky130_fd_sc_hd__clkbuf_4 _10734_ (.A(\gpout0.vpos[6] ),
    .X(_03520_));
 sky130_fd_sc_hd__o31a_1 _10735_ (.A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .B1(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__nor3_4 _10736_ (.A(_03514_),
    .B(_03516_),
    .C(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__clkbuf_4 _10737_ (.A(\gpout0.hpos[3] ),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_4 _10738_ (.A(\gpout0.hpos[4] ),
    .X(_03524_));
 sky130_fd_sc_hd__or2_1 _10739_ (.A(_03523_),
    .B(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__buf_2 _10740_ (.A(\gpout0.hpos[2] ),
    .X(_03526_));
 sky130_fd_sc_hd__buf_2 _10741_ (.A(\gpout0.hpos[1] ),
    .X(_03527_));
 sky130_fd_sc_hd__or2_1 _10742_ (.A(_03526_),
    .B(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__or2_1 _10743_ (.A(\gpout0.hpos[0] ),
    .B(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__o41a_1 _10744_ (.A1(_03461_),
    .A2(_03467_),
    .A3(_03525_),
    .A4(_03529_),
    .B1(_02902_),
    .X(_03530_));
 sky130_fd_sc_hd__or3_1 _10745_ (.A(\gpout0.vpos[7] ),
    .B(\gpout0.vpos[6] ),
    .C(_03519_),
    .X(_03531_));
 sky130_fd_sc_hd__o31a_1 _10746_ (.A1(_03517_),
    .A2(_03518_),
    .A3(_03531_),
    .B1(\gpout0.vpos[8] ),
    .X(_03532_));
 sky130_fd_sc_hd__or3b_1 _10747_ (.A(\gpout0.vpos[9] ),
    .B(_03469_),
    .C_N(net1),
    .X(_03533_));
 sky130_fd_sc_hd__nor3_2 _10748_ (.A(_03530_),
    .B(_03532_),
    .C(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__a21oi_4 _10749_ (.A1(_02902_),
    .A2(_03467_),
    .B1(\gpout0.hpos[9] ),
    .Y(_03535_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__buf_4 _10751_ (.A(net41),
    .X(_03537_));
 sky130_fd_sc_hd__inv_2 _10752_ (.A(\rbzero.row_render.side ),
    .Y(_03538_));
 sky130_fd_sc_hd__clkinv_2 _10753_ (.A(\rbzero.row_render.wall[0] ),
    .Y(_03539_));
 sky130_fd_sc_hd__nor2_1 _10754_ (.A(_03539_),
    .B(\rbzero.row_render.wall[1] ),
    .Y(_03540_));
 sky130_fd_sc_hd__nand2_1 _10755_ (.A(_03538_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__nand2_1 _10756_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .Y(_03542_));
 sky130_fd_sc_hd__or2_1 _10757_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .X(_03543_));
 sky130_fd_sc_hd__nand3_1 _10758_ (.A(\rbzero.texV[4] ),
    .B(_03542_),
    .C(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21o_1 _10759_ (.A1(_03542_),
    .A2(_03543_),
    .B1(\rbzero.texV[4] ),
    .X(_03545_));
 sky130_fd_sc_hd__nand2_1 _10760_ (.A(_03544_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__or2_1 _10761_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .X(_03547_));
 sky130_fd_sc_hd__nand2_1 _10762_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .Y(_03548_));
 sky130_fd_sc_hd__a21boi_2 _10763_ (.A1(\rbzero.texV[3] ),
    .A2(_03547_),
    .B1_N(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__nor2_1 _10764_ (.A(_03546_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand2_1 _10765_ (.A(_03548_),
    .B(_03547_),
    .Y(_03551_));
 sky130_fd_sc_hd__xor2_1 _10766_ (.A(\rbzero.texV[3] ),
    .B(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__o211a_1 _10767_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(\rbzero.texV[1] ),
    .B1(\rbzero.texV[0] ),
    .C1(\rbzero.traced_texVinit[0] ),
    .X(_03553_));
 sky130_fd_sc_hd__a221o_1 _10768_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(\rbzero.texV[1] ),
    .B2(\rbzero.traced_texVinit[1] ),
    .C1(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__o21ai_2 _10769_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__or2_2 _10770_ (.A(_03552_),
    .B(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__xnor2_1 _10771_ (.A(_03546_),
    .B(_03549_),
    .Y(_03557_));
 sky130_fd_sc_hd__nor2_2 _10772_ (.A(_03556_),
    .B(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__and2_1 _10773_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .X(_03559_));
 sky130_fd_sc_hd__nor2_1 _10774_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .Y(_03560_));
 sky130_fd_sc_hd__nor2_1 _10775_ (.A(_03559_),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__xnor2_1 _10776_ (.A(\rbzero.texV[5] ),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__a21oi_1 _10777_ (.A1(_03542_),
    .A2(_03544_),
    .B1(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__and3_1 _10778_ (.A(_03562_),
    .B(_03542_),
    .C(_03544_),
    .X(_03564_));
 sky130_fd_sc_hd__or2_1 _10779_ (.A(_03563_),
    .B(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__inv_2 _10780_ (.A(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__o21a_1 _10781_ (.A1(_03550_),
    .A2(_03558_),
    .B1(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__nand2_1 _10782_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_03568_));
 sky130_fd_sc_hd__xor2_1 _10783_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .X(_03569_));
 sky130_fd_sc_hd__xnor2_1 _10784_ (.A(_03568_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .X(_03571_));
 sky130_fd_sc_hd__nand2_1 _10786_ (.A(_03568_),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__or2_1 _10787_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .X(_03573_));
 sky130_fd_sc_hd__nand2_1 _10788_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .Y(_03574_));
 sky130_fd_sc_hd__a21boi_1 _10789_ (.A1(\rbzero.texV[8] ),
    .A2(_03573_),
    .B1_N(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__nor2_1 _10790_ (.A(_03572_),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__nand2_1 _10791_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .Y(_03577_));
 sky130_fd_sc_hd__or2_1 _10792_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .X(_03578_));
 sky130_fd_sc_hd__nand3_1 _10793_ (.A(\rbzero.texV[7] ),
    .B(_03577_),
    .C(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand2_1 _10794_ (.A(_03574_),
    .B(_03573_),
    .Y(_03580_));
 sky130_fd_sc_hd__xor2_1 _10795_ (.A(\rbzero.texV[8] ),
    .B(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__a21oi_1 _10796_ (.A1(_03577_),
    .A2(_03579_),
    .B1(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__and3_1 _10797_ (.A(_03581_),
    .B(_03577_),
    .C(_03579_),
    .X(_03583_));
 sky130_fd_sc_hd__a21o_1 _10798_ (.A1(_03577_),
    .A2(_03578_),
    .B1(\rbzero.texV[7] ),
    .X(_03584_));
 sky130_fd_sc_hd__nand2_1 _10799_ (.A(_03579_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__nand2_1 _10800_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .Y(_03586_));
 sky130_fd_sc_hd__or2_1 _10801_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .X(_03587_));
 sky130_fd_sc_hd__nand3_1 _10802_ (.A(\rbzero.texV[6] ),
    .B(_03586_),
    .C(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__nand3_1 _10803_ (.A(_03585_),
    .B(_03586_),
    .C(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__a21o_1 _10804_ (.A1(_03586_),
    .A2(_03587_),
    .B1(\rbzero.texV[6] ),
    .X(_03590_));
 sky130_fd_sc_hd__nand2_1 _10805_ (.A(_03588_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__a21oi_2 _10806_ (.A1(\rbzero.texV[5] ),
    .A2(_03561_),
    .B1(_03559_),
    .Y(_03592_));
 sky130_fd_sc_hd__xnor2_1 _10807_ (.A(_03591_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__nor2_1 _10808_ (.A(_03563_),
    .B(_03567_),
    .Y(_03594_));
 sky130_fd_sc_hd__nor2_1 _10809_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__o21bai_2 _10810_ (.A1(_03591_),
    .A2(_03592_),
    .B1_N(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__a21oi_1 _10811_ (.A1(_03586_),
    .A2(_03588_),
    .B1(_03585_),
    .Y(_03597_));
 sky130_fd_sc_hd__a21oi_1 _10812_ (.A1(_03589_),
    .A2(_03596_),
    .B1(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__nor2_1 _10813_ (.A(_03583_),
    .B(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(_03572_),
    .B(_03575_),
    .Y(_03600_));
 sky130_fd_sc_hd__o31a_1 _10815_ (.A1(_03576_),
    .A2(_03582_),
    .A3(_03599_),
    .B1(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__a21oi_1 _10816_ (.A1(_03570_),
    .A2(_03601_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_03602_));
 sky130_fd_sc_hd__o21a_4 _10817_ (.A1(_03570_),
    .A2(_03601_),
    .B1(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__nor3_1 _10818_ (.A(_03566_),
    .B(_03550_),
    .C(_03558_),
    .Y(_03604_));
 sky130_fd_sc_hd__or3_1 _10819_ (.A(_03567_),
    .B(_03603_),
    .C(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__buf_4 _10820_ (.A(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__buf_6 _10821_ (.A(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__nand2_1 _10822_ (.A(_03556_),
    .B(_03557_),
    .Y(_03608_));
 sky130_fd_sc_hd__or3b_1 _10823_ (.A(_03558_),
    .B(_03603_),
    .C_N(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__buf_4 _10824_ (.A(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__buf_4 _10825_ (.A(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__buf_6 _10826_ (.A(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__a21oi_2 _10827_ (.A1(_03552_),
    .A2(_03555_),
    .B1(_03603_),
    .Y(_03613_));
 sky130_fd_sc_hd__nand2_4 _10828_ (.A(_03556_),
    .B(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__buf_4 _10829_ (.A(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__buf_6 _10830_ (.A(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__clkbuf_8 _10831_ (.A(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__buf_4 _10832_ (.A(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__a41o_1 _10833_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_03607_),
    .A3(_03612_),
    .A4(_03618_),
    .B1(_03538_),
    .X(_03619_));
 sky130_fd_sc_hd__and2_2 _10834_ (.A(_03556_),
    .B(_03613_),
    .X(_03620_));
 sky130_fd_sc_hd__nor2_1 _10835_ (.A(\rbzero.row_render.texu[0] ),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__and2_1 _10836_ (.A(_03593_),
    .B(_03594_),
    .X(_03622_));
 sky130_fd_sc_hd__or3_1 _10837_ (.A(_03595_),
    .B(_03603_),
    .C(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__buf_6 _10838_ (.A(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__nand2_1 _10839_ (.A(\rbzero.row_render.texu[4] ),
    .B(\rbzero.row_render.texu[3] ),
    .Y(_03625_));
 sky130_fd_sc_hd__or4_1 _10840_ (.A(\rbzero.row_render.texu[2] ),
    .B(\rbzero.row_render.texu[1] ),
    .C(_03624_),
    .D(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__nor3_4 _10841_ (.A(_03595_),
    .B(_03603_),
    .C(_03622_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand2_1 _10842_ (.A(\rbzero.row_render.texu[2] ),
    .B(\rbzero.row_render.texu[1] ),
    .Y(_03628_));
 sky130_fd_sc_hd__or4_1 _10843_ (.A(\rbzero.row_render.texu[4] ),
    .B(\rbzero.row_render.texu[3] ),
    .C(_03627_),
    .D(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__a21oi_1 _10844_ (.A1(_03626_),
    .A2(_03629_),
    .B1(\rbzero.row_render.texu[0] ),
    .Y(_03630_));
 sky130_fd_sc_hd__a31o_1 _10845_ (.A1(_03606_),
    .A2(_03611_),
    .A3(_03621_),
    .B1(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__and2_1 _10846_ (.A(_03539_),
    .B(\rbzero.row_render.wall[1] ),
    .X(_03632_));
 sky130_fd_sc_hd__o21a_1 _10847_ (.A1(\rbzero.row_render.side ),
    .A2(_03631_),
    .B1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__nor3_4 _10848_ (.A(_03567_),
    .B(_03603_),
    .C(_03604_),
    .Y(_03634_));
 sky130_fd_sc_hd__nor3b_4 _10849_ (.A(_03558_),
    .B(_03603_),
    .C_N(_03608_),
    .Y(_03635_));
 sky130_fd_sc_hd__or3_1 _10850_ (.A(_03627_),
    .B(_03634_),
    .C(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__nand3_1 _10851_ (.A(\rbzero.row_render.texu[3] ),
    .B(\rbzero.row_render.texu[2] ),
    .C(\rbzero.row_render.texu[1] ),
    .Y(_03637_));
 sky130_fd_sc_hd__a21bo_1 _10852_ (.A1(_03636_),
    .A2(_03637_),
    .B1_N(\rbzero.row_render.wall[1] ),
    .X(_03638_));
 sky130_fd_sc_hd__nand2_1 _10853_ (.A(_03634_),
    .B(_03635_),
    .Y(_03639_));
 sky130_fd_sc_hd__o32a_1 _10854_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(\rbzero.row_render.texu[2] ),
    .A3(\rbzero.row_render.texu[1] ),
    .B1(_03624_),
    .B2(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__nand2_1 _10855_ (.A(\rbzero.row_render.wall[0] ),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__nor2_1 _10856_ (.A(\rbzero.row_render.side ),
    .B(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__inv_2 _10857_ (.A(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__o21ai_1 _10858_ (.A1(_03638_),
    .A2(_03641_),
    .B1(\rbzero.row_render.side ),
    .Y(_03644_));
 sky130_fd_sc_hd__o21a_1 _10859_ (.A1(_03638_),
    .A2(_03643_),
    .B1(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__nor2_1 _10860_ (.A(_03632_),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__a211o_1 _10861_ (.A1(_03619_),
    .A2(_03633_),
    .B1(_03646_),
    .C1(_03540_),
    .X(_03647_));
 sky130_fd_sc_hd__buf_4 _10862_ (.A(_03627_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_6 _10863_ (.A(_03615_),
    .X(_03649_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_03649_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_6 _10866_ (.A(_03610_),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(_03650_),
    .A1(_03651_),
    .S(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_03649_),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_03616_),
    .X(_03655_));
 sky130_fd_sc_hd__buf_6 _10870_ (.A(_03635_),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(_03654_),
    .A1(_03655_),
    .S(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(_03653_),
    .A1(_03657_),
    .S(_03607_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_4 _10873_ (.A(_03610_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_4 _10874_ (.A(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_4 _10875_ (.A(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__buf_6 _10876_ (.A(_03614_),
    .X(_03662_));
 sky130_fd_sc_hd__buf_4 _10877_ (.A(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__buf_4 _10878_ (.A(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__buf_4 _10880_ (.A(_03635_),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_03663_),
    .X(_03667_));
 sky130_fd_sc_hd__or2_1 _10882_ (.A(_03666_),
    .B(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__buf_4 _10883_ (.A(_03634_),
    .X(_03669_));
 sky130_fd_sc_hd__buf_4 _10884_ (.A(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__buf_4 _10885_ (.A(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__o211a_1 _10886_ (.A1(_03661_),
    .A2(_03665_),
    .B1(_03668_),
    .C1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__buf_6 _10887_ (.A(_03606_),
    .X(_03673_));
 sky130_fd_sc_hd__buf_6 _10888_ (.A(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_03663_),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_03663_),
    .X(_03676_));
 sky130_fd_sc_hd__buf_6 _10891_ (.A(_03635_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _10892_ (.A0(_03675_),
    .A1(_03676_),
    .S(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__buf_6 _10893_ (.A(_03624_),
    .X(_03679_));
 sky130_fd_sc_hd__a21o_1 _10894_ (.A1(_03674_),
    .A2(_03678_),
    .B1(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__inv_2 _10895_ (.A(_03589_),
    .Y(_03681_));
 sky130_fd_sc_hd__nor2_1 _10896_ (.A(_03681_),
    .B(_03597_),
    .Y(_03682_));
 sky130_fd_sc_hd__xnor2_2 _10897_ (.A(_03596_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__or2_4 _10898_ (.A(_03603_),
    .B(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__buf_6 _10899_ (.A(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__o221a_1 _10900_ (.A1(_03648_),
    .A2(_03658_),
    .B1(_03672_),
    .B2(_03680_),
    .C1(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__nor2_4 _10901_ (.A(_03603_),
    .B(_03683_),
    .Y(_03687_));
 sky130_fd_sc_hd__buf_6 _10902_ (.A(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__buf_6 _10903_ (.A(_03669_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_8 _10904_ (.A(_03615_),
    .X(_03690_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _10906_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_03649_),
    .X(_03692_));
 sky130_fd_sc_hd__buf_6 _10907_ (.A(_03635_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _10908_ (.A0(_03691_),
    .A1(_03692_),
    .S(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_03649_),
    .X(_03695_));
 sky130_fd_sc_hd__buf_4 _10910_ (.A(_03556_),
    .X(_03696_));
 sky130_fd_sc_hd__buf_4 _10911_ (.A(_03613_),
    .X(_03697_));
 sky130_fd_sc_hd__and3_1 _10912_ (.A(\rbzero.tex_r0[19] ),
    .B(_03696_),
    .C(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__buf_6 _10913_ (.A(_03614_),
    .X(_03699_));
 sky130_fd_sc_hd__buf_4 _10914_ (.A(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__a21o_1 _10915_ (.A1(\rbzero.tex_r0[18] ),
    .A2(_03700_),
    .B1(_03659_),
    .X(_03701_));
 sky130_fd_sc_hd__buf_4 _10916_ (.A(_03606_),
    .X(_03702_));
 sky130_fd_sc_hd__o221a_1 _10917_ (.A1(_03677_),
    .A2(_03695_),
    .B1(_03698_),
    .B2(_03701_),
    .C1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__buf_4 _10918_ (.A(_03627_),
    .X(_03704_));
 sky130_fd_sc_hd__a211o_1 _10919_ (.A1(_03689_),
    .A2(_03694_),
    .B1(_03703_),
    .C1(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_03690_),
    .X(_03706_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_03649_),
    .X(_03707_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(_03706_),
    .A1(_03707_),
    .S(_03693_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_4 _10923_ (.A(_03662_),
    .X(_03709_));
 sky130_fd_sc_hd__and2_1 _10924_ (.A(\rbzero.tex_r0[30] ),
    .B(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__a31o_1 _10925_ (.A1(\rbzero.tex_r0[31] ),
    .A2(_03696_),
    .A3(_03697_),
    .B1(_03659_),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_03690_),
    .X(_03712_));
 sky130_fd_sc_hd__o221a_1 _10927_ (.A1(_03710_),
    .A2(_03711_),
    .B1(_03712_),
    .B2(_03666_),
    .C1(_03670_),
    .X(_03713_));
 sky130_fd_sc_hd__a211o_1 _10928_ (.A1(_03674_),
    .A2(_03708_),
    .B1(_03713_),
    .C1(_03679_),
    .X(_03714_));
 sky130_fd_sc_hd__nor3_1 _10929_ (.A(_03583_),
    .B(_03582_),
    .C(_03598_),
    .Y(_03715_));
 sky130_fd_sc_hd__o21a_1 _10930_ (.A1(_03583_),
    .A2(_03582_),
    .B1(_03598_),
    .X(_03716_));
 sky130_fd_sc_hd__or3_1 _10931_ (.A(_03603_),
    .B(_03715_),
    .C(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__buf_6 _10932_ (.A(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__inv_4 _10933_ (.A(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__a31o_1 _10934_ (.A1(_03688_),
    .A2(_03705_),
    .A3(_03714_),
    .B1(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__buf_6 _10935_ (.A(_03624_),
    .X(_03721_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_03664_),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_03690_),
    .X(_03723_));
 sky130_fd_sc_hd__or2_1 _10938_ (.A(_03677_),
    .B(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__o211a_1 _10939_ (.A1(_03661_),
    .A2(_03722_),
    .B1(_03724_),
    .C1(_03689_),
    .X(_03725_));
 sky130_fd_sc_hd__buf_4 _10940_ (.A(_03666_),
    .X(_03726_));
 sky130_fd_sc_hd__buf_4 _10941_ (.A(_03649_),
    .X(_03727_));
 sky130_fd_sc_hd__mux2_1 _10942_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__buf_4 _10943_ (.A(_03696_),
    .X(_03729_));
 sky130_fd_sc_hd__buf_4 _10944_ (.A(_03697_),
    .X(_03730_));
 sky130_fd_sc_hd__and3_1 _10945_ (.A(\rbzero.tex_r0[43] ),
    .B(_03729_),
    .C(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__buf_4 _10946_ (.A(_03662_),
    .X(_03732_));
 sky130_fd_sc_hd__clkbuf_4 _10947_ (.A(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__a21o_1 _10948_ (.A1(\rbzero.tex_r0[42] ),
    .A2(_03733_),
    .B1(_03612_),
    .X(_03734_));
 sky130_fd_sc_hd__o221a_1 _10949_ (.A1(_03726_),
    .A2(_03728_),
    .B1(_03731_),
    .B2(_03734_),
    .C1(_03674_),
    .X(_03735_));
 sky130_fd_sc_hd__mux2_1 _10950_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_03663_),
    .X(_03736_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_03663_),
    .X(_03737_));
 sky130_fd_sc_hd__mux2_1 _10952_ (.A0(_03736_),
    .A1(_03737_),
    .S(_03677_),
    .X(_03738_));
 sky130_fd_sc_hd__buf_6 _10953_ (.A(_03635_),
    .X(_03739_));
 sky130_fd_sc_hd__buf_6 _10954_ (.A(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_03709_),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_03662_),
    .X(_03742_));
 sky130_fd_sc_hd__or2_1 _10957_ (.A(_03611_),
    .B(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__o211a_1 _10958_ (.A1(_03740_),
    .A2(_03741_),
    .B1(_03743_),
    .C1(_03670_),
    .X(_03744_));
 sky130_fd_sc_hd__a211o_1 _10959_ (.A1(_03674_),
    .A2(_03738_),
    .B1(_03744_),
    .C1(_03704_),
    .X(_03745_));
 sky130_fd_sc_hd__o311a_1 _10960_ (.A1(_03721_),
    .A2(_03725_),
    .A3(_03735_),
    .B1(_03685_),
    .C1(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_03663_),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_03690_),
    .X(_03748_));
 sky130_fd_sc_hd__mux2_1 _10963_ (.A0(_03747_),
    .A1(_03748_),
    .S(_03693_),
    .X(_03749_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_03663_),
    .X(_03750_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_03662_),
    .X(_03751_));
 sky130_fd_sc_hd__or2_1 _10966_ (.A(_03659_),
    .B(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__o211a_1 _10967_ (.A1(_03666_),
    .A2(_03750_),
    .B1(_03752_),
    .C1(_03670_),
    .X(_03753_));
 sky130_fd_sc_hd__a211o_1 _10968_ (.A1(_03674_),
    .A2(_03749_),
    .B1(_03753_),
    .C1(_03679_),
    .X(_03754_));
 sky130_fd_sc_hd__mux2_1 _10969_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_03690_),
    .X(_03755_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_03690_),
    .X(_03756_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(_03755_),
    .A1(_03756_),
    .S(_03693_),
    .X(_03757_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_03690_),
    .X(_03758_));
 sky130_fd_sc_hd__and3_1 _10973_ (.A(\rbzero.tex_r0[51] ),
    .B(_03696_),
    .C(_03697_),
    .X(_03759_));
 sky130_fd_sc_hd__a21o_1 _10974_ (.A1(\rbzero.tex_r0[50] ),
    .A2(_03700_),
    .B1(_03659_),
    .X(_03760_));
 sky130_fd_sc_hd__o221a_1 _10975_ (.A1(_03666_),
    .A2(_03758_),
    .B1(_03759_),
    .B2(_03760_),
    .C1(_03702_),
    .X(_03761_));
 sky130_fd_sc_hd__a211o_1 _10976_ (.A1(_03689_),
    .A2(_03757_),
    .B1(_03761_),
    .C1(_03704_),
    .X(_03762_));
 sky130_fd_sc_hd__a31o_1 _10977_ (.A1(_03688_),
    .A2(_03754_),
    .A3(_03762_),
    .B1(_03718_),
    .X(_03763_));
 sky130_fd_sc_hd__inv_2 _10978_ (.A(net41),
    .Y(_03764_));
 sky130_fd_sc_hd__o221a_1 _10979_ (.A1(_03686_),
    .A2(_03720_),
    .B1(_03746_),
    .B2(_03763_),
    .C1(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__a31o_1 _10980_ (.A1(_03537_),
    .A2(_03541_),
    .A3(_03647_),
    .B1(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__buf_2 _10981_ (.A(_03620_),
    .X(_03767_));
 sky130_fd_sc_hd__clkbuf_4 _10982_ (.A(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__or4_1 _10983_ (.A(_03636_),
    .B(_03719_),
    .C(_03687_),
    .D(_03535_),
    .X(_03769_));
 sky130_fd_sc_hd__inv_2 _10984_ (.A(\rbzero.row_render.size[2] ),
    .Y(_03770_));
 sky130_fd_sc_hd__nor2_1 _10985_ (.A(\rbzero.row_render.size[1] ),
    .B(\rbzero.row_render.size[0] ),
    .Y(_03771_));
 sky130_fd_sc_hd__nand2_1 _10986_ (.A(_03770_),
    .B(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__or2_1 _10987_ (.A(\rbzero.row_render.size[3] ),
    .B(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__or3_1 _10988_ (.A(\rbzero.row_render.size[5] ),
    .B(\rbzero.row_render.size[4] ),
    .C(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__and2_1 _10989_ (.A(\rbzero.row_render.size[6] ),
    .B(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__o21a_1 _10990_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_03775_),
    .B1(\rbzero.row_render.size[8] ),
    .X(_03776_));
 sky130_fd_sc_hd__xnor2_1 _10991_ (.A(\rbzero.row_render.size[7] ),
    .B(\rbzero.row_render.size[6] ),
    .Y(_03777_));
 sky130_fd_sc_hd__a21o_1 _10992_ (.A1(\rbzero.row_render.size[7] ),
    .A2(\rbzero.row_render.size[6] ),
    .B1(\rbzero.row_render.size[8] ),
    .X(_03778_));
 sky130_fd_sc_hd__nand3_1 _10993_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(\rbzero.row_render.size[6] ),
    .Y(_03779_));
 sky130_fd_sc_hd__and2_1 _10994_ (.A(_03778_),
    .B(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__inv_2 _10995_ (.A(\gpout0.hpos[5] ),
    .Y(_03781_));
 sky130_fd_sc_hd__buf_4 _10996_ (.A(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__clkinv_2 _10997_ (.A(\gpout0.hpos[2] ),
    .Y(_03783_));
 sky130_fd_sc_hd__a211o_1 _10998_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_03499_),
    .B1(_03500_),
    .C1(\rbzero.row_render.size[0] ),
    .X(_03784_));
 sky130_fd_sc_hd__o221a_1 _10999_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_03783_),
    .B1(_03499_),
    .B2(\rbzero.row_render.size[1] ),
    .C1(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__a221o_1 _11000_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_03783_),
    .B1(_03462_),
    .B2(\rbzero.row_render.size[3] ),
    .C1(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__o221a_1 _11001_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_03462_),
    .B1(_03463_),
    .B2(\rbzero.row_render.size[4] ),
    .C1(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__a221o_1 _11002_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_03463_),
    .B1(_03782_),
    .B2(\rbzero.row_render.size[5] ),
    .C1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__o2bb2a_1 _11003_ (.A1_N(\rbzero.row_render.size[6] ),
    .A2_N(_03466_),
    .B1(_03781_),
    .B2(\rbzero.row_render.size[5] ),
    .X(_03789_));
 sky130_fd_sc_hd__o22ai_1 _11004_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_03466_),
    .B1(_03777_),
    .B2(_02900_),
    .Y(_03790_));
 sky130_fd_sc_hd__a21oi_1 _11005_ (.A1(_03788_),
    .A2(_03789_),
    .B1(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__a221o_1 _11006_ (.A1(_02900_),
    .A2(_03777_),
    .B1(_03780_),
    .B2(_02902_),
    .C1(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__nor2_1 _11007_ (.A(\rbzero.row_render.size[9] ),
    .B(_03778_),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_1 _11008_ (.A(\rbzero.row_render.size[9] ),
    .B(_03778_),
    .Y(_03794_));
 sky130_fd_sc_hd__o221a_1 _11009_ (.A1(_02902_),
    .A2(_03780_),
    .B1(_03793_),
    .B2(\gpout0.hpos[9] ),
    .C1(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__nor3_1 _11010_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(_03775_),
    .Y(_03796_));
 sky130_fd_sc_hd__nor2_1 _11011_ (.A(_03776_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__xnor2_1 _11012_ (.A(\rbzero.row_render.size[7] ),
    .B(_03775_),
    .Y(_03798_));
 sky130_fd_sc_hd__a22o_1 _11013_ (.A1(_02900_),
    .A2(_03798_),
    .B1(_03797_),
    .B2(_02902_),
    .X(_03799_));
 sky130_fd_sc_hd__nor2_1 _11014_ (.A(\rbzero.row_render.size[6] ),
    .B(_03774_),
    .Y(_03800_));
 sky130_fd_sc_hd__nor2_1 _11015_ (.A(_03775_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__o21ai_1 _11016_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_03773_),
    .B1(\rbzero.row_render.size[5] ),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _11017_ (.A(_03774_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__xnor2_1 _11018_ (.A(\rbzero.row_render.size[4] ),
    .B(_03773_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand2_1 _11019_ (.A(\rbzero.row_render.size[3] ),
    .B(_03772_),
    .Y(_03805_));
 sky130_fd_sc_hd__nand2_1 _11020_ (.A(_03773_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__or2_1 _11021_ (.A(_03770_),
    .B(_03771_),
    .X(_03807_));
 sky130_fd_sc_hd__nand2_1 _11022_ (.A(_03772_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__or2_1 _11023_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .X(_03809_));
 sky130_fd_sc_hd__or2_1 _11024_ (.A(\rbzero.row_render.size[0] ),
    .B(_03527_),
    .X(_03810_));
 sky130_fd_sc_hd__a31o_1 _11025_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_03809_),
    .A3(_03810_),
    .B1(_03771_),
    .X(_03811_));
 sky130_fd_sc_hd__a211o_1 _11026_ (.A1(\rbzero.row_render.size[2] ),
    .A2(\gpout0.hpos[2] ),
    .B1(_03501_),
    .C1(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__o221a_1 _11027_ (.A1(\gpout0.hpos[3] ),
    .A2(_03806_),
    .B1(_03808_),
    .B2(_03526_),
    .C1(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__a221o_1 _11028_ (.A1(_03523_),
    .A2(_03806_),
    .B1(_03804_),
    .B2(\gpout0.hpos[4] ),
    .C1(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__o221a_1 _11029_ (.A1(\gpout0.hpos[4] ),
    .A2(_03804_),
    .B1(_03803_),
    .B2(_03460_),
    .C1(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__a221o_1 _11030_ (.A1(_03460_),
    .A2(_03803_),
    .B1(_03801_),
    .B2(_03466_),
    .C1(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__o221a_1 _11031_ (.A1(_03466_),
    .A2(_03801_),
    .B1(_03798_),
    .B2(_02900_),
    .C1(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__o221a_1 _11032_ (.A1(_02902_),
    .A2(_03797_),
    .B1(_03799_),
    .B2(_03817_),
    .C1(_02903_),
    .X(_03818_));
 sky130_fd_sc_hd__nor2_1 _11033_ (.A(_02903_),
    .B(_03793_),
    .Y(_03819_));
 sky130_fd_sc_hd__o2bb2a_1 _11034_ (.A1_N(_03792_),
    .A2_N(_03795_),
    .B1(_03818_),
    .B2(_03819_),
    .X(_03820_));
 sky130_fd_sc_hd__or4_4 _11035_ (.A(\rbzero.row_render.size[10] ),
    .B(\rbzero.row_render.size[9] ),
    .C(_03776_),
    .D(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__o31a_1 _11036_ (.A1(_03726_),
    .A2(_03768_),
    .A3(_03769_),
    .B1(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__buf_6 _11037_ (.A(_03610_),
    .X(_03823_));
 sky130_fd_sc_hd__o211a_1 _11038_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_03610_),
    .B1(_03662_),
    .C1(\rbzero.floor_leak[0] ),
    .X(_03824_));
 sky130_fd_sc_hd__a221o_1 _11039_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_03606_),
    .B1(_03823_),
    .B2(\rbzero.floor_leak[1] ),
    .C1(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__o221a_1 _11040_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_03624_),
    .B1(_03673_),
    .B2(\rbzero.floor_leak[2] ),
    .C1(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__a221o_1 _11041_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_03624_),
    .B1(_03684_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__o221a_1 _11042_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_03718_),
    .B1(_03685_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__a21oi_1 _11043_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_03718_),
    .B1(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__o21a_2 _11044_ (.A1(\rbzero.row_render.vinf ),
    .A2(_03822_),
    .B1(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(_03536_),
    .A1(_03766_),
    .S(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__xor2_1 _11046_ (.A(\gpout0.vpos[5] ),
    .B(\rbzero.debug_overlay.playerY[2] ),
    .X(_03832_));
 sky130_fd_sc_hd__xor2_1 _11047_ (.A(_03517_),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .X(_03833_));
 sky130_fd_sc_hd__buf_4 _11048_ (.A(\gpout0.vpos[4] ),
    .X(_03834_));
 sky130_fd_sc_hd__xnor2_1 _11049_ (.A(_03834_),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .Y(_03835_));
 sky130_fd_sc_hd__o221a_1 _11050_ (.A1(\gpout0.vpos[6] ),
    .A2(_03347_),
    .B1(\rbzero.debug_overlay.playerX[0] ),
    .B2(_03462_),
    .C1(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__or3b_1 _11051_ (.A(_03832_),
    .B(_03833_),
    .C_N(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__buf_4 _11052_ (.A(_03466_),
    .X(_03838_));
 sky130_fd_sc_hd__inv_2 _11053_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .Y(_03839_));
 sky130_fd_sc_hd__clkinv_2 _11054_ (.A(\gpout0.vpos[7] ),
    .Y(_03840_));
 sky130_fd_sc_hd__a22o_1 _11055_ (.A1(_03840_),
    .A2(\rbzero.debug_overlay.playerY[4] ),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .B2(_03782_),
    .X(_03841_));
 sky130_fd_sc_hd__a221o_1 _11056_ (.A1(\gpout0.vpos[6] ),
    .A2(_03347_),
    .B1(_03363_),
    .B2(_03460_),
    .C1(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__a221o_1 _11057_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03463_),
    .B1(_03838_),
    .B2(_03839_),
    .C1(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__a221o_1 _11058_ (.A1(_03515_),
    .A2(_03344_),
    .B1(_03342_),
    .B2(_03524_),
    .C1(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__xor2_1 _11059_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_02901_),
    .X(_03845_));
 sky130_fd_sc_hd__a221o_1 _11060_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03462_),
    .B1(_03474_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .C1(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__or3_2 _11061_ (.A(_03837_),
    .B(_03844_),
    .C(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__and3_1 _11062_ (.A(_03518_),
    .B(_03529_),
    .C(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__inv_2 _11063_ (.A(\gpout0.vpos[5] ),
    .Y(_03849_));
 sky130_fd_sc_hd__xnor2_1 _11064_ (.A(_03834_),
    .B(\rbzero.map_overlay.i_mapdy[1] ),
    .Y(_03850_));
 sky130_fd_sc_hd__o221a_1 _11065_ (.A1(\gpout0.vpos[6] ),
    .A2(_03447_),
    .B1(\rbzero.map_overlay.i_mapdy[2] ),
    .B2(_03849_),
    .C1(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__buf_4 _11066_ (.A(_03849_),
    .X(_03852_));
 sky130_fd_sc_hd__o2bb2a_1 _11067_ (.A1_N(\rbzero.map_overlay.i_mapdy[2] ),
    .A2_N(_03852_),
    .B1(\gpout0.vpos[7] ),
    .B2(_03451_),
    .X(_03853_));
 sky130_fd_sc_hd__inv_2 _11068_ (.A(\gpout0.vpos[3] ),
    .Y(_03854_));
 sky130_fd_sc_hd__or4_1 _11069_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_overlay.i_mapdy[2] ),
    .C(\rbzero.map_overlay.i_mapdy[1] ),
    .D(\rbzero.map_overlay.i_mapdy[0] ),
    .X(_03855_));
 sky130_fd_sc_hd__o21a_1 _11070_ (.A1(\rbzero.map_overlay.i_mapdy[5] ),
    .A2(_03855_),
    .B1(_03840_),
    .X(_03856_));
 sky130_fd_sc_hd__inv_2 _11071_ (.A(\gpout0.vpos[6] ),
    .Y(_03857_));
 sky130_fd_sc_hd__o2bb2a_1 _11072_ (.A1_N(_03854_),
    .A2_N(\rbzero.map_overlay.i_mapdy[0] ),
    .B1(\rbzero.map_overlay.i_mapdy[3] ),
    .B2(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__o221a_1 _11073_ (.A1(_03854_),
    .A2(\rbzero.map_overlay.i_mapdy[0] ),
    .B1(_03856_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__and3_1 _11074_ (.A(_03851_),
    .B(_03853_),
    .C(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__xor2_1 _11075_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_03838_),
    .X(_03861_));
 sky130_fd_sc_hd__xor2_1 _11076_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_03460_),
    .X(_03862_));
 sky130_fd_sc_hd__a221o_1 _11077_ (.A1(_03425_),
    .A2(_03523_),
    .B1(_03464_),
    .B2(\rbzero.map_overlay.i_mapdx[1] ),
    .C1(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__o21a_1 _11078_ (.A1(\rbzero.map_overlay.i_mapdx[5] ),
    .A2(_03421_),
    .B1(_03420_),
    .X(_03864_));
 sky130_fd_sc_hd__clkinv_4 _11079_ (.A(_02900_),
    .Y(_03865_));
 sky130_fd_sc_hd__o22a_1 _11080_ (.A1(\rbzero.map_overlay.i_mapdx[1] ),
    .A2(_03463_),
    .B1(_03865_),
    .B2(\rbzero.map_overlay.i_mapdx[4] ),
    .X(_03866_));
 sky130_fd_sc_hd__o221a_1 _11081_ (.A1(_03425_),
    .A2(_03523_),
    .B1(_02900_),
    .B2(_03864_),
    .C1(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__or3b_2 _11082_ (.A(_03861_),
    .B(_03863_),
    .C_N(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__xor2_1 _11083_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_02900_),
    .X(_03869_));
 sky130_fd_sc_hd__a221o_1 _11084_ (.A1(\rbzero.map_overlay.i_otherx[0] ),
    .A2(_03462_),
    .B1(_03474_),
    .B2(\rbzero.map_overlay.i_otherx[3] ),
    .C1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__inv_2 _11085_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .Y(_03871_));
 sky130_fd_sc_hd__inv_2 _11086_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .Y(_03872_));
 sky130_fd_sc_hd__inv_2 _11087_ (.A(\rbzero.map_overlay.i_othery[3] ),
    .Y(_03873_));
 sky130_fd_sc_hd__inv_2 _11088_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .Y(_03874_));
 sky130_fd_sc_hd__a22o_1 _11089_ (.A1(_03840_),
    .A2(\rbzero.map_overlay.i_othery[4] ),
    .B1(\rbzero.map_overlay.i_otherx[2] ),
    .B2(_03781_),
    .X(_03875_));
 sky130_fd_sc_hd__a221o_1 _11090_ (.A1(\gpout0.vpos[6] ),
    .A2(_03873_),
    .B1(_03874_),
    .B2(_03460_),
    .C1(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__a221o_1 _11091_ (.A1(\rbzero.map_overlay.i_otherx[1] ),
    .A2(_03463_),
    .B1(_03466_),
    .B2(_03872_),
    .C1(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__a221o_1 _11092_ (.A1(\gpout0.vpos[7] ),
    .A2(_03871_),
    .B1(_03430_),
    .B2(_03524_),
    .C1(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_1 _11093_ (.A(_03517_),
    .B(\rbzero.map_overlay.i_othery[0] ),
    .Y(_03879_));
 sky130_fd_sc_hd__or2_1 _11094_ (.A(\gpout0.vpos[3] ),
    .B(\rbzero.map_overlay.i_othery[0] ),
    .X(_03880_));
 sky130_fd_sc_hd__inv_2 _11095_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .Y(_03881_));
 sky130_fd_sc_hd__xor2_1 _11096_ (.A(\gpout0.vpos[4] ),
    .B(\rbzero.map_overlay.i_othery[1] ),
    .X(_03882_));
 sky130_fd_sc_hd__a221o_1 _11097_ (.A1(_03857_),
    .A2(\rbzero.map_overlay.i_othery[3] ),
    .B1(_03881_),
    .B2(_03523_),
    .C1(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__xor2_1 _11098_ (.A(\gpout0.vpos[5] ),
    .B(\rbzero.map_overlay.i_othery[2] ),
    .X(_03884_));
 sky130_fd_sc_hd__a211o_1 _11099_ (.A1(_03879_),
    .A2(_03880_),
    .B1(_03883_),
    .C1(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__or3_1 _11100_ (.A(_03870_),
    .B(_03878_),
    .C(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__a21bo_1 _11101_ (.A1(_03860_),
    .A2(_03868_),
    .B1_N(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__xnor2_1 _11102_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(\gpout0.hpos[0] ),
    .Y(_03888_));
 sky130_fd_sc_hd__xnor2_1 _11103_ (.A(\gpout0.vpos[1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .Y(_03889_));
 sky130_fd_sc_hd__inv_2 _11104_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .Y(_03890_));
 sky130_fd_sc_hd__xnor2_1 _11105_ (.A(\gpout0.vpos[2] ),
    .B(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_03891_));
 sky130_fd_sc_hd__o221a_1 _11106_ (.A1(\gpout0.vpos[0] ),
    .A2(_03890_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .B2(_03783_),
    .C1(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__xor2_1 _11107_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_03527_),
    .X(_03893_));
 sky130_fd_sc_hd__a221o_1 _11108_ (.A1(\gpout0.vpos[0] ),
    .A2(_03890_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .B2(_03783_),
    .C1(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__nor2_1 _11109_ (.A(_03847_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__or3_2 _11110_ (.A(_03530_),
    .B(_03532_),
    .C(_03533_),
    .X(_03896_));
 sky130_fd_sc_hd__a41o_1 _11111_ (.A1(_03888_),
    .A2(_03889_),
    .A3(_03892_),
    .A4(_03895_),
    .B1(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__a21o_1 _11112_ (.A1(_03848_),
    .A2(_03887_),
    .B1(_03897_),
    .X(_03898_));
 sky130_fd_sc_hd__o21a_1 _11113_ (.A1(_03534_),
    .A2(_03831_),
    .B1(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__or2_2 _11114_ (.A(\gpout0.vpos[4] ),
    .B(\gpout0.vpos[3] ),
    .X(_03900_));
 sky130_fd_sc_hd__nand2_4 _11115_ (.A(_03834_),
    .B(\gpout0.vpos[3] ),
    .Y(_03901_));
 sky130_fd_sc_hd__buf_4 _11116_ (.A(\gpout0.vpos[5] ),
    .X(_03902_));
 sky130_fd_sc_hd__nand2_1 _11117_ (.A(_03902_),
    .B(_03834_),
    .Y(_03903_));
 sky130_fd_sc_hd__nand2_1 _11118_ (.A(_03502_),
    .B(_03518_),
    .Y(_03904_));
 sky130_fd_sc_hd__a41o_1 _11119_ (.A1(_03519_),
    .A2(_03900_),
    .A3(_03901_),
    .A4(_03903_),
    .B1(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__clkbuf_4 _11120_ (.A(\gpout0.vpos[8] ),
    .X(_03906_));
 sky130_fd_sc_hd__nand2_1 _11121_ (.A(\gpout0.vpos[7] ),
    .B(\gpout0.vpos[6] ),
    .Y(_03907_));
 sky130_fd_sc_hd__nor2_1 _11122_ (.A(_03849_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__clkbuf_4 _11123_ (.A(\gpout0.vpos[9] ),
    .X(_03909_));
 sky130_fd_sc_hd__a21o_4 _11124_ (.A1(_03906_),
    .A2(_03908_),
    .B1(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__clkbuf_8 _11125_ (.A(_03504_),
    .X(_03911_));
 sky130_fd_sc_hd__a211oi_4 _11126_ (.A1(_03522_),
    .A2(_03905_),
    .B1(_03910_),
    .C1(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__o21ai_4 _11127_ (.A1(_03522_),
    .A2(_03899_),
    .B1(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__inv_2 _11128_ (.A(_03913_),
    .Y(net66));
 sky130_fd_sc_hd__or2b_1 _11129_ (.A(\rbzero.color_floor[1] ),
    .B_N(_03535_),
    .X(_03914_));
 sky130_fd_sc_hd__o21ai_1 _11130_ (.A1(\rbzero.color_sky[1] ),
    .A2(_03535_),
    .B1(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__or2_1 _11131_ (.A(\rbzero.tex_r1[54] ),
    .B(_03767_),
    .X(_03916_));
 sky130_fd_sc_hd__clkbuf_8 _11132_ (.A(_03693_),
    .X(_03917_));
 sky130_fd_sc_hd__o211a_1 _11133_ (.A1(\rbzero.tex_r1[55] ),
    .A2(_03618_),
    .B1(_03916_),
    .C1(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__clkbuf_4 _11134_ (.A(_03823_),
    .X(_03919_));
 sky130_fd_sc_hd__clkbuf_4 _11135_ (.A(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__a31o_1 _11136_ (.A1(\rbzero.tex_r1[53] ),
    .A2(_03652_),
    .A3(_03767_),
    .B1(_03673_),
    .X(_03921_));
 sky130_fd_sc_hd__a31o_1 _11137_ (.A1(\rbzero.tex_r1[52] ),
    .A2(_03920_),
    .A3(_03618_),
    .B1(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__or2_1 _11138_ (.A(\rbzero.tex_r1[50] ),
    .B(_03767_),
    .X(_03923_));
 sky130_fd_sc_hd__o211a_1 _11139_ (.A1(\rbzero.tex_r1[51] ),
    .A2(_03618_),
    .B1(_03923_),
    .C1(_03917_),
    .X(_03924_));
 sky130_fd_sc_hd__clkbuf_4 _11140_ (.A(_03733_),
    .X(_03925_));
 sky130_fd_sc_hd__clkbuf_4 _11141_ (.A(_03620_),
    .X(_03926_));
 sky130_fd_sc_hd__a31o_1 _11142_ (.A1(\rbzero.tex_r1[49] ),
    .A2(_03919_),
    .A3(_03926_),
    .B1(_03669_),
    .X(_03927_));
 sky130_fd_sc_hd__a31o_1 _11143_ (.A1(\rbzero.tex_r1[48] ),
    .A2(_03920_),
    .A3(_03925_),
    .B1(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__o221a_1 _11144_ (.A1(_03918_),
    .A2(_03922_),
    .B1(_03924_),
    .B2(_03928_),
    .C1(_03721_),
    .X(_03929_));
 sky130_fd_sc_hd__or2_1 _11145_ (.A(\rbzero.tex_r1[62] ),
    .B(_03767_),
    .X(_03930_));
 sky130_fd_sc_hd__o211a_1 _11146_ (.A1(\rbzero.tex_r1[63] ),
    .A2(_03925_),
    .B1(_03930_),
    .C1(_03917_),
    .X(_03931_));
 sky130_fd_sc_hd__a31o_1 _11147_ (.A1(\rbzero.tex_r1[61] ),
    .A2(_03919_),
    .A3(_03926_),
    .B1(_03673_),
    .X(_03932_));
 sky130_fd_sc_hd__a31o_1 _11148_ (.A1(\rbzero.tex_r1[60] ),
    .A2(_03920_),
    .A3(_03925_),
    .B1(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__or2_1 _11149_ (.A(\rbzero.tex_r1[58] ),
    .B(_03926_),
    .X(_03934_));
 sky130_fd_sc_hd__o211a_1 _11150_ (.A1(\rbzero.tex_r1[59] ),
    .A2(_03925_),
    .B1(_03934_),
    .C1(_03726_),
    .X(_03935_));
 sky130_fd_sc_hd__buf_4 _11151_ (.A(_03733_),
    .X(_03936_));
 sky130_fd_sc_hd__a31o_1 _11152_ (.A1(\rbzero.tex_r1[57] ),
    .A2(_03919_),
    .A3(_03768_),
    .B1(_03670_),
    .X(_03937_));
 sky130_fd_sc_hd__a31o_1 _11153_ (.A1(\rbzero.tex_r1[56] ),
    .A2(_03661_),
    .A3(_03936_),
    .B1(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__o221a_1 _11154_ (.A1(_03931_),
    .A2(_03933_),
    .B1(_03935_),
    .B2(_03938_),
    .C1(_03648_),
    .X(_03939_));
 sky130_fd_sc_hd__or2_1 _11155_ (.A(\rbzero.tex_r1[46] ),
    .B(_03620_),
    .X(_03940_));
 sky130_fd_sc_hd__o211a_1 _11156_ (.A1(\rbzero.tex_r1[47] ),
    .A2(_03664_),
    .B1(_03940_),
    .C1(_03677_),
    .X(_03941_));
 sky130_fd_sc_hd__a31o_1 _11157_ (.A1(\rbzero.tex_r1[45] ),
    .A2(_03919_),
    .A3(_03926_),
    .B1(_03673_),
    .X(_03942_));
 sky130_fd_sc_hd__a311o_1 _11158_ (.A1(\rbzero.tex_r1[44] ),
    .A2(_03920_),
    .A3(_03925_),
    .B1(_03941_),
    .C1(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__or2_1 _11159_ (.A(\rbzero.tex_r1[42] ),
    .B(_03620_),
    .X(_03944_));
 sky130_fd_sc_hd__o211a_1 _11160_ (.A1(\rbzero.tex_r1[43] ),
    .A2(_03664_),
    .B1(_03944_),
    .C1(_03677_),
    .X(_03945_));
 sky130_fd_sc_hd__a31o_1 _11161_ (.A1(\rbzero.tex_r1[41] ),
    .A2(_03919_),
    .A3(_03926_),
    .B1(_03669_),
    .X(_03946_));
 sky130_fd_sc_hd__a311o_1 _11162_ (.A1(\rbzero.tex_r1[40] ),
    .A2(_03920_),
    .A3(_03618_),
    .B1(_03945_),
    .C1(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__or2_1 _11163_ (.A(\rbzero.tex_r1[38] ),
    .B(_03767_),
    .X(_03948_));
 sky130_fd_sc_hd__o211a_1 _11164_ (.A1(\rbzero.tex_r1[39] ),
    .A2(_03733_),
    .B1(_03948_),
    .C1(_03666_),
    .X(_03949_));
 sky130_fd_sc_hd__a31o_1 _11165_ (.A1(\rbzero.tex_r1[37] ),
    .A2(_03659_),
    .A3(_03767_),
    .B1(_03606_),
    .X(_03950_));
 sky130_fd_sc_hd__a31o_1 _11166_ (.A1(\rbzero.tex_r1[36] ),
    .A2(_03919_),
    .A3(_03733_),
    .B1(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__or2_1 _11167_ (.A(\rbzero.tex_r1[34] ),
    .B(_03767_),
    .X(_03952_));
 sky130_fd_sc_hd__o211a_1 _11168_ (.A1(\rbzero.tex_r1[35] ),
    .A2(_03733_),
    .B1(_03952_),
    .C1(_03666_),
    .X(_03953_));
 sky130_fd_sc_hd__a31o_1 _11169_ (.A1(\rbzero.tex_r1[33] ),
    .A2(_03659_),
    .A3(_03767_),
    .B1(_03634_),
    .X(_03954_));
 sky130_fd_sc_hd__a31o_1 _11170_ (.A1(\rbzero.tex_r1[32] ),
    .A2(_03660_),
    .A3(_03733_),
    .B1(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__o221a_1 _11171_ (.A1(_03949_),
    .A2(_03951_),
    .B1(_03953_),
    .B2(_03955_),
    .C1(_03679_),
    .X(_03956_));
 sky130_fd_sc_hd__a311o_1 _11172_ (.A1(_03648_),
    .A2(_03943_),
    .A3(_03947_),
    .B1(_03687_),
    .C1(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__o311a_1 _11173_ (.A1(_03685_),
    .A2(_03929_),
    .A3(_03939_),
    .B1(_03957_),
    .C1(_03719_),
    .X(_03958_));
 sky130_fd_sc_hd__or2_1 _11174_ (.A(\rbzero.tex_r1[6] ),
    .B(_03926_),
    .X(_03959_));
 sky130_fd_sc_hd__o211a_1 _11175_ (.A1(\rbzero.tex_r1[7] ),
    .A2(_03925_),
    .B1(_03959_),
    .C1(_03726_),
    .X(_03960_));
 sky130_fd_sc_hd__a31o_1 _11176_ (.A1(\rbzero.tex_r1[5] ),
    .A2(_03919_),
    .A3(_03926_),
    .B1(_03673_),
    .X(_03961_));
 sky130_fd_sc_hd__a31o_1 _11177_ (.A1(\rbzero.tex_r1[4] ),
    .A2(_03661_),
    .A3(_03936_),
    .B1(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__or2_1 _11178_ (.A(\rbzero.tex_r1[2] ),
    .B(_03926_),
    .X(_03963_));
 sky130_fd_sc_hd__o211a_1 _11179_ (.A1(\rbzero.tex_r1[3] ),
    .A2(_03936_),
    .B1(_03963_),
    .C1(_03726_),
    .X(_03964_));
 sky130_fd_sc_hd__a31o_1 _11180_ (.A1(\rbzero.tex_r1[1] ),
    .A2(_03660_),
    .A3(_03768_),
    .B1(_03670_),
    .X(_03965_));
 sky130_fd_sc_hd__a31o_1 _11181_ (.A1(\rbzero.tex_r1[0] ),
    .A2(_03661_),
    .A3(_03936_),
    .B1(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__o221a_1 _11182_ (.A1(_03960_),
    .A2(_03962_),
    .B1(_03964_),
    .B2(_03966_),
    .C1(_03721_),
    .X(_03967_));
 sky130_fd_sc_hd__or2_1 _11183_ (.A(\rbzero.tex_r1[14] ),
    .B(_03620_),
    .X(_03968_));
 sky130_fd_sc_hd__o211a_1 _11184_ (.A1(\rbzero.tex_r1[15] ),
    .A2(_03664_),
    .B1(_03968_),
    .C1(_03677_),
    .X(_03969_));
 sky130_fd_sc_hd__a31o_1 _11185_ (.A1(\rbzero.tex_r1[13] ),
    .A2(_03919_),
    .A3(_03768_),
    .B1(_03673_),
    .X(_03970_));
 sky130_fd_sc_hd__a311o_1 _11186_ (.A1(\rbzero.tex_r1[12] ),
    .A2(_03920_),
    .A3(_03925_),
    .B1(_03969_),
    .C1(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__or2_1 _11187_ (.A(\rbzero.tex_r1[10] ),
    .B(_03620_),
    .X(_03972_));
 sky130_fd_sc_hd__o211a_1 _11188_ (.A1(\rbzero.tex_r1[11] ),
    .A2(_03664_),
    .B1(_03972_),
    .C1(_03677_),
    .X(_03973_));
 sky130_fd_sc_hd__a31o_1 _11189_ (.A1(\rbzero.tex_r1[9] ),
    .A2(_03919_),
    .A3(_03926_),
    .B1(_03670_),
    .X(_03974_));
 sky130_fd_sc_hd__a311o_1 _11190_ (.A1(\rbzero.tex_r1[8] ),
    .A2(_03920_),
    .A3(_03925_),
    .B1(_03973_),
    .C1(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__a31o_1 _11191_ (.A1(_03648_),
    .A2(_03971_),
    .A3(_03975_),
    .B1(_03687_),
    .X(_03976_));
 sky130_fd_sc_hd__or2_1 _11192_ (.A(\rbzero.tex_r1[30] ),
    .B(_03926_),
    .X(_03977_));
 sky130_fd_sc_hd__o211a_1 _11193_ (.A1(\rbzero.tex_r1[31] ),
    .A2(_03936_),
    .B1(_03977_),
    .C1(_03726_),
    .X(_03978_));
 sky130_fd_sc_hd__a31o_1 _11194_ (.A1(\rbzero.tex_r1[29] ),
    .A2(_03660_),
    .A3(_03768_),
    .B1(_03702_),
    .X(_03979_));
 sky130_fd_sc_hd__a31o_1 _11195_ (.A1(\rbzero.tex_r1[28] ),
    .A2(_03661_),
    .A3(_03936_),
    .B1(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__or2_1 _11196_ (.A(\rbzero.tex_r1[26] ),
    .B(_03768_),
    .X(_03981_));
 sky130_fd_sc_hd__o211a_1 _11197_ (.A1(\rbzero.tex_r1[27] ),
    .A2(_03936_),
    .B1(_03981_),
    .C1(_03726_),
    .X(_03982_));
 sky130_fd_sc_hd__a31o_1 _11198_ (.A1(\rbzero.tex_r1[25] ),
    .A2(_03660_),
    .A3(_03768_),
    .B1(_03670_),
    .X(_03983_));
 sky130_fd_sc_hd__a31o_1 _11199_ (.A1(\rbzero.tex_r1[24] ),
    .A2(_03661_),
    .A3(_03936_),
    .B1(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__o221a_1 _11200_ (.A1(_03978_),
    .A2(_03980_),
    .B1(_03982_),
    .B2(_03984_),
    .C1(_03648_),
    .X(_03985_));
 sky130_fd_sc_hd__or2_1 _11201_ (.A(\rbzero.tex_r1[22] ),
    .B(_03767_),
    .X(_03986_));
 sky130_fd_sc_hd__o211a_1 _11202_ (.A1(\rbzero.tex_r1[23] ),
    .A2(_03733_),
    .B1(_03986_),
    .C1(_03666_),
    .X(_03987_));
 sky130_fd_sc_hd__a31o_1 _11203_ (.A1(\rbzero.tex_r1[21] ),
    .A2(_03660_),
    .A3(_03768_),
    .B1(_03702_),
    .X(_03988_));
 sky130_fd_sc_hd__a311o_1 _11204_ (.A1(\rbzero.tex_r1[20] ),
    .A2(_03920_),
    .A3(_03936_),
    .B1(_03987_),
    .C1(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__or2_1 _11205_ (.A(\rbzero.tex_r1[18] ),
    .B(_03620_),
    .X(_03990_));
 sky130_fd_sc_hd__o211a_1 _11206_ (.A1(\rbzero.tex_r1[19] ),
    .A2(_03664_),
    .B1(_03990_),
    .C1(_03677_),
    .X(_03991_));
 sky130_fd_sc_hd__a31o_1 _11207_ (.A1(\rbzero.tex_r1[17] ),
    .A2(_03660_),
    .A3(_03768_),
    .B1(_03670_),
    .X(_03992_));
 sky130_fd_sc_hd__a311o_1 _11208_ (.A1(\rbzero.tex_r1[16] ),
    .A2(_03920_),
    .A3(_03925_),
    .B1(_03991_),
    .C1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__a31o_1 _11209_ (.A1(_03721_),
    .A2(_03989_),
    .A3(_03993_),
    .B1(_03685_),
    .X(_03994_));
 sky130_fd_sc_hd__o221a_1 _11210_ (.A1(_03967_),
    .A2(_03976_),
    .B1(_03985_),
    .B2(_03994_),
    .C1(_03718_),
    .X(_03995_));
 sky130_fd_sc_hd__or2_1 _11211_ (.A(_03539_),
    .B(\rbzero.row_render.wall[1] ),
    .X(_03996_));
 sky130_fd_sc_hd__a21oi_1 _11212_ (.A1(\rbzero.row_render.side ),
    .A2(_03631_),
    .B1(\rbzero.row_render.wall[0] ),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_1 _11213_ (.A(\rbzero.row_render.wall[1] ),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__o21a_1 _11214_ (.A1(_03638_),
    .A2(_03643_),
    .B1(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__or2_1 _11215_ (.A(\rbzero.row_render.texu[4] ),
    .B(_03687_),
    .X(_04000_));
 sky130_fd_sc_hd__a21oi_1 _11216_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_03688_),
    .B1(_03996_),
    .Y(_04001_));
 sky130_fd_sc_hd__a221o_1 _11217_ (.A1(_03996_),
    .A2(_03999_),
    .B1(_04000_),
    .B2(_04001_),
    .C1(_03764_),
    .X(_04002_));
 sky130_fd_sc_hd__o31ai_2 _11218_ (.A1(_03537_),
    .A2(_03958_),
    .A3(_03995_),
    .B1(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(_03915_),
    .A1(_04003_),
    .S(_03830_),
    .X(_04004_));
 sky130_fd_sc_hd__nand2_1 _11220_ (.A(_03886_),
    .B(_03868_),
    .Y(_04005_));
 sky130_fd_sc_hd__nor3_1 _11221_ (.A(_03460_),
    .B(_03467_),
    .C(_03525_),
    .Y(_04006_));
 sky130_fd_sc_hd__a31o_1 _11222_ (.A1(_02901_),
    .A2(_03838_),
    .A3(_03476_),
    .B1(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__nor2_1 _11223_ (.A(\gpout0.vpos[3] ),
    .B(_03523_),
    .Y(_04008_));
 sky130_fd_sc_hd__a21oi_1 _11224_ (.A1(_03900_),
    .A2(_03901_),
    .B1(_03464_),
    .Y(_04009_));
 sky130_fd_sc_hd__o211a_1 _11225_ (.A1(_04008_),
    .A2(_04009_),
    .B1(_03902_),
    .C1(_03461_),
    .X(_04010_));
 sky130_fd_sc_hd__nor2_1 _11226_ (.A(\gpout0.vpos[3] ),
    .B(_03531_),
    .Y(_04011_));
 sky130_fd_sc_hd__a31o_1 _11227_ (.A1(_03834_),
    .A2(_03517_),
    .A3(_03908_),
    .B1(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__a31o_1 _11228_ (.A1(_03852_),
    .A2(_03782_),
    .A3(_04008_),
    .B1(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__a2bb2o_1 _11229_ (.A1_N(\gpout0.vpos[4] ),
    .A2_N(_03524_),
    .B1(_03523_),
    .B2(\gpout0.vpos[3] ),
    .X(_04014_));
 sky130_fd_sc_hd__a221o_1 _11230_ (.A1(_03834_),
    .A2(_03524_),
    .B1(_03782_),
    .B2(_03849_),
    .C1(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__or4_1 _11231_ (.A(\gpout0.vpos[6] ),
    .B(_03838_),
    .C(_04008_),
    .D(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__a21oi_1 _11232_ (.A1(_03902_),
    .A2(_03461_),
    .B1(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__or4_1 _11233_ (.A(_04007_),
    .B(_04010_),
    .C(_04013_),
    .D(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__nor2_1 _11234_ (.A(_03461_),
    .B(_02901_),
    .Y(_04019_));
 sky130_fd_sc_hd__clkbuf_4 _11235_ (.A(_03523_),
    .X(_04020_));
 sky130_fd_sc_hd__nor4_1 _11236_ (.A(\gpout0.vpos[5] ),
    .B(_03517_),
    .C(_04020_),
    .D(_03524_),
    .Y(_04021_));
 sky130_fd_sc_hd__and4_1 _11237_ (.A(_03840_),
    .B(_03520_),
    .C(_03834_),
    .D(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__xnor2_1 _11238_ (.A(\gpout0.vpos[6] ),
    .B(_03460_),
    .Y(_04023_));
 sky130_fd_sc_hd__a221o_1 _11239_ (.A1(\gpout0.vpos[5] ),
    .A2(_03523_),
    .B1(_03524_),
    .B2(_03517_),
    .C1(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__xor2_1 _11240_ (.A(_03834_),
    .B(_03466_),
    .X(_04025_));
 sky130_fd_sc_hd__o221a_1 _11241_ (.A1(\gpout0.vpos[5] ),
    .A2(_03523_),
    .B1(_03524_),
    .B2(_03517_),
    .C1(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__and2b_1 _11242_ (.A_N(_04024_),
    .B(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__a31o_1 _11243_ (.A1(_03838_),
    .A2(_04019_),
    .A3(_04022_),
    .B1(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__and3b_1 _11244_ (.A_N(_03860_),
    .B(_04018_),
    .C(_04028_),
    .X(_04029_));
 sky130_fd_sc_hd__o21a_1 _11245_ (.A1(_04005_),
    .A2(_04029_),
    .B1(_03848_),
    .X(_04030_));
 sky130_fd_sc_hd__o2bb2a_1 _11246_ (.A1_N(_03896_),
    .A2_N(_04004_),
    .B1(_04030_),
    .B2(_03897_),
    .X(_04031_));
 sky130_fd_sc_hd__nand2_1 _11247_ (.A(\gpout0.hpos[2] ),
    .B(\gpout0.hpos[1] ),
    .Y(_04032_));
 sky130_fd_sc_hd__nor2_1 _11248_ (.A(_03500_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__and2_2 _11249_ (.A(_03476_),
    .B(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__xnor2_4 _11250_ (.A(_03466_),
    .B(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__nor2_1 _11251_ (.A(\gpout0.hpos[7] ),
    .B(_03512_),
    .Y(_04036_));
 sky130_fd_sc_hd__or2_1 _11252_ (.A(_03513_),
    .B(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_1 _11253_ (.A(\gpout0.hpos[3] ),
    .B(_04033_),
    .Y(_04038_));
 sky130_fd_sc_hd__or2_1 _11254_ (.A(_03503_),
    .B(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__buf_2 _11255_ (.A(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__nor2_1 _11256_ (.A(\gpout0.hpos[4] ),
    .B(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__and3b_1 _11257_ (.A_N(_03511_),
    .B(_03473_),
    .C(_03781_),
    .X(_04042_));
 sky130_fd_sc_hd__nor2_1 _11258_ (.A(_03512_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__or3b_1 _11259_ (.A(_04041_),
    .B(_04043_),
    .C_N(_04035_),
    .X(_04044_));
 sky130_fd_sc_hd__or2_1 _11260_ (.A(_04037_),
    .B(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__nand2_1 _11261_ (.A(\gpout0.hpos[5] ),
    .B(_03466_),
    .Y(_04046_));
 sky130_fd_sc_hd__o21ai_1 _11262_ (.A1(_04041_),
    .A2(_04043_),
    .B1(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__o21ba_1 _11263_ (.A1(_04037_),
    .A2(_04047_),
    .B1_N(_03513_),
    .X(_04048_));
 sky130_fd_sc_hd__xnor2_1 _11264_ (.A(\gpout0.hpos[8] ),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__xor2_1 _11265_ (.A(_04045_),
    .B(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__nand2_4 _11266_ (.A(_04035_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__or3b_2 _11267_ (.A(_03504_),
    .B(_03514_),
    .C_N(_04045_),
    .X(_04052_));
 sky130_fd_sc_hd__and3_1 _11268_ (.A(\gpout0.hpos[3] ),
    .B(\gpout0.hpos[4] ),
    .C(_04033_),
    .X(_04053_));
 sky130_fd_sc_hd__nand2b_1 _11269_ (.A_N(_04053_),
    .B(_03511_),
    .Y(_04054_));
 sky130_fd_sc_hd__nor2_1 _11270_ (.A(_04052_),
    .B(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__and4bb_4 _11271_ (.A_N(_03782_),
    .B_N(_04051_),
    .C(_04055_),
    .D(_04040_),
    .X(_04056_));
 sky130_fd_sc_hd__or3_1 _11272_ (.A(\gpout0.hpos[4] ),
    .B(_04040_),
    .C(_04052_),
    .X(_04057_));
 sky130_fd_sc_hd__or2_1 _11273_ (.A(_03460_),
    .B(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__nor2_1 _11274_ (.A(_04051_),
    .B(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__nand3b_2 _11275_ (.A_N(_04052_),
    .B(_04054_),
    .C(_04040_),
    .Y(_04060_));
 sky130_fd_sc_hd__nor2_1 _11276_ (.A(\gpout0.hpos[5] ),
    .B(_04053_),
    .Y(_04061_));
 sky130_fd_sc_hd__or2_2 _11277_ (.A(_04034_),
    .B(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__or2b_1 _11278_ (.A(_04060_),
    .B_N(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__nor2_1 _11279_ (.A(_04051_),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__or4b_2 _11280_ (.A(_03463_),
    .B(_04040_),
    .C(_04052_),
    .D_N(_04062_),
    .X(_04065_));
 sky130_fd_sc_hd__nor2_1 _11281_ (.A(_04051_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__or4b_2 _11282_ (.A(\gpout0.hpos[5] ),
    .B(_04052_),
    .C(_04054_),
    .D_N(_04040_),
    .X(_04067_));
 sky130_fd_sc_hd__nor2_1 _11283_ (.A(_04051_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__or3_1 _11284_ (.A(_04064_),
    .B(_04066_),
    .C(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__or2_2 _11285_ (.A(_04035_),
    .B(_04049_),
    .X(_04070_));
 sky130_fd_sc_hd__nand2_1 _11286_ (.A(_03460_),
    .B(_04040_),
    .Y(_04071_));
 sky130_fd_sc_hd__a21bo_1 _11287_ (.A1(_04070_),
    .A2(_04071_),
    .B1_N(_04055_),
    .X(_04072_));
 sky130_fd_sc_hd__or3_1 _11288_ (.A(_03474_),
    .B(_04062_),
    .C(_04060_),
    .X(_04073_));
 sky130_fd_sc_hd__or2_1 _11289_ (.A(_04046_),
    .B(_04057_),
    .X(_04074_));
 sky130_fd_sc_hd__nand2_1 _11290_ (.A(_04044_),
    .B(_04047_),
    .Y(_04075_));
 sky130_fd_sc_hd__xnor2_2 _11291_ (.A(_04037_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__a31o_1 _11292_ (.A1(_04072_),
    .A2(_04073_),
    .A3(_04074_),
    .B1(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__or3b_4 _11293_ (.A(_04059_),
    .B(_04069_),
    .C_N(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__nor3_4 _11294_ (.A(_04051_),
    .B(_04062_),
    .C(_04060_),
    .Y(_04079_));
 sky130_fd_sc_hd__or2b_2 _11295_ (.A(_04049_),
    .B_N(_04076_),
    .X(_04080_));
 sky130_fd_sc_hd__nor2_4 _11296_ (.A(_04074_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__or2_2 _11297_ (.A(_04035_),
    .B(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__nor2_4 _11298_ (.A(_04065_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__nor2_4 _11299_ (.A(_04067_),
    .B(_04082_),
    .Y(_04084_));
 sky130_fd_sc_hd__nor2_4 _11300_ (.A(_04058_),
    .B(_04070_),
    .Y(_04085_));
 sky130_fd_sc_hd__a211o_1 _11301_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_04085_),
    .B1(_03900_),
    .C1(_03849_),
    .X(_04086_));
 sky130_fd_sc_hd__a221o_1 _11302_ (.A1(\rbzero.debug_overlay.facingY[-7] ),
    .A2(_04083_),
    .B1(_04084_),
    .B2(\rbzero.debug_overlay.facingY[-6] ),
    .C1(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__a221o_1 _11303_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_04079_),
    .B1(_04081_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .C1(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__nor2_4 _11304_ (.A(_04063_),
    .B(_04070_),
    .Y(_04089_));
 sky130_fd_sc_hd__nor2_4 _11305_ (.A(_04073_),
    .B(_04080_),
    .Y(_04090_));
 sky130_fd_sc_hd__or4_2 _11306_ (.A(_03463_),
    .B(_04040_),
    .C(_04062_),
    .D(_04052_),
    .X(_04091_));
 sky130_fd_sc_hd__nor2_4 _11307_ (.A(_04051_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__nor3_4 _11308_ (.A(_03782_),
    .B(_04051_),
    .C(_04057_),
    .Y(_04093_));
 sky130_fd_sc_hd__a22o_1 _11309_ (.A1(\rbzero.debug_overlay.facingY[-3] ),
    .A2(_04092_),
    .B1(_04093_),
    .B2(\rbzero.debug_overlay.facingY[-1] ),
    .X(_04094_));
 sky130_fd_sc_hd__a221o_1 _11310_ (.A1(\rbzero.debug_overlay.facingY[-4] ),
    .A2(_04089_),
    .B1(_04090_),
    .B2(\rbzero.debug_overlay.facingY[-8] ),
    .C1(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__a211o_1 _11311_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_04078_),
    .B1(_04088_),
    .C1(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__a21oi_1 _11312_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(_04056_),
    .B1(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__a221o_1 _11313_ (.A1(\rbzero.debug_overlay.vplaneX[-7] ),
    .A2(_04083_),
    .B1(_04084_),
    .B2(\rbzero.debug_overlay.vplaneX[-6] ),
    .C1(\gpout0.vpos[3] ),
    .X(_04098_));
 sky130_fd_sc_hd__a221o_1 _11314_ (.A1(\rbzero.debug_overlay.vplaneX[-1] ),
    .A2(_04093_),
    .B1(_04056_),
    .B2(\rbzero.debug_overlay.vplaneX[-2] ),
    .C1(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__clkbuf_4 _11315_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_04100_));
 sky130_fd_sc_hd__a22o_1 _11316_ (.A1(\rbzero.debug_overlay.vplaneX[-8] ),
    .A2(_04090_),
    .B1(_04085_),
    .B2(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_4 _11317_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_04102_));
 sky130_fd_sc_hd__a22o_1 _11318_ (.A1(\rbzero.debug_overlay.vplaneX[-9] ),
    .A2(_04081_),
    .B1(_04089_),
    .B2(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__a211o_1 _11319_ (.A1(\rbzero.debug_overlay.vplaneX[-3] ),
    .A2(_04092_),
    .B1(_04101_),
    .C1(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__a211o_1 _11320_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_04079_),
    .B1(_04099_),
    .C1(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__a21oi_2 _11321_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_04078_),
    .B1(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a22o_1 _11322_ (.A1(\rbzero.debug_overlay.vplaneY[-4] ),
    .A2(_04089_),
    .B1(_04085_),
    .B2(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_04107_));
 sky130_fd_sc_hd__a221o_1 _11323_ (.A1(\rbzero.debug_overlay.vplaneY[-3] ),
    .A2(_04092_),
    .B1(_04090_),
    .B2(\rbzero.debug_overlay.vplaneY[-8] ),
    .C1(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_4 _11324_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_04109_));
 sky130_fd_sc_hd__a221o_1 _11325_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_04081_),
    .B1(_04084_),
    .B2(\rbzero.debug_overlay.vplaneY[-6] ),
    .C1(_03854_),
    .X(_04110_));
 sky130_fd_sc_hd__a21o_1 _11326_ (.A1(\rbzero.debug_overlay.vplaneY[-7] ),
    .A2(_04083_),
    .B1(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__a221o_1 _11327_ (.A1(\rbzero.debug_overlay.vplaneY[-1] ),
    .A2(_04093_),
    .B1(_04056_),
    .B2(_04109_),
    .C1(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__a211o_1 _11328_ (.A1(\rbzero.debug_overlay.vplaneY[0] ),
    .A2(_04079_),
    .B1(_04108_),
    .C1(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__a21oi_1 _11329_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(_04078_),
    .B1(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__o32a_1 _11330_ (.A1(_03903_),
    .A2(_04106_),
    .A3(_04114_),
    .B1(_03900_),
    .B2(_03852_),
    .X(_04115_));
 sky130_fd_sc_hd__o22a_1 _11331_ (.A1(_03902_),
    .A2(_03901_),
    .B1(_04097_),
    .B2(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__a211o_1 _11332_ (.A1(\rbzero.debug_overlay.facingX[-6] ),
    .A2(_04084_),
    .B1(_03901_),
    .C1(\gpout0.vpos[5] ),
    .X(_04117_));
 sky130_fd_sc_hd__a221o_1 _11333_ (.A1(\rbzero.debug_overlay.facingX[-7] ),
    .A2(_04083_),
    .B1(_04085_),
    .B2(\rbzero.debug_overlay.facingX[-5] ),
    .C1(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__a221o_1 _11334_ (.A1(\rbzero.debug_overlay.facingX[0] ),
    .A2(_04079_),
    .B1(_04081_),
    .B2(\rbzero.debug_overlay.facingX[-9] ),
    .C1(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__a22o_1 _11335_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_04089_),
    .B1(_04090_),
    .B2(\rbzero.debug_overlay.facingX[-8] ),
    .X(_04120_));
 sky130_fd_sc_hd__a221o_1 _11336_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_04092_),
    .B1(_04056_),
    .B2(\rbzero.debug_overlay.facingX[-2] ),
    .C1(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__a211o_1 _11337_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_04078_),
    .B1(_04119_),
    .C1(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__a21oi_1 _11338_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(_04093_),
    .B1(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__or2_1 _11339_ (.A(_04116_),
    .B(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__nor2_1 _11340_ (.A(_04076_),
    .B(_04091_),
    .Y(_04125_));
 sky130_fd_sc_hd__a211o_1 _11341_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_04125_),
    .B1(_03519_),
    .C1(\gpout0.vpos[3] ),
    .X(_04126_));
 sky130_fd_sc_hd__a221o_1 _11342_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_04083_),
    .B1(_04085_),
    .B2(\rbzero.debug_overlay.playerX[-5] ),
    .C1(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__a221o_1 _11343_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_04093_),
    .B1(_04084_),
    .B2(\rbzero.debug_overlay.playerX[-6] ),
    .C1(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__a22o_1 _11344_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_04068_),
    .B1(_04092_),
    .B2(\rbzero.debug_overlay.playerX[-3] ),
    .X(_04129_));
 sky130_fd_sc_hd__a22o_1 _11345_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(_04081_),
    .B1(_04089_),
    .B2(\rbzero.debug_overlay.playerX[-4] ),
    .X(_04130_));
 sky130_fd_sc_hd__a221o_1 _11346_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_04059_),
    .B1(_04090_),
    .B2(\rbzero.debug_overlay.playerX[-8] ),
    .C1(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__a221o_1 _11347_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_04064_),
    .B1(_04079_),
    .B2(\rbzero.debug_overlay.playerX[0] ),
    .C1(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__a211o_1 _11348_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_04066_),
    .B1(_04129_),
    .C1(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__a211o_1 _11349_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_04056_),
    .B1(_04128_),
    .C1(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__a211o_1 _11350_ (.A1(\rbzero.debug_overlay.playerY[5] ),
    .A2(_04125_),
    .B1(_03519_),
    .C1(_03854_),
    .X(_04135_));
 sky130_fd_sc_hd__a221o_1 _11351_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_04089_),
    .B1(_04083_),
    .B2(\rbzero.debug_overlay.playerY[-7] ),
    .C1(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__a221o_1 _11352_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_04056_),
    .B1(_04084_),
    .B2(\rbzero.debug_overlay.playerY[-6] ),
    .C1(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__a22o_1 _11353_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_04066_),
    .B1(_04068_),
    .B2(\rbzero.debug_overlay.playerY[2] ),
    .X(_04138_));
 sky130_fd_sc_hd__a22o_1 _11354_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(_04090_),
    .B1(_04085_),
    .B2(\rbzero.debug_overlay.playerY[-5] ),
    .X(_04139_));
 sky130_fd_sc_hd__a221o_1 _11355_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_04079_),
    .B1(_04081_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .C1(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__a221o_1 _11356_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_04064_),
    .B1(_04092_),
    .B2(\rbzero.debug_overlay.playerY[-3] ),
    .C1(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__a211o_1 _11357_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_04059_),
    .B1(_04138_),
    .C1(_04141_),
    .X(_04142_));
 sky130_fd_sc_hd__a211o_1 _11358_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_04093_),
    .B1(_04137_),
    .C1(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__and3b_1 _11359_ (.A_N(_03904_),
    .B(_04134_),
    .C(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__a21bo_1 _11360_ (.A1(_03519_),
    .A2(_04124_),
    .B1_N(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__nand2_1 _11361_ (.A(_03461_),
    .B(_02904_),
    .Y(_04146_));
 sky130_fd_sc_hd__or4_1 _11362_ (.A(_03467_),
    .B(_03502_),
    .C(_03525_),
    .D(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__a311oi_4 _11363_ (.A1(_03522_),
    .A2(_04145_),
    .A3(_04147_),
    .B1(_03910_),
    .C1(_03911_),
    .Y(_04148_));
 sky130_fd_sc_hd__o21a_1 _11364_ (.A1(_03522_),
    .A2(_04031_),
    .B1(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__buf_4 _11365_ (.A(_04149_),
    .X(net67));
 sky130_fd_sc_hd__mux2_1 _11366_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_03535_),
    .X(_04150_));
 sky130_fd_sc_hd__mux2_1 _11367_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_03709_),
    .X(_04151_));
 sky130_fd_sc_hd__mux2_1 _11368_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_03709_),
    .X(_04152_));
 sky130_fd_sc_hd__mux2_1 _11369_ (.A0(_04151_),
    .A1(_04152_),
    .S(_03666_),
    .X(_04153_));
 sky130_fd_sc_hd__mux2_1 _11370_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_03663_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_4 _11371_ (.A(_03696_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_4 _11372_ (.A(_03697_),
    .X(_04156_));
 sky130_fd_sc_hd__and3_1 _11373_ (.A(\rbzero.tex_g0[19] ),
    .B(_04155_),
    .C(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__a21o_1 _11374_ (.A1(\rbzero.tex_g0[18] ),
    .A2(_03617_),
    .B1(_03611_),
    .X(_04158_));
 sky130_fd_sc_hd__o221a_1 _11375_ (.A1(_03740_),
    .A2(_04154_),
    .B1(_04157_),
    .B2(_04158_),
    .C1(_03702_),
    .X(_04159_));
 sky130_fd_sc_hd__a211o_1 _11376_ (.A1(_03671_),
    .A2(_04153_),
    .B1(_04159_),
    .C1(_03704_),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_03709_),
    .X(_04161_));
 sky130_fd_sc_hd__mux2_1 _11378_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_03709_),
    .X(_04162_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(_04161_),
    .A1(_04162_),
    .S(_03677_),
    .X(_04163_));
 sky130_fd_sc_hd__and2_1 _11380_ (.A(\rbzero.tex_g0[30] ),
    .B(_03700_),
    .X(_04164_));
 sky130_fd_sc_hd__a31o_1 _11381_ (.A1(\rbzero.tex_g0[31] ),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_03659_),
    .X(_04165_));
 sky130_fd_sc_hd__mux2_1 _11382_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_03709_),
    .X(_04166_));
 sky130_fd_sc_hd__o221a_1 _11383_ (.A1(_04164_),
    .A2(_04165_),
    .B1(_04166_),
    .B2(_03740_),
    .C1(_03670_),
    .X(_04167_));
 sky130_fd_sc_hd__a211o_1 _11384_ (.A1(_03674_),
    .A2(_04163_),
    .B1(_04167_),
    .C1(_03679_),
    .X(_04168_));
 sky130_fd_sc_hd__mux2_1 _11385_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_03615_),
    .X(_04169_));
 sky130_fd_sc_hd__mux2_1 _11386_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_03615_),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _11387_ (.A0(_04169_),
    .A1(_04170_),
    .S(_03823_),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _11388_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_03615_),
    .X(_04172_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_03615_),
    .X(_04173_));
 sky130_fd_sc_hd__mux2_1 _11390_ (.A0(_04172_),
    .A1(_04173_),
    .S(_03635_),
    .X(_04174_));
 sky130_fd_sc_hd__mux2_1 _11391_ (.A0(_04171_),
    .A1(_04174_),
    .S(_03702_),
    .X(_04175_));
 sky130_fd_sc_hd__mux2_1 _11392_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_03709_),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _11393_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_03662_),
    .X(_04177_));
 sky130_fd_sc_hd__or2_1 _11394_ (.A(_03739_),
    .B(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__buf_4 _11395_ (.A(_03669_),
    .X(_04179_));
 sky130_fd_sc_hd__o211a_1 _11396_ (.A1(_03612_),
    .A2(_04176_),
    .B1(_04178_),
    .C1(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__mux2_1 _11397_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_03662_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _11398_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_03662_),
    .X(_04182_));
 sky130_fd_sc_hd__mux2_1 _11399_ (.A0(_04181_),
    .A1(_04182_),
    .S(_03635_),
    .X(_04183_));
 sky130_fd_sc_hd__a21o_1 _11400_ (.A1(_03702_),
    .A2(_04183_),
    .B1(_03624_),
    .X(_04184_));
 sky130_fd_sc_hd__o221a_1 _11401_ (.A1(_03704_),
    .A2(_04175_),
    .B1(_04180_),
    .B2(_04184_),
    .C1(_03684_),
    .X(_04185_));
 sky130_fd_sc_hd__a311o_1 _11402_ (.A1(_03688_),
    .A2(_04160_),
    .A3(_04168_),
    .B1(_04185_),
    .C1(_03719_),
    .X(_04186_));
 sky130_fd_sc_hd__mux2_1 _11403_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_03700_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_8 _11404_ (.A(_03614_),
    .X(_04188_));
 sky130_fd_sc_hd__buf_6 _11405_ (.A(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__mux2_1 _11406_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__mux2_1 _11407_ (.A0(_04187_),
    .A1(_04190_),
    .S(_03740_),
    .X(_04191_));
 sky130_fd_sc_hd__buf_4 _11408_ (.A(_03656_),
    .X(_04192_));
 sky130_fd_sc_hd__mux2_1 _11409_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04189_),
    .X(_04193_));
 sky130_fd_sc_hd__and3_1 _11410_ (.A(\rbzero.tex_g0[51] ),
    .B(_03729_),
    .C(_03730_),
    .X(_04194_));
 sky130_fd_sc_hd__a21o_1 _11411_ (.A1(\rbzero.tex_g0[50] ),
    .A2(_03727_),
    .B1(_03652_),
    .X(_04195_));
 sky130_fd_sc_hd__o221a_1 _11412_ (.A1(_04192_),
    .A2(_04193_),
    .B1(_04194_),
    .B2(_04195_),
    .C1(_03607_),
    .X(_04196_));
 sky130_fd_sc_hd__a211o_1 _11413_ (.A1(_03671_),
    .A2(_04191_),
    .B1(_04196_),
    .C1(_03648_),
    .X(_04197_));
 sky130_fd_sc_hd__buf_4 _11414_ (.A(_03607_),
    .X(_04198_));
 sky130_fd_sc_hd__mux2_1 _11415_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_03700_),
    .X(_04199_));
 sky130_fd_sc_hd__mux2_1 _11416_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04189_),
    .X(_04200_));
 sky130_fd_sc_hd__mux2_1 _11417_ (.A0(_04199_),
    .A1(_04200_),
    .S(_03740_),
    .X(_04201_));
 sky130_fd_sc_hd__mux2_1 _11418_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_03700_),
    .X(_04202_));
 sky130_fd_sc_hd__mux2_1 _11419_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_03699_),
    .X(_04203_));
 sky130_fd_sc_hd__or2_1 _11420_ (.A(_03652_),
    .B(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__o211a_1 _11421_ (.A1(_03917_),
    .A2(_04202_),
    .B1(_04204_),
    .C1(_03689_),
    .X(_04205_));
 sky130_fd_sc_hd__a211o_1 _11422_ (.A1(_04198_),
    .A2(_04201_),
    .B1(_04205_),
    .C1(_03721_),
    .X(_04206_));
 sky130_fd_sc_hd__mux2_1 _11423_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_03699_),
    .X(_04207_));
 sky130_fd_sc_hd__mux2_1 _11424_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04188_),
    .X(_04208_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(_04207_),
    .A1(_04208_),
    .S(_03739_),
    .X(_04209_));
 sky130_fd_sc_hd__mux2_1 _11426_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_03699_),
    .X(_04210_));
 sky130_fd_sc_hd__mux2_1 _11427_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_03614_),
    .X(_04211_));
 sky130_fd_sc_hd__or2_1 _11428_ (.A(_03610_),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__o211a_1 _11429_ (.A1(_03656_),
    .A2(_04210_),
    .B1(_04212_),
    .C1(_03669_),
    .X(_04213_));
 sky130_fd_sc_hd__a211o_1 _11430_ (.A1(_03607_),
    .A2(_04209_),
    .B1(_04213_),
    .C1(_03627_),
    .X(_04214_));
 sky130_fd_sc_hd__mux2_1 _11431_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_04188_),
    .X(_04215_));
 sky130_fd_sc_hd__mux2_1 _11432_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04188_),
    .X(_04216_));
 sky130_fd_sc_hd__mux2_1 _11433_ (.A0(_04215_),
    .A1(_04216_),
    .S(_03739_),
    .X(_04217_));
 sky130_fd_sc_hd__mux2_1 _11434_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04188_),
    .X(_04218_));
 sky130_fd_sc_hd__and3_1 _11435_ (.A(\rbzero.tex_g0[43] ),
    .B(_03696_),
    .C(_03697_),
    .X(_04219_));
 sky130_fd_sc_hd__a21o_1 _11436_ (.A1(\rbzero.tex_g0[42] ),
    .A2(_03649_),
    .B1(_03610_),
    .X(_04220_));
 sky130_fd_sc_hd__o221a_1 _11437_ (.A1(_03656_),
    .A2(_04218_),
    .B1(_04219_),
    .B2(_04220_),
    .C1(_03606_),
    .X(_04221_));
 sky130_fd_sc_hd__a211o_1 _11438_ (.A1(_04179_),
    .A2(_04217_),
    .B1(_04221_),
    .C1(_03624_),
    .X(_04222_));
 sky130_fd_sc_hd__a31o_1 _11439_ (.A1(_03685_),
    .A2(_04214_),
    .A3(_04222_),
    .B1(_03718_),
    .X(_04223_));
 sky130_fd_sc_hd__a31o_1 _11440_ (.A1(_03688_),
    .A2(_04197_),
    .A3(_04206_),
    .B1(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__o31ai_1 _11441_ (.A1(_03538_),
    .A2(_03539_),
    .A3(_03640_),
    .B1(_03996_),
    .Y(_04225_));
 sky130_fd_sc_hd__nor3_1 _11442_ (.A(_03936_),
    .B(_03630_),
    .C(_03639_),
    .Y(_04226_));
 sky130_fd_sc_hd__o21a_1 _11443_ (.A1(_03619_),
    .A2(_04226_),
    .B1(_03633_),
    .X(_04227_));
 sky130_fd_sc_hd__o211a_1 _11444_ (.A1(_04225_),
    .A2(_04227_),
    .B1(net41),
    .C1(_03541_),
    .X(_04228_));
 sky130_fd_sc_hd__a31o_1 _11445_ (.A1(_03764_),
    .A2(_04186_),
    .A3(_04224_),
    .B1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(_04150_),
    .A1(_04229_),
    .S(_03830_),
    .X(_04230_));
 sky130_fd_sc_hd__or2_1 _11447_ (.A(_03896_),
    .B(_03847_),
    .X(_04231_));
 sky130_fd_sc_hd__inv_2 _11448_ (.A(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__a211o_1 _11449_ (.A1(_03896_),
    .A2(_04230_),
    .B1(_04232_),
    .C1(_03522_),
    .X(_04233_));
 sky130_fd_sc_hd__and2_1 _11450_ (.A(_03912_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__buf_4 _11451_ (.A(_04234_),
    .X(net62));
 sky130_fd_sc_hd__mux2_1 _11452_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_03535_),
    .X(_04235_));
 sky130_fd_sc_hd__nor2_2 _11453_ (.A(_03540_),
    .B(_03632_),
    .Y(_04236_));
 sky130_fd_sc_hd__or2_1 _11454_ (.A(\rbzero.row_render.texu[2] ),
    .B(_04198_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_1 _11455_ (.A(\rbzero.row_render.texu[2] ),
    .B(_04198_),
    .Y(_04238_));
 sky130_fd_sc_hd__a311o_1 _11456_ (.A1(_03540_),
    .A2(_04237_),
    .A3(_04238_),
    .B1(_03997_),
    .C1(_03764_),
    .X(_04239_));
 sky130_fd_sc_hd__mux2_1 _11457_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_03617_),
    .X(_04240_));
 sky130_fd_sc_hd__mux2_1 _11458_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_03700_),
    .X(_04241_));
 sky130_fd_sc_hd__mux2_1 _11459_ (.A0(_04240_),
    .A1(_04241_),
    .S(_03612_),
    .X(_04242_));
 sky130_fd_sc_hd__mux2_1 _11460_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_03700_),
    .X(_04243_));
 sky130_fd_sc_hd__mux2_1 _11461_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_03700_),
    .X(_04244_));
 sky130_fd_sc_hd__mux2_1 _11462_ (.A0(_04243_),
    .A1(_04244_),
    .S(_03740_),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_1 _11463_ (.A0(_04242_),
    .A1(_04245_),
    .S(_03671_),
    .X(_04246_));
 sky130_fd_sc_hd__buf_6 _11464_ (.A(_03649_),
    .X(_04247_));
 sky130_fd_sc_hd__mux2_1 _11465_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__mux2_1 _11466_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04247_),
    .X(_04249_));
 sky130_fd_sc_hd__mux2_1 _11467_ (.A0(_04248_),
    .A1(_04249_),
    .S(_03612_),
    .X(_04250_));
 sky130_fd_sc_hd__and2_1 _11468_ (.A(\rbzero.tex_g1[26] ),
    .B(_03664_),
    .X(_04251_));
 sky130_fd_sc_hd__a31o_1 _11469_ (.A1(\rbzero.tex_g1[27] ),
    .A2(_03729_),
    .A3(_03730_),
    .B1(_03652_),
    .X(_04252_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04247_),
    .X(_04253_));
 sky130_fd_sc_hd__o221a_1 _11471_ (.A1(_04251_),
    .A2(_04252_),
    .B1(_04253_),
    .B2(_03917_),
    .C1(_03674_),
    .X(_04254_));
 sky130_fd_sc_hd__a211o_1 _11472_ (.A1(_03671_),
    .A2(_04250_),
    .B1(_04254_),
    .C1(_03721_),
    .X(_04255_));
 sky130_fd_sc_hd__o211a_1 _11473_ (.A1(_03648_),
    .A2(_04246_),
    .B1(_04255_),
    .C1(_03688_),
    .X(_04256_));
 sky130_fd_sc_hd__mux2_1 _11474_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_03618_),
    .X(_04257_));
 sky130_fd_sc_hd__and2_1 _11475_ (.A(\rbzero.tex_g1[14] ),
    .B(_03618_),
    .X(_04258_));
 sky130_fd_sc_hd__a31o_1 _11476_ (.A1(\rbzero.tex_g1[15] ),
    .A2(_03729_),
    .A3(_03730_),
    .B1(_03612_),
    .X(_04259_));
 sky130_fd_sc_hd__o221a_1 _11477_ (.A1(_03726_),
    .A2(_04257_),
    .B1(_04258_),
    .B2(_04259_),
    .C1(_03671_),
    .X(_04260_));
 sky130_fd_sc_hd__mux2_1 _11478_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_03618_),
    .X(_04261_));
 sky130_fd_sc_hd__and2_1 _11479_ (.A(\rbzero.tex_g1[8] ),
    .B(_03618_),
    .X(_04262_));
 sky130_fd_sc_hd__a31o_1 _11480_ (.A1(\rbzero.tex_g1[9] ),
    .A2(_03729_),
    .A3(_03730_),
    .B1(_03917_),
    .X(_04263_));
 sky130_fd_sc_hd__o221a_1 _11481_ (.A1(_03661_),
    .A2(_04261_),
    .B1(_04262_),
    .B2(_04263_),
    .C1(_04198_),
    .X(_04264_));
 sky130_fd_sc_hd__mux2_1 _11482_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_04247_),
    .X(_04265_));
 sky130_fd_sc_hd__mux2_1 _11483_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_04247_),
    .X(_04266_));
 sky130_fd_sc_hd__mux2_1 _11484_ (.A0(_04265_),
    .A1(_04266_),
    .S(_03612_),
    .X(_04267_));
 sky130_fd_sc_hd__and2_1 _11485_ (.A(\rbzero.tex_g1[2] ),
    .B(_03664_),
    .X(_04268_));
 sky130_fd_sc_hd__a31o_1 _11486_ (.A1(\rbzero.tex_g1[3] ),
    .A2(_03729_),
    .A3(_03730_),
    .B1(_03652_),
    .X(_04269_));
 sky130_fd_sc_hd__mux2_1 _11487_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[0] ),
    .S(_03727_),
    .X(_04270_));
 sky130_fd_sc_hd__o221a_1 _11488_ (.A1(_04268_),
    .A2(_04269_),
    .B1(_04270_),
    .B2(_03917_),
    .C1(_03674_),
    .X(_04271_));
 sky130_fd_sc_hd__a211o_1 _11489_ (.A1(_03671_),
    .A2(_04267_),
    .B1(_04271_),
    .C1(_03648_),
    .X(_04272_));
 sky130_fd_sc_hd__o311a_1 _11490_ (.A1(_03721_),
    .A2(_04260_),
    .A3(_04264_),
    .B1(_04272_),
    .C1(_03685_),
    .X(_04273_));
 sky130_fd_sc_hd__mux2_1 _11491_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04247_),
    .X(_04274_));
 sky130_fd_sc_hd__mux2_1 _11492_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04247_),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_1 _11493_ (.A0(_04274_),
    .A1(_04275_),
    .S(_03612_),
    .X(_04276_));
 sky130_fd_sc_hd__mux2_1 _11494_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04247_),
    .X(_04277_));
 sky130_fd_sc_hd__mux2_1 _11495_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_03617_),
    .X(_04278_));
 sky130_fd_sc_hd__mux2_1 _11496_ (.A0(_04277_),
    .A1(_04278_),
    .S(_03917_),
    .X(_04279_));
 sky130_fd_sc_hd__mux2_1 _11497_ (.A0(_04276_),
    .A1(_04279_),
    .S(_03671_),
    .X(_04280_));
 sky130_fd_sc_hd__and2_1 _11498_ (.A(\rbzero.tex_g1[62] ),
    .B(_03925_),
    .X(_04281_));
 sky130_fd_sc_hd__a31o_1 _11499_ (.A1(\rbzero.tex_g1[63] ),
    .A2(_03729_),
    .A3(_03730_),
    .B1(_03661_),
    .X(_04282_));
 sky130_fd_sc_hd__mux2_1 _11500_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_03618_),
    .X(_04283_));
 sky130_fd_sc_hd__o221a_1 _11501_ (.A1(_04281_),
    .A2(_04282_),
    .B1(_04283_),
    .B2(_03726_),
    .C1(_03671_),
    .X(_04284_));
 sky130_fd_sc_hd__mux2_1 _11502_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_03664_),
    .X(_04285_));
 sky130_fd_sc_hd__mux2_1 _11503_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_03727_),
    .X(_04286_));
 sky130_fd_sc_hd__mux2_1 _11504_ (.A0(_04285_),
    .A1(_04286_),
    .S(_03917_),
    .X(_04287_));
 sky130_fd_sc_hd__a21o_1 _11505_ (.A1(_04198_),
    .A2(_04287_),
    .B1(_03721_),
    .X(_04288_));
 sky130_fd_sc_hd__o221a_1 _11506_ (.A1(_03648_),
    .A2(_04280_),
    .B1(_04284_),
    .B2(_04288_),
    .C1(_03688_),
    .X(_04289_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_03727_),
    .X(_04290_));
 sky130_fd_sc_hd__mux2_1 _11508_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_03727_),
    .X(_04291_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(_04290_),
    .A1(_04291_),
    .S(_03920_),
    .X(_04292_));
 sky130_fd_sc_hd__and3_1 _11510_ (.A(\rbzero.tex_g1[39] ),
    .B(_03729_),
    .C(_03730_),
    .X(_04293_));
 sky130_fd_sc_hd__a21o_1 _11511_ (.A1(\rbzero.tex_g1[38] ),
    .A2(_03733_),
    .B1(_03660_),
    .X(_04294_));
 sky130_fd_sc_hd__mux2_1 _11512_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_03727_),
    .X(_04295_));
 sky130_fd_sc_hd__o221a_1 _11513_ (.A1(_04293_),
    .A2(_04294_),
    .B1(_04295_),
    .B2(_03726_),
    .C1(_03689_),
    .X(_04296_));
 sky130_fd_sc_hd__a211o_1 _11514_ (.A1(_04198_),
    .A2(_04292_),
    .B1(_04296_),
    .C1(_03648_),
    .X(_04297_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_03727_),
    .X(_04298_));
 sky130_fd_sc_hd__mux2_1 _11516_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_03727_),
    .X(_04299_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(_04298_),
    .A1(_04299_),
    .S(_03612_),
    .X(_04300_));
 sky130_fd_sc_hd__and2_1 _11518_ (.A(\rbzero.tex_g1[46] ),
    .B(_03733_),
    .X(_04301_));
 sky130_fd_sc_hd__a31o_1 _11519_ (.A1(\rbzero.tex_g1[47] ),
    .A2(_03729_),
    .A3(_03730_),
    .B1(_03660_),
    .X(_04302_));
 sky130_fd_sc_hd__mux2_1 _11520_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_03727_),
    .X(_04303_));
 sky130_fd_sc_hd__o221a_1 _11521_ (.A1(_04301_),
    .A2(_04302_),
    .B1(_04303_),
    .B2(_03917_),
    .C1(_03689_),
    .X(_04304_));
 sky130_fd_sc_hd__a211o_1 _11522_ (.A1(_04198_),
    .A2(_04300_),
    .B1(_04304_),
    .C1(_03721_),
    .X(_04305_));
 sky130_fd_sc_hd__a31o_1 _11523_ (.A1(_03685_),
    .A2(_04297_),
    .A3(_04305_),
    .B1(_03718_),
    .X(_04306_));
 sky130_fd_sc_hd__o32a_1 _11524_ (.A1(_03719_),
    .A2(_04256_),
    .A3(_04273_),
    .B1(_04289_),
    .B2(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__a2bb2o_1 _11525_ (.A1_N(_04236_),
    .A2_N(_04239_),
    .B1(_03764_),
    .B2(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_1 _11526_ (.A0(_04235_),
    .A1(_04308_),
    .S(_03830_),
    .X(_04309_));
 sky130_fd_sc_hd__inv_2 _11527_ (.A(_04028_),
    .Y(_04310_));
 sky130_fd_sc_hd__nor2_1 _11528_ (.A(_03860_),
    .B(_04005_),
    .Y(_04311_));
 sky130_fd_sc_hd__a41o_1 _11529_ (.A1(_03848_),
    .A2(_04018_),
    .A3(_04310_),
    .A4(_04311_),
    .B1(_03897_),
    .X(_04312_));
 sky130_fd_sc_hd__o21a_1 _11530_ (.A1(_03534_),
    .A2(_04309_),
    .B1(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__o21ai_4 _11531_ (.A1(_03522_),
    .A2(_04313_),
    .B1(_04148_),
    .Y(_04314_));
 sky130_fd_sc_hd__clkinv_2 _11532_ (.A(_04314_),
    .Y(net63));
 sky130_fd_sc_hd__mux2_1 _11533_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_03535_),
    .X(_04315_));
 sky130_fd_sc_hd__mux2_1 _11534_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_04189_),
    .X(_04316_));
 sky130_fd_sc_hd__mux2_1 _11535_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_03732_),
    .X(_04317_));
 sky130_fd_sc_hd__mux2_1 _11536_ (.A0(_04316_),
    .A1(_04317_),
    .S(_03740_),
    .X(_04318_));
 sky130_fd_sc_hd__and2_1 _11537_ (.A(\rbzero.tex_b0[62] ),
    .B(_03617_),
    .X(_04319_));
 sky130_fd_sc_hd__a31o_1 _11538_ (.A1(\rbzero.tex_b0[63] ),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_03611_),
    .X(_04320_));
 sky130_fd_sc_hd__mux2_1 _11539_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_04189_),
    .X(_04321_));
 sky130_fd_sc_hd__o221a_1 _11540_ (.A1(_04319_),
    .A2(_04320_),
    .B1(_04321_),
    .B2(_04192_),
    .C1(_04179_),
    .X(_04322_));
 sky130_fd_sc_hd__a211o_1 _11541_ (.A1(_04198_),
    .A2(_04318_),
    .B1(_04322_),
    .C1(_03721_),
    .X(_04323_));
 sky130_fd_sc_hd__mux2_1 _11542_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_03732_),
    .X(_04324_));
 sky130_fd_sc_hd__mux2_1 _11543_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_03732_),
    .X(_04325_));
 sky130_fd_sc_hd__mux2_1 _11544_ (.A0(_04324_),
    .A1(_04325_),
    .S(_03660_),
    .X(_04326_));
 sky130_fd_sc_hd__mux2_1 _11545_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_03732_),
    .X(_04327_));
 sky130_fd_sc_hd__and3_1 _11546_ (.A(\rbzero.tex_b0[55] ),
    .B(_04155_),
    .C(_04156_),
    .X(_04328_));
 sky130_fd_sc_hd__a21o_1 _11547_ (.A1(\rbzero.tex_b0[54] ),
    .A2(_04247_),
    .B1(_03652_),
    .X(_04329_));
 sky130_fd_sc_hd__o221a_1 _11548_ (.A1(_04192_),
    .A2(_04327_),
    .B1(_04328_),
    .B2(_04329_),
    .C1(_04179_),
    .X(_04330_));
 sky130_fd_sc_hd__a211o_1 _11549_ (.A1(_03674_),
    .A2(_04326_),
    .B1(_04330_),
    .C1(_03704_),
    .X(_04331_));
 sky130_fd_sc_hd__mux2_1 _11550_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_03709_),
    .X(_04332_));
 sky130_fd_sc_hd__and3_1 _11551_ (.A(\rbzero.tex_b0[35] ),
    .B(_04155_),
    .C(_04156_),
    .X(_04333_));
 sky130_fd_sc_hd__a21o_1 _11552_ (.A1(\rbzero.tex_b0[34] ),
    .A2(_04247_),
    .B1(_03652_),
    .X(_04334_));
 sky130_fd_sc_hd__o221a_1 _11553_ (.A1(_03740_),
    .A2(_04332_),
    .B1(_04333_),
    .B2(_04334_),
    .C1(_03702_),
    .X(_04335_));
 sky130_fd_sc_hd__and2_1 _11554_ (.A(\rbzero.tex_b0[38] ),
    .B(_03617_),
    .X(_04336_));
 sky130_fd_sc_hd__a31o_1 _11555_ (.A1(\rbzero.tex_b0[39] ),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_03611_),
    .X(_04337_));
 sky130_fd_sc_hd__mux2_1 _11556_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04189_),
    .X(_04338_));
 sky130_fd_sc_hd__o221a_1 _11557_ (.A1(_04336_),
    .A2(_04337_),
    .B1(_04338_),
    .B2(_04192_),
    .C1(_04179_),
    .X(_04339_));
 sky130_fd_sc_hd__mux2_1 _11558_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_03699_),
    .X(_04340_));
 sky130_fd_sc_hd__mux2_1 _11559_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_04188_),
    .X(_04341_));
 sky130_fd_sc_hd__mux2_1 _11560_ (.A0(_04340_),
    .A1(_04341_),
    .S(_03659_),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _11561_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_04188_),
    .X(_04343_));
 sky130_fd_sc_hd__and3_1 _11562_ (.A(\rbzero.tex_b0[43] ),
    .B(_03696_),
    .C(_03697_),
    .X(_04344_));
 sky130_fd_sc_hd__a21o_1 _11563_ (.A1(\rbzero.tex_b0[42] ),
    .A2(_03649_),
    .B1(_03823_),
    .X(_04345_));
 sky130_fd_sc_hd__o221a_1 _11564_ (.A1(_03656_),
    .A2(_04343_),
    .B1(_04344_),
    .B2(_04345_),
    .C1(_03606_),
    .X(_04346_));
 sky130_fd_sc_hd__a211o_1 _11565_ (.A1(_04179_),
    .A2(_04342_),
    .B1(_04346_),
    .C1(_03624_),
    .X(_04347_));
 sky130_fd_sc_hd__o311a_1 _11566_ (.A1(_03704_),
    .A2(_04335_),
    .A3(_04339_),
    .B1(_04347_),
    .C1(_03684_),
    .X(_04348_));
 sky130_fd_sc_hd__a311o_1 _11567_ (.A1(_03688_),
    .A2(_04323_),
    .A3(_04331_),
    .B1(_04348_),
    .C1(_03718_),
    .X(_04349_));
 sky130_fd_sc_hd__mux2_1 _11568_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04189_),
    .X(_04350_));
 sky130_fd_sc_hd__mux2_1 _11569_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_03732_),
    .X(_04351_));
 sky130_fd_sc_hd__mux2_1 _11570_ (.A0(_04350_),
    .A1(_04351_),
    .S(_03740_),
    .X(_04352_));
 sky130_fd_sc_hd__and2_1 _11571_ (.A(\rbzero.tex_b0[22] ),
    .B(_03617_),
    .X(_04353_));
 sky130_fd_sc_hd__a31o_1 _11572_ (.A1(\rbzero.tex_b0[23] ),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_03611_),
    .X(_04354_));
 sky130_fd_sc_hd__mux2_1 _11573_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04189_),
    .X(_04355_));
 sky130_fd_sc_hd__o221a_1 _11574_ (.A1(_04353_),
    .A2(_04354_),
    .B1(_04355_),
    .B2(_04192_),
    .C1(_04179_),
    .X(_04356_));
 sky130_fd_sc_hd__a211o_1 _11575_ (.A1(_04198_),
    .A2(_04352_),
    .B1(_04356_),
    .C1(_03704_),
    .X(_04357_));
 sky130_fd_sc_hd__mux2_1 _11576_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_03732_),
    .X(_04358_));
 sky130_fd_sc_hd__mux2_1 _11577_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_03732_),
    .X(_04359_));
 sky130_fd_sc_hd__mux2_1 _11578_ (.A0(_04358_),
    .A1(_04359_),
    .S(_03666_),
    .X(_04360_));
 sky130_fd_sc_hd__and2_1 _11579_ (.A(\rbzero.tex_b0[26] ),
    .B(_03617_),
    .X(_04361_));
 sky130_fd_sc_hd__a31o_1 _11580_ (.A1(\rbzero.tex_b0[27] ),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_03611_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_1 _11581_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04189_),
    .X(_04363_));
 sky130_fd_sc_hd__o221a_1 _11582_ (.A1(_04361_),
    .A2(_04362_),
    .B1(_04363_),
    .B2(_04192_),
    .C1(_03607_),
    .X(_04364_));
 sky130_fd_sc_hd__a211o_1 _11583_ (.A1(_03671_),
    .A2(_04360_),
    .B1(_04364_),
    .C1(_03679_),
    .X(_04365_));
 sky130_fd_sc_hd__and2_1 _11584_ (.A(\rbzero.tex_b0[10] ),
    .B(_03700_),
    .X(_04366_));
 sky130_fd_sc_hd__a31o_1 _11585_ (.A1(\rbzero.tex_b0[11] ),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_03659_),
    .X(_04367_));
 sky130_fd_sc_hd__mux2_1 _11586_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_03709_),
    .X(_04368_));
 sky130_fd_sc_hd__o221a_1 _11587_ (.A1(_04366_),
    .A2(_04367_),
    .B1(_04368_),
    .B2(_03740_),
    .C1(_03702_),
    .X(_04369_));
 sky130_fd_sc_hd__and2_1 _11588_ (.A(\rbzero.tex_b0[14] ),
    .B(_03617_),
    .X(_04370_));
 sky130_fd_sc_hd__a31o_1 _11589_ (.A1(\rbzero.tex_b0[15] ),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_03611_),
    .X(_04371_));
 sky130_fd_sc_hd__mux2_1 _11590_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_03732_),
    .X(_04372_));
 sky130_fd_sc_hd__o221a_1 _11591_ (.A1(_04370_),
    .A2(_04371_),
    .B1(_04372_),
    .B2(_04192_),
    .C1(_04179_),
    .X(_04373_));
 sky130_fd_sc_hd__mux2_1 _11592_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_03699_),
    .X(_04374_));
 sky130_fd_sc_hd__or2_1 _11593_ (.A(_03652_),
    .B(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__buf_4 _11594_ (.A(_03615_),
    .X(_04376_));
 sky130_fd_sc_hd__mux2_1 _11595_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__o21a_1 _11596_ (.A1(_03656_),
    .A2(_04377_),
    .B1(_03669_),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_1 _11597_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04188_),
    .X(_04379_));
 sky130_fd_sc_hd__mux2_1 _11598_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_04188_),
    .X(_04380_));
 sky130_fd_sc_hd__mux2_1 _11599_ (.A0(_04379_),
    .A1(_04380_),
    .S(_03739_),
    .X(_04381_));
 sky130_fd_sc_hd__a221o_1 _11600_ (.A1(_04375_),
    .A2(_04378_),
    .B1(_04381_),
    .B2(_03607_),
    .C1(_03627_),
    .X(_04382_));
 sky130_fd_sc_hd__o311a_1 _11601_ (.A1(_03679_),
    .A2(_04369_),
    .A3(_04373_),
    .B1(_03684_),
    .C1(_04382_),
    .X(_04383_));
 sky130_fd_sc_hd__a311o_1 _11602_ (.A1(_03688_),
    .A2(_04357_),
    .A3(_04365_),
    .B1(_04383_),
    .C1(_03719_),
    .X(_04384_));
 sky130_fd_sc_hd__a311o_1 _11603_ (.A1(_04179_),
    .A2(_04192_),
    .A3(_03768_),
    .B1(_03631_),
    .C1(\rbzero.row_render.side ),
    .X(_04385_));
 sky130_fd_sc_hd__and3_1 _11604_ (.A(\rbzero.row_render.wall[1] ),
    .B(_03997_),
    .C(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__o311a_1 _11605_ (.A1(_03642_),
    .A2(_04225_),
    .A3(_04386_),
    .B1(_03541_),
    .C1(_03537_),
    .X(_04387_));
 sky130_fd_sc_hd__a31o_1 _11606_ (.A1(_03764_),
    .A2(_04349_),
    .A3(_04384_),
    .B1(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__mux2_1 _11607_ (.A0(_04315_),
    .A1(_04388_),
    .S(_03830_),
    .X(_04389_));
 sky130_fd_sc_hd__o21a_1 _11608_ (.A1(_04018_),
    .A2(_04028_),
    .B1(_04311_),
    .X(_04390_));
 sky130_fd_sc_hd__or4bb_1 _11609_ (.A(_03896_),
    .B(_04390_),
    .C_N(_03518_),
    .D_N(_03529_),
    .X(_04391_));
 sky130_fd_sc_hd__o211a_1 _11610_ (.A1(_03534_),
    .A2(_04389_),
    .B1(_04391_),
    .C1(_04231_),
    .X(_04392_));
 sky130_fd_sc_hd__o21ai_4 _11611_ (.A1(_03522_),
    .A2(_04392_),
    .B1(_03912_),
    .Y(_04393_));
 sky130_fd_sc_hd__inv_2 _11612_ (.A(_04393_),
    .Y(net64));
 sky130_fd_sc_hd__mux2_1 _11613_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_03535_),
    .X(_04394_));
 sky130_fd_sc_hd__a21oi_1 _11614_ (.A1(_04198_),
    .A2(_03661_),
    .B1(_03630_),
    .Y(_04395_));
 sky130_fd_sc_hd__o211a_1 _11615_ (.A1(_04395_),
    .A2(_03998_),
    .B1(_03643_),
    .C1(\rbzero.row_render.wall[1] ),
    .X(_04396_));
 sky130_fd_sc_hd__a31o_1 _11616_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_03729_),
    .A3(_03730_),
    .B1(_03996_),
    .X(_04397_));
 sky130_fd_sc_hd__nor2_1 _11617_ (.A(_03621_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__mux2_1 _11618_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_03732_),
    .X(_04399_));
 sky130_fd_sc_hd__mux2_1 _11619_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_03662_),
    .X(_04400_));
 sky130_fd_sc_hd__or2_1 _11620_ (.A(_03611_),
    .B(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__o211a_1 _11621_ (.A1(_04192_),
    .A2(_04399_),
    .B1(_04401_),
    .C1(_03702_),
    .X(_04402_));
 sky130_fd_sc_hd__mux2_1 _11622_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_04189_),
    .X(_04403_));
 sky130_fd_sc_hd__mux2_1 _11623_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04188_),
    .X(_04404_));
 sky130_fd_sc_hd__or2_1 _11624_ (.A(_03652_),
    .B(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__o211a_1 _11625_ (.A1(_04192_),
    .A2(_04403_),
    .B1(_04405_),
    .C1(_04179_),
    .X(_04406_));
 sky130_fd_sc_hd__mux2_1 _11626_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_03617_),
    .X(_04407_));
 sky130_fd_sc_hd__mux2_1 _11627_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_03616_),
    .X(_04408_));
 sky130_fd_sc_hd__or2_1 _11628_ (.A(_03693_),
    .B(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__o211a_1 _11629_ (.A1(_03612_),
    .A2(_04407_),
    .B1(_04409_),
    .C1(_03689_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _11630_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_03616_),
    .X(_04411_));
 sky130_fd_sc_hd__mux2_1 _11631_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_03616_),
    .X(_04412_));
 sky130_fd_sc_hd__mux2_1 _11632_ (.A0(_04411_),
    .A1(_04412_),
    .S(_03656_),
    .X(_04413_));
 sky130_fd_sc_hd__a21o_1 _11633_ (.A1(_03674_),
    .A2(_04413_),
    .B1(_03704_),
    .X(_04414_));
 sky130_fd_sc_hd__o32a_1 _11634_ (.A1(_03679_),
    .A2(_04402_),
    .A3(_04406_),
    .B1(_04410_),
    .B2(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__mux2_1 _11635_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_03616_),
    .X(_04416_));
 sky130_fd_sc_hd__mux2_1 _11636_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_03616_),
    .X(_04417_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(_04416_),
    .A1(_04417_),
    .S(_03656_),
    .X(_04418_));
 sky130_fd_sc_hd__mux2_1 _11638_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_04376_),
    .X(_04419_));
 sky130_fd_sc_hd__and3_1 _11639_ (.A(\rbzero.tex_b1[59] ),
    .B(_03696_),
    .C(_03697_),
    .X(_04420_));
 sky130_fd_sc_hd__a21o_1 _11640_ (.A1(\rbzero.tex_b1[58] ),
    .A2(_03663_),
    .B1(_03823_),
    .X(_04421_));
 sky130_fd_sc_hd__o221a_1 _11641_ (.A1(_03693_),
    .A2(_04419_),
    .B1(_04420_),
    .B2(_04421_),
    .C1(_03673_),
    .X(_04422_));
 sky130_fd_sc_hd__a211o_1 _11642_ (.A1(_03689_),
    .A2(_04418_),
    .B1(_04422_),
    .C1(_03679_),
    .X(_04423_));
 sky130_fd_sc_hd__mux2_1 _11643_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04376_),
    .X(_04424_));
 sky130_fd_sc_hd__mux2_1 _11644_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04376_),
    .X(_04425_));
 sky130_fd_sc_hd__mux2_1 _11645_ (.A0(_04424_),
    .A1(_04425_),
    .S(_03739_),
    .X(_04426_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_03616_),
    .X(_04427_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_03615_),
    .X(_04428_));
 sky130_fd_sc_hd__or2_1 _11648_ (.A(_03823_),
    .B(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__o211a_1 _11649_ (.A1(_03693_),
    .A2(_04427_),
    .B1(_04429_),
    .C1(_03669_),
    .X(_04430_));
 sky130_fd_sc_hd__a211o_1 _11650_ (.A1(_03607_),
    .A2(_04426_),
    .B1(_04430_),
    .C1(_03704_),
    .X(_04431_));
 sky130_fd_sc_hd__a21o_1 _11651_ (.A1(_04423_),
    .A2(_04431_),
    .B1(_03685_),
    .X(_04432_));
 sky130_fd_sc_hd__o211a_1 _11652_ (.A1(_03688_),
    .A2(_04415_),
    .B1(_04432_),
    .C1(_03719_),
    .X(_04433_));
 sky130_fd_sc_hd__mux2_1 _11653_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_04376_),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_04376_),
    .X(_04435_));
 sky130_fd_sc_hd__mux2_1 _11655_ (.A0(_04434_),
    .A1(_04435_),
    .S(_03739_),
    .X(_04436_));
 sky130_fd_sc_hd__mux2_1 _11656_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_04376_),
    .X(_04437_));
 sky130_fd_sc_hd__and3_1 _11657_ (.A(\rbzero.tex_b1[27] ),
    .B(_03696_),
    .C(_03697_),
    .X(_04438_));
 sky130_fd_sc_hd__a21o_1 _11658_ (.A1(\rbzero.tex_b1[26] ),
    .A2(_03690_),
    .B1(_03823_),
    .X(_04439_));
 sky130_fd_sc_hd__o221a_1 _11659_ (.A1(_03656_),
    .A2(_04437_),
    .B1(_04438_),
    .B2(_04439_),
    .C1(_03673_),
    .X(_04440_));
 sky130_fd_sc_hd__a211o_1 _11660_ (.A1(_03689_),
    .A2(_04436_),
    .B1(_04440_),
    .C1(_03679_),
    .X(_04441_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04376_),
    .X(_04442_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_03699_),
    .X(_04443_));
 sky130_fd_sc_hd__mux2_1 _11663_ (.A0(_04442_),
    .A1(_04443_),
    .S(_03739_),
    .X(_04444_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_03616_),
    .X(_04445_));
 sky130_fd_sc_hd__mux2_1 _11665_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_03614_),
    .X(_04446_));
 sky130_fd_sc_hd__or2_1 _11666_ (.A(_03823_),
    .B(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__o211a_1 _11667_ (.A1(_03693_),
    .A2(_04445_),
    .B1(_04447_),
    .C1(_03669_),
    .X(_04448_));
 sky130_fd_sc_hd__a211o_1 _11668_ (.A1(_03607_),
    .A2(_04444_),
    .B1(_04448_),
    .C1(_03627_),
    .X(_04449_));
 sky130_fd_sc_hd__a21o_1 _11669_ (.A1(_04441_),
    .A2(_04449_),
    .B1(_03685_),
    .X(_04450_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04376_),
    .X(_04451_));
 sky130_fd_sc_hd__mux2_1 _11671_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04376_),
    .X(_04452_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(_04451_),
    .A1(_04452_),
    .S(_03739_),
    .X(_04453_));
 sky130_fd_sc_hd__mux2_1 _11673_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_03616_),
    .X(_04454_));
 sky130_fd_sc_hd__mux2_1 _11674_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_03615_),
    .X(_04455_));
 sky130_fd_sc_hd__or2_1 _11675_ (.A(_03823_),
    .B(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__o211a_1 _11676_ (.A1(_03693_),
    .A2(_04454_),
    .B1(_04456_),
    .C1(_03669_),
    .X(_04457_));
 sky130_fd_sc_hd__a211o_1 _11677_ (.A1(_03607_),
    .A2(_04453_),
    .B1(_04457_),
    .C1(_03624_),
    .X(_04458_));
 sky130_fd_sc_hd__mux2_1 _11678_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_03699_),
    .X(_04459_));
 sky130_fd_sc_hd__mux2_1 _11679_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_03699_),
    .X(_04460_));
 sky130_fd_sc_hd__mux2_1 _11680_ (.A0(_04459_),
    .A1(_04460_),
    .S(_03739_),
    .X(_04461_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_03699_),
    .X(_04462_));
 sky130_fd_sc_hd__and3_1 _11682_ (.A(\rbzero.tex_b1[3] ),
    .B(_03696_),
    .C(_03697_),
    .X(_04463_));
 sky130_fd_sc_hd__a21o_1 _11683_ (.A1(\rbzero.tex_b1[2] ),
    .A2(_03690_),
    .B1(_03823_),
    .X(_04464_));
 sky130_fd_sc_hd__o221a_1 _11684_ (.A1(_03656_),
    .A2(_04462_),
    .B1(_04463_),
    .B2(_04464_),
    .C1(_03673_),
    .X(_04465_));
 sky130_fd_sc_hd__a211o_1 _11685_ (.A1(_03689_),
    .A2(_04461_),
    .B1(_04465_),
    .C1(_03627_),
    .X(_04466_));
 sky130_fd_sc_hd__a21o_1 _11686_ (.A1(_04458_),
    .A2(_04466_),
    .B1(_03687_),
    .X(_04467_));
 sky130_fd_sc_hd__a31o_1 _11687_ (.A1(_03718_),
    .A2(_04450_),
    .A3(_04467_),
    .B1(_03537_),
    .X(_04468_));
 sky130_fd_sc_hd__o32a_1 _11688_ (.A1(_03764_),
    .A2(_04396_),
    .A3(_04398_),
    .B1(_04433_),
    .B2(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__mux2_1 _11689_ (.A0(_04394_),
    .A1(_04469_),
    .S(_03830_),
    .X(_04470_));
 sky130_fd_sc_hd__and2_1 _11690_ (.A(_03896_),
    .B(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__a31o_1 _11691_ (.A1(_03534_),
    .A2(_03848_),
    .A3(_04390_),
    .B1(_03522_),
    .X(_04472_));
 sky130_fd_sc_hd__o21a_1 _11692_ (.A1(_04471_),
    .A2(_04472_),
    .B1(_04148_),
    .X(_04473_));
 sky130_fd_sc_hd__buf_6 _11693_ (.A(_04473_),
    .X(net65));
 sky130_fd_sc_hd__nand4_1 _11694_ (.A(_03838_),
    .B(_03465_),
    .C(_04019_),
    .D(_03529_),
    .Y(_04474_));
 sky130_fd_sc_hd__a31o_1 _11695_ (.A1(_02899_),
    .A2(_04032_),
    .A3(_03528_),
    .B1(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__or3_1 _11696_ (.A(_04020_),
    .B(_03464_),
    .C(_03528_),
    .X(_04476_));
 sky130_fd_sc_hd__inv_2 _11697_ (.A(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(\rbzero.row_render.texu[1] ),
    .A1(\rbzero.row_render.texu[0] ),
    .S(_02899_),
    .X(_04478_));
 sky130_fd_sc_hd__mux4_1 _11699_ (.A0(\rbzero.row_render.texu[3] ),
    .A1(\rbzero.row_render.texu[2] ),
    .A2(_03539_),
    .A3(\rbzero.row_render.side ),
    .S0(_02899_),
    .S1(_03783_),
    .X(_04479_));
 sky130_fd_sc_hd__or2b_1 _11700_ (.A(\rbzero.row_render.texu[4] ),
    .B_N(_02899_),
    .X(_04480_));
 sky130_fd_sc_hd__o211a_1 _11701_ (.A1(\rbzero.row_render.texu[5] ),
    .A2(_02899_),
    .B1(_04480_),
    .C1(_03526_),
    .X(_04481_));
 sky130_fd_sc_hd__a311o_1 _11702_ (.A1(_03783_),
    .A2(_02899_),
    .A3(_04236_),
    .B1(_04481_),
    .C1(_03527_),
    .X(_04482_));
 sky130_fd_sc_hd__inv_2 _11703_ (.A(_03505_),
    .Y(_04483_));
 sky130_fd_sc_hd__o2111a_1 _11704_ (.A1(_03499_),
    .A2(_04479_),
    .B1(_04482_),
    .C1(_04020_),
    .D1(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__a21oi_1 _11705_ (.A1(_04477_),
    .A2(_04478_),
    .B1(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__o22ai_4 _11706_ (.A1(_03471_),
    .A2(_04475_),
    .B1(_04485_),
    .B2(net69),
    .Y(net70));
 sky130_fd_sc_hd__buf_1 _11707_ (.A(clknet_leaf_29_i_clk),
    .X(_04486_));
 sky130_fd_sc_hd__inv_2 _19253__3 (.A(clknet_1_0__leaf__02433_),
    .Y(net125));
 sky130_fd_sc_hd__buf_2 _11709_ (.A(net3),
    .X(_04487_));
 sky130_fd_sc_hd__nor2_1 _11710_ (.A(_04487_),
    .B(_03913_),
    .Y(_04488_));
 sky130_fd_sc_hd__a211o_1 _11711_ (.A1(_04487_),
    .A2(net67),
    .B1(_04488_),
    .C1(net7),
    .X(_04489_));
 sky130_fd_sc_hd__nand2_1 _11712_ (.A(_04487_),
    .B(_04314_),
    .Y(_04490_));
 sky130_fd_sc_hd__or2_1 _11713_ (.A(_04487_),
    .B(net62),
    .X(_04491_));
 sky130_fd_sc_hd__a31o_1 _11714_ (.A1(net7),
    .A2(_04490_),
    .A3(_04491_),
    .B1(net6),
    .X(_04492_));
 sky130_fd_sc_hd__nor2_1 _11715_ (.A(_04487_),
    .B(_04393_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2_1 _11716_ (.A(net6),
    .B(net7),
    .Y(_04494_));
 sky130_fd_sc_hd__a211o_1 _11717_ (.A1(_04487_),
    .A2(net65),
    .B1(_04493_),
    .C1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__buf_2 _11718_ (.A(net5),
    .X(_04496_));
 sky130_fd_sc_hd__and4b_1 _11719_ (.A_N(net8),
    .B(_04495_),
    .C(net4),
    .D(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__and3_1 _11720_ (.A(_04489_),
    .B(_04492_),
    .C(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__buf_2 _11721_ (.A(\gpout0.vpos[0] ),
    .X(_04499_));
 sky130_fd_sc_hd__buf_2 _11722_ (.A(\gpout0.vpos[1] ),
    .X(_04500_));
 sky130_fd_sc_hd__mux4_1 _11723_ (.A0(_03906_),
    .A1(_04499_),
    .A2(_03909_),
    .A3(_04500_),
    .S0(_04494_),
    .S1(_04487_),
    .X(_04501_));
 sky130_fd_sc_hd__nand2_1 _11724_ (.A(_04496_),
    .B(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__clkbuf_4 _11725_ (.A(_03834_),
    .X(_04503_));
 sky130_fd_sc_hd__nor2_1 _11726_ (.A(_04503_),
    .B(_04487_),
    .Y(_04504_));
 sky130_fd_sc_hd__a211o_1 _11727_ (.A1(_03852_),
    .A2(_04487_),
    .B1(_04496_),
    .C1(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__nand3_1 _11728_ (.A(net4),
    .B(_04502_),
    .C(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__clkbuf_4 _11729_ (.A(\gpout0.vpos[2] ),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_4 _11730_ (.A(_03517_),
    .X(_04508_));
 sky130_fd_sc_hd__mux4_1 _11731_ (.A0(_04507_),
    .A1(_04508_),
    .A2(_03520_),
    .A3(_03515_),
    .S0(_04487_),
    .S1(_04496_),
    .X(_04509_));
 sky130_fd_sc_hd__a21o_1 _11732_ (.A1(net4),
    .A2(_04496_),
    .B1(net6),
    .X(_04510_));
 sky130_fd_sc_hd__o2111a_1 _11733_ (.A1(net4),
    .A2(_04509_),
    .B1(_04510_),
    .C1(net7),
    .D1(net8),
    .X(_04511_));
 sky130_fd_sc_hd__nor2_1 _11734_ (.A(net4),
    .B(net3),
    .Y(_04512_));
 sky130_fd_sc_hd__nor2_2 _11735_ (.A(net6),
    .B(_04496_),
    .Y(_04513_));
 sky130_fd_sc_hd__and2_1 _11736_ (.A(_04512_),
    .B(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__and2_1 _11737_ (.A(net4),
    .B(net3),
    .X(_04515_));
 sky130_fd_sc_hd__and2b_1 _11738_ (.A_N(net3),
    .B(net4),
    .X(_04516_));
 sky130_fd_sc_hd__and3_2 _11739_ (.A(clknet_leaf_31_i_clk),
    .B(_04516_),
    .C(_04513_),
    .X(_04517_));
 sky130_fd_sc_hd__a31o_2 _11740_ (.A1(\gpout0.clk_div[1] ),
    .A2(_04515_),
    .A3(_04513_),
    .B1(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__and2b_1 _11741_ (.A_N(net4),
    .B(net3),
    .X(_04519_));
 sky130_fd_sc_hd__a22o_1 _11742_ (.A1(net51),
    .A2(_04519_),
    .B1(_04516_),
    .B2(net53),
    .X(_04520_));
 sky130_fd_sc_hd__a21o_1 _11743_ (.A1(net50),
    .A2(_04512_),
    .B1(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__and2b_1 _11744_ (.A_N(net6),
    .B(net5),
    .X(_04522_));
 sky130_fd_sc_hd__a32o_1 _11745_ (.A1(_02981_),
    .A2(_04519_),
    .A3(_04513_),
    .B1(_04521_),
    .B2(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__or3_2 _11746_ (.A(_04514_),
    .B(_04518_),
    .C(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__nor2_1 _11747_ (.A(net8),
    .B(net7),
    .Y(_04525_));
 sky130_fd_sc_hd__a22o_2 _11748_ (.A1(_04506_),
    .A2(_04511_),
    .B1(_04524_),
    .B2(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__inv_2 _11749_ (.A(net7),
    .Y(_04527_));
 sky130_fd_sc_hd__a22o_1 _11750_ (.A1(_03910_),
    .A2(_04512_),
    .B1(_04519_),
    .B2(net69),
    .X(_04528_));
 sky130_fd_sc_hd__a22o_1 _11751_ (.A1(net49),
    .A2(_04512_),
    .B1(_04519_),
    .B2(net39),
    .X(_04529_));
 sky130_fd_sc_hd__a221o_1 _11752_ (.A1(_03537_),
    .A2(_04515_),
    .B1(_04516_),
    .B2(net40),
    .C1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__and3b_1 _11753_ (.A_N(_04496_),
    .B(_04530_),
    .C(net6),
    .X(_04531_));
 sky130_fd_sc_hd__buf_4 _11754_ (.A(net52),
    .X(_04532_));
 sky130_fd_sc_hd__and4_1 _11755_ (.A(_04532_),
    .B(_04522_),
    .C(_04515_),
    .D(_04525_),
    .X(_04533_));
 sky130_fd_sc_hd__a31o_1 _11756_ (.A1(net44),
    .A2(_04519_),
    .A3(_04513_),
    .B1(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__a22o_1 _11757_ (.A1(net48),
    .A2(_04515_),
    .B1(_04516_),
    .B2(net47),
    .X(_04535_));
 sky130_fd_sc_hd__and3_1 _11758_ (.A(net43),
    .B(_04516_),
    .C(_04513_),
    .X(_04536_));
 sky130_fd_sc_hd__a221o_1 _11759_ (.A1(_04522_),
    .A2(_04535_),
    .B1(_04514_),
    .B2(net42),
    .C1(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__a311o_1 _11760_ (.A1(_03911_),
    .A2(_04515_),
    .A3(_04513_),
    .B1(_04534_),
    .C1(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__a211o_1 _11761_ (.A1(_04522_),
    .A2(_04528_),
    .B1(_04531_),
    .C1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__a22o_1 _11762_ (.A1(_03782_),
    .A2(_04519_),
    .B1(_04515_),
    .B2(_03865_),
    .X(_04540_));
 sky130_fd_sc_hd__a221o_1 _11763_ (.A1(_03464_),
    .A2(_04512_),
    .B1(_04516_),
    .B2(_03474_),
    .C1(_04496_),
    .X(_04541_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(_03459_),
    .A1(_03469_),
    .S(net3),
    .X(_04542_));
 sky130_fd_sc_hd__mux4_1 _11765_ (.A0(\gpout0.hpos[0] ),
    .A1(_03527_),
    .A2(_03526_),
    .A3(_04020_),
    .S0(net3),
    .S1(net4),
    .X(_04543_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(_04542_),
    .A1(_04543_),
    .S(net6),
    .X(_04544_));
 sky130_fd_sc_hd__nand2_1 _11767_ (.A(_04496_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__o21ai_1 _11768_ (.A1(_04540_),
    .A2(_04541_),
    .B1(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__nand2_1 _11769_ (.A(net7),
    .B(_04510_),
    .Y(_04547_));
 sky130_fd_sc_hd__a21o_1 _11770_ (.A1(net6),
    .A2(_04496_),
    .B1(net7),
    .X(_04548_));
 sky130_fd_sc_hd__and4_1 _11771_ (.A(net8),
    .B(_04546_),
    .C(_04547_),
    .D(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__a311o_1 _11772_ (.A1(net8),
    .A2(_04527_),
    .A3(_04539_),
    .B1(_04549_),
    .C1(_04533_),
    .X(_04550_));
 sky130_fd_sc_hd__or4b_1 _11773_ (.A(net8),
    .B(net7),
    .C(net62),
    .D_N(_04514_),
    .X(_04551_));
 sky130_fd_sc_hd__o31a_2 _11774_ (.A1(_04498_),
    .A2(_04526_),
    .A3(_04550_),
    .B1(_04551_),
    .X(net54));
 sky130_fd_sc_hd__buf_2 _11775_ (.A(net15),
    .X(_04552_));
 sky130_fd_sc_hd__nor2_1 _11776_ (.A(_04552_),
    .B(_03913_),
    .Y(_04553_));
 sky130_fd_sc_hd__a211o_1 _11777_ (.A1(_04552_),
    .A2(net67),
    .B1(_04553_),
    .C1(net19),
    .X(_04554_));
 sky130_fd_sc_hd__nand2_1 _11778_ (.A(_04552_),
    .B(_04314_),
    .Y(_04555_));
 sky130_fd_sc_hd__or2_1 _11779_ (.A(_04552_),
    .B(net62),
    .X(_04556_));
 sky130_fd_sc_hd__a31o_1 _11780_ (.A1(net19),
    .A2(_04555_),
    .A3(_04556_),
    .B1(net18),
    .X(_04557_));
 sky130_fd_sc_hd__nor2_1 _11781_ (.A(_04552_),
    .B(_04393_),
    .Y(_04558_));
 sky130_fd_sc_hd__nand2_1 _11782_ (.A(net18),
    .B(net19),
    .Y(_04559_));
 sky130_fd_sc_hd__a211o_1 _11783_ (.A1(_04552_),
    .A2(net65),
    .B1(_04558_),
    .C1(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__and4b_1 _11784_ (.A_N(net20),
    .B(_04560_),
    .C(net16),
    .D(net17),
    .X(_04561_));
 sky130_fd_sc_hd__and3_1 _11785_ (.A(_04554_),
    .B(_04557_),
    .C(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__inv_2 _11786_ (.A(net19),
    .Y(_04563_));
 sky130_fd_sc_hd__inv_2 _11787_ (.A(net17),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_1 _11788_ (.A(net18),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__nor2_1 _11789_ (.A(net16),
    .B(net15),
    .Y(_04566_));
 sky130_fd_sc_hd__inv_2 _11790_ (.A(net16),
    .Y(_04567_));
 sky130_fd_sc_hd__and2_1 _11791_ (.A(_04567_),
    .B(net15),
    .X(_04568_));
 sky130_fd_sc_hd__nor2_2 _11792_ (.A(_04567_),
    .B(net15),
    .Y(_04569_));
 sky130_fd_sc_hd__and2_1 _11793_ (.A(net16),
    .B(net15),
    .X(_04570_));
 sky130_fd_sc_hd__nor2_1 _11794_ (.A(net20),
    .B(net19),
    .Y(_04571_));
 sky130_fd_sc_hd__a21o_1 _11795_ (.A1(_04532_),
    .A2(_04571_),
    .B1(net48),
    .X(_04572_));
 sky130_fd_sc_hd__a22o_1 _11796_ (.A1(net47),
    .A2(_04569_),
    .B1(_04570_),
    .B2(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__a221o_1 _11797_ (.A1(_03910_),
    .A2(_04566_),
    .B1(_04568_),
    .B2(net69),
    .C1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__a22o_1 _11798_ (.A1(net49),
    .A2(_04566_),
    .B1(_04568_),
    .B2(net39),
    .X(_04575_));
 sky130_fd_sc_hd__a221o_1 _11799_ (.A1(net40),
    .A2(_04569_),
    .B1(_04570_),
    .B2(_03537_),
    .C1(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__nor2_2 _11800_ (.A(net18),
    .B(net17),
    .Y(_04577_));
 sky130_fd_sc_hd__and3_1 _11801_ (.A(net43),
    .B(_04569_),
    .C(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__and2_1 _11802_ (.A(_04566_),
    .B(_04577_),
    .X(_04579_));
 sky130_fd_sc_hd__a32o_1 _11803_ (.A1(_03911_),
    .A2(_04577_),
    .A3(_04570_),
    .B1(_04579_),
    .B2(net42),
    .X(_04580_));
 sky130_fd_sc_hd__a311o_1 _11804_ (.A1(net44),
    .A2(_04568_),
    .A3(_04577_),
    .B1(_04578_),
    .C1(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__a31o_1 _11805_ (.A1(net18),
    .A2(_04564_),
    .A3(_04576_),
    .B1(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__a21o_1 _11806_ (.A1(_04565_),
    .A2(_04574_),
    .B1(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__a21o_1 _11807_ (.A1(net16),
    .A2(net17),
    .B1(net18),
    .X(_04584_));
 sky130_fd_sc_hd__nand2_1 _11808_ (.A(net19),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(_03459_),
    .A1(_03469_),
    .S(net15),
    .X(_04586_));
 sky130_fd_sc_hd__mux4_1 _11810_ (.A0(\gpout0.hpos[0] ),
    .A1(_03527_),
    .A2(_03526_),
    .A3(_04020_),
    .S0(net15),
    .S1(net16),
    .X(_04587_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(_04586_),
    .A1(_04587_),
    .S(net18),
    .X(_04588_));
 sky130_fd_sc_hd__a22o_1 _11812_ (.A1(_03782_),
    .A2(_04568_),
    .B1(_04570_),
    .B2(_03865_),
    .X(_04589_));
 sky130_fd_sc_hd__a211o_1 _11813_ (.A1(_03474_),
    .A2(_04569_),
    .B1(_04589_),
    .C1(net17),
    .X(_04590_));
 sky130_fd_sc_hd__a21oi_1 _11814_ (.A1(_03464_),
    .A2(_04566_),
    .B1(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a21o_1 _11815_ (.A1(net17),
    .A2(_04588_),
    .B1(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__a21o_1 _11816_ (.A1(net18),
    .A2(net17),
    .B1(net19),
    .X(_04593_));
 sky130_fd_sc_hd__and4_1 _11817_ (.A(net20),
    .B(_04585_),
    .C(_04592_),
    .D(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__a41o_1 _11818_ (.A1(_04532_),
    .A2(_04571_),
    .A3(_04565_),
    .A4(_04570_),
    .B1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__and3_1 _11819_ (.A(\gpout2.clk_div[1] ),
    .B(_04577_),
    .C(_04570_),
    .X(_04596_));
 sky130_fd_sc_hd__a31o_1 _11820_ (.A1(net45),
    .A2(_04568_),
    .A3(_04577_),
    .B1(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__and2_1 _11821_ (.A(net50),
    .B(_04566_),
    .X(_04598_));
 sky130_fd_sc_hd__a221o_1 _11822_ (.A1(net53),
    .A2(_04569_),
    .B1(_04568_),
    .B2(net51),
    .C1(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__a32o_2 _11823_ (.A1(clknet_1_0__leaf__04486_),
    .A2(_04569_),
    .A3(_04577_),
    .B1(_04565_),
    .B2(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__o31a_2 _11824_ (.A1(_04579_),
    .A2(_04597_),
    .A3(_04600_),
    .B1(_04571_),
    .X(_04601_));
 sky130_fd_sc_hd__mux4_1 _11825_ (.A0(_03906_),
    .A1(_04499_),
    .A2(_03909_),
    .A3(\gpout0.vpos[1] ),
    .S0(_04559_),
    .S1(_04552_),
    .X(_04602_));
 sky130_fd_sc_hd__nand2_1 _11826_ (.A(net17),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__nor2_1 _11827_ (.A(_04503_),
    .B(_04552_),
    .Y(_04604_));
 sky130_fd_sc_hd__a211o_1 _11828_ (.A1(_03852_),
    .A2(_04552_),
    .B1(net17),
    .C1(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__mux4_1 _11829_ (.A0(_04507_),
    .A1(_04508_),
    .A2(_03520_),
    .A3(_03515_),
    .S0(_04552_),
    .S1(net17),
    .X(_04606_));
 sky130_fd_sc_hd__o2111ai_1 _11830_ (.A1(net16),
    .A2(_04606_),
    .B1(_04584_),
    .C1(net20),
    .D1(net19),
    .Y(_04607_));
 sky130_fd_sc_hd__a31o_1 _11831_ (.A1(net16),
    .A2(_04603_),
    .A3(_04605_),
    .B1(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__or3b_2 _11832_ (.A(_04595_),
    .B(_04601_),
    .C_N(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__a31o_2 _11833_ (.A1(net20),
    .A2(_04563_),
    .A3(_04583_),
    .B1(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__nand2_1 _11834_ (.A(_04571_),
    .B(_04579_),
    .Y(_04611_));
 sky130_fd_sc_hd__o22a_2 _11835_ (.A1(_04562_),
    .A2(_04610_),
    .B1(_04611_),
    .B2(net66),
    .X(net56));
 sky130_fd_sc_hd__buf_2 _11836_ (.A(net9),
    .X(_04612_));
 sky130_fd_sc_hd__nand2_1 _11837_ (.A(_04612_),
    .B(_04314_),
    .Y(_04613_));
 sky130_fd_sc_hd__o211a_1 _11838_ (.A1(_04612_),
    .A2(net62),
    .B1(_04613_),
    .C1(net13),
    .X(_04614_));
 sky130_fd_sc_hd__nor2_1 _11839_ (.A(_04612_),
    .B(_04393_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand2_1 _11840_ (.A(net12),
    .B(net13),
    .Y(_04616_));
 sky130_fd_sc_hd__a211o_1 _11841_ (.A1(_04612_),
    .A2(net65),
    .B1(_04615_),
    .C1(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__and4b_1 _11842_ (.A_N(net14),
    .B(_04617_),
    .C(net10),
    .D(net11),
    .X(_04618_));
 sky130_fd_sc_hd__nor2_1 _11843_ (.A(_04612_),
    .B(_03913_),
    .Y(_04619_));
 sky130_fd_sc_hd__a211o_1 _11844_ (.A1(_04612_),
    .A2(net67),
    .B1(_04619_),
    .C1(net13),
    .X(_04620_));
 sky130_fd_sc_hd__o211a_1 _11845_ (.A1(net12),
    .A2(_04614_),
    .B1(_04618_),
    .C1(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__nor2_1 _11846_ (.A(net10),
    .B(net9),
    .Y(_04622_));
 sky130_fd_sc_hd__nor2_1 _11847_ (.A(net12),
    .B(net11),
    .Y(_04623_));
 sky130_fd_sc_hd__inv_2 _11848_ (.A(net11),
    .Y(_04624_));
 sky130_fd_sc_hd__and2b_1 _11849_ (.A_N(net10),
    .B(net9),
    .X(_04625_));
 sky130_fd_sc_hd__and2b_1 _11850_ (.A_N(net9),
    .B(net10),
    .X(_04626_));
 sky130_fd_sc_hd__and2_1 _11851_ (.A(net10),
    .B(net9),
    .X(_04627_));
 sky130_fd_sc_hd__a22o_1 _11852_ (.A1(net40),
    .A2(_04626_),
    .B1(_04627_),
    .B2(_03537_),
    .X(_04628_));
 sky130_fd_sc_hd__a221o_1 _11853_ (.A1(net49),
    .A2(_04622_),
    .B1(_04625_),
    .B2(net39),
    .C1(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__and3_1 _11854_ (.A(net12),
    .B(_04624_),
    .C(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__a31o_1 _11855_ (.A1(net42),
    .A2(_04622_),
    .A3(_04623_),
    .B1(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__nor2_1 _11856_ (.A(net14),
    .B(net13),
    .Y(_04632_));
 sky130_fd_sc_hd__a21o_1 _11857_ (.A1(_04532_),
    .A2(_04632_),
    .B1(net48),
    .X(_04633_));
 sky130_fd_sc_hd__a22o_1 _11858_ (.A1(net47),
    .A2(_04626_),
    .B1(_04627_),
    .B2(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__nor2_2 _11859_ (.A(net12),
    .B(_04624_),
    .Y(_04635_));
 sky130_fd_sc_hd__a32o_1 _11860_ (.A1(net44),
    .A2(_04625_),
    .A3(_04623_),
    .B1(_04634_),
    .B2(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__a31o_1 _11861_ (.A1(_04532_),
    .A2(_04635_),
    .A3(_04627_),
    .B1(net14),
    .X(_04637_));
 sky130_fd_sc_hd__o21ai_1 _11862_ (.A1(_04631_),
    .A2(_04636_),
    .B1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand2_2 _11863_ (.A(net124),
    .B(_04626_),
    .Y(_04639_));
 sky130_fd_sc_hd__or2b_1 _11864_ (.A(\gpout1.clk_div[1] ),
    .B_N(_04627_),
    .X(_04640_));
 sky130_fd_sc_hd__a22o_1 _11865_ (.A1(net51),
    .A2(_04625_),
    .B1(_04626_),
    .B2(net53),
    .X(_04641_));
 sky130_fd_sc_hd__a21o_1 _11866_ (.A1(net50),
    .A2(_04622_),
    .B1(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__a32o_2 _11867_ (.A1(_04639_),
    .A2(_04623_),
    .A3(_04640_),
    .B1(_04635_),
    .B2(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__a2bb2o_2 _11868_ (.A1_N(net13),
    .A2_N(_04638_),
    .B1(_04643_),
    .B2(_04632_),
    .X(_04644_));
 sky130_fd_sc_hd__a21o_1 _11869_ (.A1(net10),
    .A2(net11),
    .B1(net12),
    .X(_04645_));
 sky130_fd_sc_hd__mux4_1 _11870_ (.A0(\gpout0.hpos[0] ),
    .A1(_03527_),
    .A2(_03526_),
    .A3(_04020_),
    .S0(net9),
    .S1(net10),
    .X(_04646_));
 sky130_fd_sc_hd__and3_1 _11871_ (.A(net12),
    .B(net11),
    .C(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__mux4_1 _11872_ (.A0(_03524_),
    .A1(_03461_),
    .A2(_03838_),
    .A3(_02901_),
    .S0(net9),
    .S1(net10),
    .X(_04648_));
 sky130_fd_sc_hd__mux2_1 _11873_ (.A0(_03459_),
    .A1(_03469_),
    .S(_04612_),
    .X(_04649_));
 sky130_fd_sc_hd__a22o_1 _11874_ (.A1(_04624_),
    .A2(_04648_),
    .B1(_04649_),
    .B2(_04635_),
    .X(_04650_));
 sky130_fd_sc_hd__nor2_1 _11875_ (.A(_04647_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(_04503_),
    .A1(_03902_),
    .S(_04612_),
    .X(_04652_));
 sky130_fd_sc_hd__mux4_1 _11877_ (.A0(_03906_),
    .A1(_04499_),
    .A2(_03909_),
    .A3(_04500_),
    .S0(_04616_),
    .S1(_04612_),
    .X(_04653_));
 sky130_fd_sc_hd__a21bo_1 _11878_ (.A1(net11),
    .A2(_04653_),
    .B1_N(net10),
    .X(_04654_));
 sky130_fd_sc_hd__a21oi_1 _11879_ (.A1(_04624_),
    .A2(_04652_),
    .B1(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__mux4_1 _11880_ (.A0(_04507_),
    .A1(_04508_),
    .A2(_03520_),
    .A3(_03515_),
    .S0(_04612_),
    .S1(net11),
    .X(_04656_));
 sky130_fd_sc_hd__o21ai_1 _11881_ (.A1(net10),
    .A2(_04656_),
    .B1(_04645_),
    .Y(_04657_));
 sky130_fd_sc_hd__o221a_1 _11882_ (.A1(_04645_),
    .A2(_04651_),
    .B1(_04655_),
    .B2(_04657_),
    .C1(net13),
    .X(_04658_));
 sky130_fd_sc_hd__a22o_1 _11883_ (.A1(_03910_),
    .A2(_04622_),
    .B1(_04625_),
    .B2(net69),
    .X(_04659_));
 sky130_fd_sc_hd__a22o_1 _11884_ (.A1(net43),
    .A2(_04626_),
    .B1(_04627_),
    .B2(_03911_),
    .X(_04660_));
 sky130_fd_sc_hd__a211o_1 _11885_ (.A1(_04623_),
    .A2(_04660_),
    .B1(_04647_),
    .C1(net13),
    .X(_04661_));
 sky130_fd_sc_hd__a21o_1 _11886_ (.A1(_04635_),
    .A2(_04659_),
    .B1(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__and3b_1 _11887_ (.A_N(_04658_),
    .B(net14),
    .C(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__nand4_1 _11888_ (.A(_04314_),
    .B(_04622_),
    .C(_04623_),
    .D(_04632_),
    .Y(_04664_));
 sky130_fd_sc_hd__o31a_2 _11889_ (.A1(_04621_),
    .A2(_04644_),
    .A3(_04663_),
    .B1(_04664_),
    .X(net55));
 sky130_fd_sc_hd__and2b_1 _11890_ (.A_N(net22),
    .B(net21),
    .X(_04665_));
 sky130_fd_sc_hd__and2_1 _11891_ (.A(net22),
    .B(net21),
    .X(_04666_));
 sky130_fd_sc_hd__a22o_1 _11892_ (.A1(_03782_),
    .A2(_04665_),
    .B1(_04666_),
    .B2(_03865_),
    .X(_04667_));
 sky130_fd_sc_hd__and2b_1 _11893_ (.A_N(net21),
    .B(net22),
    .X(_04668_));
 sky130_fd_sc_hd__nor2_1 _11894_ (.A(net22),
    .B(net21),
    .Y(_04669_));
 sky130_fd_sc_hd__buf_2 _11895_ (.A(net23),
    .X(_04670_));
 sky130_fd_sc_hd__a221o_1 _11896_ (.A1(_03474_),
    .A2(_04668_),
    .B1(_04669_),
    .B2(_03464_),
    .C1(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__buf_2 _11897_ (.A(net21),
    .X(_04672_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(_03459_),
    .A1(_03469_),
    .S(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__mux4_1 _11899_ (.A0(_02899_),
    .A1(_03527_),
    .A2(_03526_),
    .A3(_04020_),
    .S0(net21),
    .S1(net22),
    .X(_04674_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(_04673_),
    .A1(_04674_),
    .S(net24),
    .X(_04675_));
 sky130_fd_sc_hd__nand2_1 _11901_ (.A(_04670_),
    .B(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__o21a_1 _11902_ (.A1(_04667_),
    .A2(_04671_),
    .B1(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__a21o_1 _11903_ (.A1(net22),
    .A2(_04670_),
    .B1(net24),
    .X(_04678_));
 sky130_fd_sc_hd__a21oi_1 _11904_ (.A1(net24),
    .A2(_04670_),
    .B1(net25),
    .Y(_04679_));
 sky130_fd_sc_hd__inv_2 _11905_ (.A(net26),
    .Y(_04680_));
 sky130_fd_sc_hd__a211o_1 _11906_ (.A1(net25),
    .A2(_04678_),
    .B1(_04679_),
    .C1(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__and2b_1 _11907_ (.A_N(net24),
    .B(_04670_),
    .X(_04682_));
 sky130_fd_sc_hd__a22o_1 _11908_ (.A1(net51),
    .A2(_04665_),
    .B1(_04669_),
    .B2(net50),
    .X(_04683_));
 sky130_fd_sc_hd__a221o_1 _11909_ (.A1(_04532_),
    .A2(_04666_),
    .B1(_04668_),
    .B2(net53),
    .C1(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__nor2_2 _11910_ (.A(net24),
    .B(net23),
    .Y(_04685_));
 sky130_fd_sc_hd__and2_1 _11911_ (.A(_04669_),
    .B(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__and3_1 _11912_ (.A(net46),
    .B(_04665_),
    .C(_04685_),
    .X(_04687_));
 sky130_fd_sc_hd__a31o_1 _11913_ (.A1(\gpout3.clk_div[1] ),
    .A2(_04666_),
    .A3(_04685_),
    .B1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__a311o_2 _11914_ (.A1(clknet_1_0__leaf__04486_),
    .A2(_04668_),
    .A3(_04685_),
    .B1(_04686_),
    .C1(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__a21oi_2 _11915_ (.A1(_04682_),
    .A2(_04684_),
    .B1(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2_1 _11916_ (.A(net24),
    .B(net25),
    .Y(_04691_));
 sky130_fd_sc_hd__mux4_1 _11917_ (.A0(_03906_),
    .A1(_04499_),
    .A2(_03909_),
    .A3(_04500_),
    .S0(_04691_),
    .S1(_04672_),
    .X(_04692_));
 sky130_fd_sc_hd__nand2_1 _11918_ (.A(_04670_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__nor2_1 _11919_ (.A(_04503_),
    .B(_04672_),
    .Y(_04694_));
 sky130_fd_sc_hd__a211o_1 _11920_ (.A1(_03852_),
    .A2(_04672_),
    .B1(_04670_),
    .C1(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__mux4_1 _11921_ (.A0(_04507_),
    .A1(_04508_),
    .A2(_03520_),
    .A3(_03515_),
    .S0(net21),
    .S1(_04670_),
    .X(_04696_));
 sky130_fd_sc_hd__o2111ai_1 _11922_ (.A1(net22),
    .A2(_04696_),
    .B1(_04678_),
    .C1(net26),
    .D1(net25),
    .Y(_04697_));
 sky130_fd_sc_hd__a31o_1 _11923_ (.A1(net22),
    .A2(_04693_),
    .A3(_04695_),
    .B1(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__o31a_2 _11924_ (.A1(net25),
    .A2(net26),
    .A3(_04690_),
    .B1(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__o21ai_2 _11925_ (.A1(_04677_),
    .A2(_04681_),
    .B1(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__nand2_1 _11926_ (.A(_04672_),
    .B(_04314_),
    .Y(_04701_));
 sky130_fd_sc_hd__or2_1 _11927_ (.A(_04672_),
    .B(net62),
    .X(_04702_));
 sky130_fd_sc_hd__a31o_1 _11928_ (.A1(net25),
    .A2(_04701_),
    .A3(_04702_),
    .B1(net24),
    .X(_04703_));
 sky130_fd_sc_hd__nor2_1 _11929_ (.A(_04672_),
    .B(_04393_),
    .Y(_04704_));
 sky130_fd_sc_hd__a211o_1 _11930_ (.A1(_04672_),
    .A2(net65),
    .B1(_04704_),
    .C1(_04691_),
    .X(_04705_));
 sky130_fd_sc_hd__nor2_1 _11931_ (.A(_04672_),
    .B(_03913_),
    .Y(_04706_));
 sky130_fd_sc_hd__a211o_1 _11932_ (.A1(_04672_),
    .A2(net67),
    .B1(_04706_),
    .C1(net25),
    .X(_04707_));
 sky130_fd_sc_hd__and4_1 _11933_ (.A(net22),
    .B(_04670_),
    .C(_04680_),
    .D(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__inv_2 _11934_ (.A(net25),
    .Y(_04709_));
 sky130_fd_sc_hd__a31o_1 _11935_ (.A1(_04532_),
    .A2(_04709_),
    .A3(_04680_),
    .B1(net48),
    .X(_04710_));
 sky130_fd_sc_hd__a22o_1 _11936_ (.A1(net47),
    .A2(_04668_),
    .B1(_04710_),
    .B2(_04666_),
    .X(_04711_));
 sky130_fd_sc_hd__a221o_1 _11937_ (.A1(net69),
    .A2(_04665_),
    .B1(_04669_),
    .B2(_03910_),
    .C1(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__a22o_1 _11938_ (.A1(net39),
    .A2(_04665_),
    .B1(_04669_),
    .B2(net49),
    .X(_04713_));
 sky130_fd_sc_hd__a221o_1 _11939_ (.A1(_03537_),
    .A2(_04666_),
    .B1(_04668_),
    .B2(net40),
    .C1(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__and3b_1 _11940_ (.A_N(_04670_),
    .B(_04714_),
    .C(net24),
    .X(_04715_));
 sky130_fd_sc_hd__a32o_1 _11941_ (.A1(_03911_),
    .A2(_04666_),
    .A3(_04685_),
    .B1(_04686_),
    .B2(net42),
    .X(_04716_));
 sky130_fd_sc_hd__and3_1 _11942_ (.A(net44),
    .B(_04665_),
    .C(_04685_),
    .X(_04717_));
 sky130_fd_sc_hd__a311o_1 _11943_ (.A1(net43),
    .A2(_04668_),
    .A3(_04685_),
    .B1(_04716_),
    .C1(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__a211o_1 _11944_ (.A1(_04682_),
    .A2(_04712_),
    .B1(_04715_),
    .C1(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__and3b_1 _11945_ (.A_N(net25),
    .B(net26),
    .C(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__a31o_1 _11946_ (.A1(_04703_),
    .A2(_04705_),
    .A3(_04708_),
    .B1(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__or4b_1 _11947_ (.A(net25),
    .B(net26),
    .C(net67),
    .D_N(_04686_),
    .X(_04722_));
 sky130_fd_sc_hd__o21a_2 _11948_ (.A1(_04700_),
    .A2(_04721_),
    .B1(_04722_),
    .X(net57));
 sky130_fd_sc_hd__nor2_1 _11949_ (.A(net31),
    .B(net32),
    .Y(_04723_));
 sky130_fd_sc_hd__nor2_1 _11950_ (.A(net28),
    .B(net27),
    .Y(_04724_));
 sky130_fd_sc_hd__nor2_2 _11951_ (.A(net30),
    .B(net29),
    .Y(_04725_));
 sky130_fd_sc_hd__and2_1 _11952_ (.A(_04724_),
    .B(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(_03459_),
    .A1(_03469_),
    .S(net27),
    .X(_04727_));
 sky130_fd_sc_hd__mux4_1 _11954_ (.A0(\gpout0.hpos[0] ),
    .A1(_03527_),
    .A2(_03526_),
    .A3(_04020_),
    .S0(net27),
    .S1(net28),
    .X(_04728_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(_04727_),
    .A1(_04728_),
    .S(net30),
    .X(_04729_));
 sky130_fd_sc_hd__nor2b_2 _11956_ (.A(net27),
    .B_N(net28),
    .Y(_04730_));
 sky130_fd_sc_hd__and2b_1 _11957_ (.A_N(net28),
    .B(net27),
    .X(_04731_));
 sky130_fd_sc_hd__and2_1 _11958_ (.A(net28),
    .B(net27),
    .X(_04732_));
 sky130_fd_sc_hd__and2_1 _11959_ (.A(_03464_),
    .B(_04724_),
    .X(_04733_));
 sky130_fd_sc_hd__a221o_1 _11960_ (.A1(_03782_),
    .A2(_04731_),
    .B1(_04732_),
    .B2(_03865_),
    .C1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__a211oi_1 _11961_ (.A1(_03474_),
    .A2(_04730_),
    .B1(_04734_),
    .C1(net29),
    .Y(_04735_));
 sky130_fd_sc_hd__a21oi_1 _11962_ (.A1(net29),
    .A2(_04729_),
    .B1(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__nand2_1 _11963_ (.A(net30),
    .B(net31),
    .Y(_04737_));
 sky130_fd_sc_hd__inv_2 _11964_ (.A(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__a31o_1 _11965_ (.A1(net28),
    .A2(net29),
    .A3(net31),
    .B1(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__a21oi_1 _11966_ (.A1(net30),
    .A2(net29),
    .B1(net31),
    .Y(_04740_));
 sky130_fd_sc_hd__or4b_1 _11967_ (.A(_04736_),
    .B(_04739_),
    .C(_04740_),
    .D_N(net32),
    .X(_04741_));
 sky130_fd_sc_hd__inv_2 _11968_ (.A(net29),
    .Y(_04742_));
 sky130_fd_sc_hd__nor2_1 _11969_ (.A(net30),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__a22o_1 _11970_ (.A1(net53),
    .A2(_04730_),
    .B1(_04724_),
    .B2(net50),
    .X(_04744_));
 sky130_fd_sc_hd__a221o_1 _11971_ (.A1(net51),
    .A2(_04731_),
    .B1(_04732_),
    .B2(_04532_),
    .C1(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__and3_1 _11972_ (.A(net2),
    .B(_04731_),
    .C(_04725_),
    .X(_04746_));
 sky130_fd_sc_hd__a31o_1 _11973_ (.A1(\gpout4.clk_div[1] ),
    .A2(_04732_),
    .A3(_04725_),
    .B1(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__a31o_2 _11974_ (.A1(clknet_1_0__leaf__04486_),
    .A2(_04730_),
    .A3(_04725_),
    .B1(_04726_),
    .X(_04748_));
 sky130_fd_sc_hd__a211o_2 _11975_ (.A1(_04743_),
    .A2(_04745_),
    .B1(_04747_),
    .C1(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__buf_2 _11976_ (.A(net27),
    .X(_04750_));
 sky130_fd_sc_hd__mux4_1 _11977_ (.A0(_03906_),
    .A1(_04499_),
    .A2(_03909_),
    .A3(_04500_),
    .S0(_04737_),
    .S1(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__nand2_1 _11978_ (.A(net29),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nor2_1 _11979_ (.A(_04503_),
    .B(_04750_),
    .Y(_04753_));
 sky130_fd_sc_hd__a211o_1 _11980_ (.A1(_03852_),
    .A2(_04750_),
    .B1(net29),
    .C1(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__mux4_1 _11981_ (.A0(_04507_),
    .A1(_04508_),
    .A2(_03520_),
    .A3(_03515_),
    .S0(_04750_),
    .S1(net29),
    .X(_04755_));
 sky130_fd_sc_hd__o211ai_1 _11982_ (.A1(net28),
    .A2(_04755_),
    .B1(_04739_),
    .C1(net32),
    .Y(_04756_));
 sky130_fd_sc_hd__a31o_1 _11983_ (.A1(net28),
    .A2(_04752_),
    .A3(_04754_),
    .B1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a21boi_2 _11984_ (.A1(_04723_),
    .A2(_04749_),
    .B1_N(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__a21o_1 _11985_ (.A1(net52),
    .A2(_04723_),
    .B1(net48),
    .X(_04759_));
 sky130_fd_sc_hd__a22o_1 _11986_ (.A1(net47),
    .A2(_04730_),
    .B1(_04732_),
    .B2(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__a221o_1 _11987_ (.A1(net69),
    .A2(_04731_),
    .B1(_04724_),
    .B2(_03910_),
    .C1(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__a22o_1 _11988_ (.A1(net39),
    .A2(_04731_),
    .B1(_04724_),
    .B2(net49),
    .X(_04762_));
 sky130_fd_sc_hd__a221o_1 _11989_ (.A1(net40),
    .A2(_04730_),
    .B1(_04732_),
    .B2(_03537_),
    .C1(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__a32o_1 _11990_ (.A1(net43),
    .A2(_04730_),
    .A3(_04725_),
    .B1(_04726_),
    .B2(net42),
    .X(_04764_));
 sky130_fd_sc_hd__and3_1 _11991_ (.A(net44),
    .B(_04731_),
    .C(_04725_),
    .X(_04765_));
 sky130_fd_sc_hd__a31o_1 _11992_ (.A1(_03911_),
    .A2(_04732_),
    .A3(_04725_),
    .B1(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__a311o_1 _11993_ (.A1(net30),
    .A2(_04742_),
    .A3(_04763_),
    .B1(_04764_),
    .C1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__a21oi_1 _11994_ (.A1(_04743_),
    .A2(_04761_),
    .B1(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__or3b_1 _11995_ (.A(net31),
    .B(_04768_),
    .C_N(net32),
    .X(_04769_));
 sky130_fd_sc_hd__and3_2 _11996_ (.A(_04741_),
    .B(_04758_),
    .C(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__nand2_1 _11997_ (.A(_04750_),
    .B(_04314_),
    .Y(_04771_));
 sky130_fd_sc_hd__o211a_1 _11998_ (.A1(_04750_),
    .A2(net62),
    .B1(_04771_),
    .C1(net31),
    .X(_04772_));
 sky130_fd_sc_hd__nor2_1 _11999_ (.A(_04750_),
    .B(_04393_),
    .Y(_04773_));
 sky130_fd_sc_hd__a211o_1 _12000_ (.A1(_04750_),
    .A2(net65),
    .B1(_04737_),
    .C1(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__and4b_1 _12001_ (.A_N(net32),
    .B(_04774_),
    .C(net28),
    .D(net29),
    .X(_04775_));
 sky130_fd_sc_hd__nor2_1 _12002_ (.A(_04750_),
    .B(_03913_),
    .Y(_04776_));
 sky130_fd_sc_hd__a211o_1 _12003_ (.A1(_04750_),
    .A2(net67),
    .B1(_04776_),
    .C1(net31),
    .X(_04777_));
 sky130_fd_sc_hd__o211ai_1 _12004_ (.A1(net30),
    .A2(_04772_),
    .B1(_04775_),
    .C1(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__a32oi_2 _12005_ (.A1(_04393_),
    .A2(_04723_),
    .A3(_04726_),
    .B1(_04770_),
    .B2(_04778_),
    .Y(net58));
 sky130_fd_sc_hd__buf_2 _12006_ (.A(net33),
    .X(_04779_));
 sky130_fd_sc_hd__or4_1 _12007_ (.A(net36),
    .B(net37),
    .C(net38),
    .D(net65),
    .X(_04780_));
 sky130_fd_sc_hd__nor2_1 _12008_ (.A(_04779_),
    .B(_03913_),
    .Y(_04781_));
 sky130_fd_sc_hd__a211o_1 _12009_ (.A1(_04779_),
    .A2(net67),
    .B1(_04781_),
    .C1(net37),
    .X(_04782_));
 sky130_fd_sc_hd__nand2_1 _12010_ (.A(_04779_),
    .B(_04314_),
    .Y(_04783_));
 sky130_fd_sc_hd__or2_1 _12011_ (.A(_04779_),
    .B(net62),
    .X(_04784_));
 sky130_fd_sc_hd__a31o_1 _12012_ (.A1(net37),
    .A2(_04783_),
    .A3(_04784_),
    .B1(net36),
    .X(_04785_));
 sky130_fd_sc_hd__nor2_1 _12013_ (.A(_04779_),
    .B(_04393_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2_1 _12014_ (.A(net36),
    .B(net37),
    .Y(_04787_));
 sky130_fd_sc_hd__a211o_1 _12015_ (.A1(_04779_),
    .A2(net65),
    .B1(_04786_),
    .C1(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__and4b_1 _12016_ (.A_N(net38),
    .B(_04788_),
    .C(net34),
    .D(net35),
    .X(_04789_));
 sky130_fd_sc_hd__clkbuf_4 _12017_ (.A(net33),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_1 _12018_ (.A(net34),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__inv_2 _12019_ (.A(net34),
    .Y(_04792_));
 sky130_fd_sc_hd__and3_1 _12020_ (.A(net44),
    .B(_04792_),
    .C(_04790_),
    .X(_04793_));
 sky130_fd_sc_hd__nor2_1 _12021_ (.A(_04792_),
    .B(net33),
    .Y(_04794_));
 sky130_fd_sc_hd__a211o_1 _12022_ (.A1(net43),
    .A2(_04794_),
    .B1(net35),
    .C1(net36),
    .X(_04795_));
 sky130_fd_sc_hd__a211o_1 _12023_ (.A1(net42),
    .A2(_04791_),
    .B1(_04793_),
    .C1(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__a31o_1 _12024_ (.A1(net34),
    .A2(_04779_),
    .A3(_03911_),
    .B1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__inv_2 _12025_ (.A(net36),
    .Y(_04798_));
 sky130_fd_sc_hd__mux4_1 _12026_ (.A0(net47),
    .A1(net48),
    .A2(_03910_),
    .A3(net69),
    .S0(_04790_),
    .S1(_04792_),
    .X(_04799_));
 sky130_fd_sc_hd__mux4_1 _12027_ (.A0(net49),
    .A1(net40),
    .A2(net39),
    .A3(_03537_),
    .S0(net34),
    .S1(_04790_),
    .X(_04800_));
 sky130_fd_sc_hd__inv_2 _12028_ (.A(net35),
    .Y(_04801_));
 sky130_fd_sc_hd__o21a_1 _12029_ (.A1(_04798_),
    .A2(_04800_),
    .B1(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__a21o_1 _12030_ (.A1(_04798_),
    .A2(_04799_),
    .B1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__mux4_1 _12031_ (.A0(\gpout0.hpos[0] ),
    .A1(_03527_),
    .A2(_03526_),
    .A3(_04020_),
    .S0(_04790_),
    .S1(net34),
    .X(_04804_));
 sky130_fd_sc_hd__a31o_1 _12032_ (.A1(net36),
    .A2(net35),
    .A3(_04804_),
    .B1(net37),
    .X(_04805_));
 sky130_fd_sc_hd__a21o_1 _12033_ (.A1(_04797_),
    .A2(_04803_),
    .B1(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__mux4_1 _12034_ (.A0(_04507_),
    .A1(_04508_),
    .A2(_03520_),
    .A3(_03515_),
    .S0(_04790_),
    .S1(net35),
    .X(_04807_));
 sky130_fd_sc_hd__nor2_1 _12035_ (.A(_04792_),
    .B(net35),
    .Y(_04808_));
 sky130_fd_sc_hd__mux2_1 _12036_ (.A0(_04503_),
    .A1(_03902_),
    .S(_04790_),
    .X(_04809_));
 sky130_fd_sc_hd__a221o_1 _12037_ (.A1(_04792_),
    .A2(_04807_),
    .B1(_04808_),
    .B2(_04809_),
    .C1(_04798_),
    .X(_04810_));
 sky130_fd_sc_hd__mux4_1 _12038_ (.A0(_03524_),
    .A1(_03461_),
    .A2(_03459_),
    .A3(_03469_),
    .S0(_04790_),
    .S1(net35),
    .X(_04811_));
 sky130_fd_sc_hd__mux2_1 _12039_ (.A0(_03838_),
    .A1(_02901_),
    .S(_04779_),
    .X(_04812_));
 sky130_fd_sc_hd__a221o_1 _12040_ (.A1(_04792_),
    .A2(_04811_),
    .B1(_04812_),
    .B2(_04808_),
    .C1(net36),
    .X(_04813_));
 sky130_fd_sc_hd__mux2_1 _12041_ (.A0(\gpout0.vpos[0] ),
    .A1(\gpout0.vpos[1] ),
    .S(_04790_),
    .X(_04814_));
 sky130_fd_sc_hd__or2b_1 _12042_ (.A(_04814_),
    .B_N(_04787_),
    .X(_04815_));
 sky130_fd_sc_hd__mux2_1 _12043_ (.A0(_03906_),
    .A1(_03909_),
    .S(_04790_),
    .X(_04816_));
 sky130_fd_sc_hd__o211a_1 _12044_ (.A1(_04787_),
    .A2(_04816_),
    .B1(net34),
    .C1(net35),
    .X(_04817_));
 sky130_fd_sc_hd__a21bo_1 _12045_ (.A1(_04815_),
    .A2(_04817_),
    .B1_N(net37),
    .X(_04818_));
 sky130_fd_sc_hd__a21o_1 _12046_ (.A1(_04810_),
    .A2(_04813_),
    .B1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__mux4_1 _12047_ (.A0(net50),
    .A1(net51),
    .A2(net53),
    .A3(_04532_),
    .S0(_04779_),
    .S1(net34),
    .X(_04820_));
 sky130_fd_sc_hd__and3_1 _12048_ (.A(net34),
    .B(net33),
    .C(\gpout5.clk_div[1] ),
    .X(_04821_));
 sky130_fd_sc_hd__a2111oi_2 _12049_ (.A1(clknet_leaf_27_i_clk),
    .A2(_04794_),
    .B1(_04791_),
    .C1(_04821_),
    .D1(net35),
    .Y(_04822_));
 sky130_fd_sc_hd__or4_2 _12050_ (.A(net36),
    .B(net37),
    .C(net38),
    .D(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__o21ba_2 _12051_ (.A1(_04801_),
    .A2(_04820_),
    .B1_N(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__a31o_2 _12052_ (.A1(net38),
    .A2(_04806_),
    .A3(_04819_),
    .B1(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__a31o_2 _12053_ (.A1(_04782_),
    .A2(_04785_),
    .A3(_04789_),
    .B1(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__o41a_2 _12054_ (.A1(net34),
    .A2(_04779_),
    .A3(net35),
    .A4(_04780_),
    .B1(_04826_),
    .X(net59));
 sky130_fd_sc_hd__inv_2 _12055_ (.A(\rbzero.hsync ),
    .Y(net60));
 sky130_fd_sc_hd__buf_4 _12056_ (.A(_02907_),
    .X(_04827_));
 sky130_fd_sc_hd__buf_6 _12057_ (.A(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__and3_1 _12058_ (.A(net72),
    .B(\rbzero.wall_tracer.state[2] ),
    .C(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__clkbuf_1 _12059_ (.A(_04829_),
    .X(_00006_));
 sky130_fd_sc_hd__clkinv_2 _12060_ (.A(\rbzero.wall_tracer.state[3] ),
    .Y(_04830_));
 sky130_fd_sc_hd__clkbuf_4 _12061_ (.A(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__buf_4 _12062_ (.A(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__nor2_1 _12063_ (.A(_04832_),
    .B(_03486_),
    .Y(_00007_));
 sky130_fd_sc_hd__and3_2 _12064_ (.A(net72),
    .B(\rbzero.wall_tracer.state[4] ),
    .C(_02907_),
    .X(_04833_));
 sky130_fd_sc_hd__buf_4 _12065_ (.A(_04833_),
    .X(_00008_));
 sky130_fd_sc_hd__buf_6 _12066_ (.A(_04827_),
    .X(_04834_));
 sky130_fd_sc_hd__and3_1 _12067_ (.A(net72),
    .B(\rbzero.wall_tracer.state[7] ),
    .C(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _12068_ (.A(_04835_),
    .X(_00002_));
 sky130_fd_sc_hd__nor2_1 _12069_ (.A(_03481_),
    .B(_03486_),
    .Y(_00003_));
 sky130_fd_sc_hd__and3_2 _12070_ (.A(net72),
    .B(\rbzero.wall_tracer.state[9] ),
    .C(_02907_),
    .X(_04836_));
 sky130_fd_sc_hd__buf_4 _12071_ (.A(_04836_),
    .X(_00004_));
 sky130_fd_sc_hd__and3_1 _12072_ (.A(net72),
    .B(\rbzero.wall_tracer.state[12] ),
    .C(_04834_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_1 _12073_ (.A(_04837_),
    .X(_00001_));
 sky130_fd_sc_hd__inv_4 _12074_ (.A(\rbzero.wall_tracer.state[6] ),
    .Y(_04838_));
 sky130_fd_sc_hd__clkbuf_4 _12075_ (.A(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__clkbuf_4 _12076_ (.A(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__buf_4 _12077_ (.A(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__nor2_1 _12078_ (.A(_04841_),
    .B(_03486_),
    .Y(_00010_));
 sky130_fd_sc_hd__and3_1 _12079_ (.A(net72),
    .B(\rbzero.wall_tracer.state[5] ),
    .C(_04834_),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_1 _12080_ (.A(_04842_),
    .X(_00009_));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_04843_));
 sky130_fd_sc_hd__or2_1 _12082_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_04844_));
 sky130_fd_sc_hd__nand2_1 _12083_ (.A(_04843_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_04846_));
 sky130_fd_sc_hd__or2_1 _12085_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_04847_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(_04846_),
    .B(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__or2_1 _12087_ (.A(_04845_),
    .B(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__and2_1 _12088_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_04850_));
 sky130_fd_sc_hd__nor2_1 _12089_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_04851_));
 sky130_fd_sc_hd__nor2_1 _12090_ (.A(_04850_),
    .B(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__nor2_1 _12091_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_04853_));
 sky130_fd_sc_hd__nand2_1 _12092_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_04854_));
 sky130_fd_sc_hd__and2b_1 _12093_ (.A_N(_04853_),
    .B(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__nand2_1 _12094_ (.A(_04852_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__or2_1 _12095_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_04857_));
 sky130_fd_sc_hd__or2_1 _12096_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_04858_));
 sky130_fd_sc_hd__nand2_1 _12097_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_04859_));
 sky130_fd_sc_hd__xnor2_1 _12098_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_04860_));
 sky130_fd_sc_hd__nand2_1 _12099_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_04861_));
 sky130_fd_sc_hd__o21ai_1 _12100_ (.A1(_04859_),
    .A2(_04860_),
    .B1(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__and2_1 _12101_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_04863_));
 sky130_fd_sc_hd__a221o_1 _12102_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_04858_),
    .B2(_04862_),
    .C1(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__or4bb_1 _12103_ (.A(_04849_),
    .B(_04856_),
    .C_N(_04857_),
    .D_N(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__and2b_1 _12104_ (.A_N(_04850_),
    .B(_04854_),
    .X(_04866_));
 sky130_fd_sc_hd__or2_1 _12105_ (.A(_04853_),
    .B(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__or2b_1 _12106_ (.A(_04846_),
    .B_N(_04844_),
    .X(_04868_));
 sky130_fd_sc_hd__o211a_1 _12107_ (.A1(_04849_),
    .A2(_04867_),
    .B1(_04868_),
    .C1(_04843_),
    .X(_04869_));
 sky130_fd_sc_hd__and2_1 _12108_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_04870_));
 sky130_fd_sc_hd__nor2_1 _12109_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_04871_));
 sky130_fd_sc_hd__or2_1 _12110_ (.A(_04870_),
    .B(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__a21oi_2 _12111_ (.A1(_04865_),
    .A2(_04869_),
    .B1(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__nand2_1 _12112_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_04874_));
 sky130_fd_sc_hd__or2b_1 _12113_ (.A(_04870_),
    .B_N(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__or2_1 _12114_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_04876_));
 sky130_fd_sc_hd__o221a_1 _12115_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(\rbzero.wall_tracer.rayAddendY[9] ),
    .B1(_04873_),
    .B2(_04875_),
    .C1(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__and2_1 _12116_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_04878_));
 sky130_fd_sc_hd__nor2_1 _12117_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_04879_));
 sky130_fd_sc_hd__nand2_1 _12118_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_04880_));
 sky130_fd_sc_hd__o31a_1 _12119_ (.A1(_04877_),
    .A2(_04878_),
    .A3(_04879_),
    .B1(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__or2_1 _12120_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_04882_));
 sky130_fd_sc_hd__nand2_1 _12121_ (.A(_04880_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__o21bai_1 _12122_ (.A1(_04877_),
    .A2(_04878_),
    .B1_N(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__or3b_1 _12123_ (.A(_04877_),
    .B(_04878_),
    .C_N(_04883_),
    .X(_04885_));
 sky130_fd_sc_hd__and2_1 _12124_ (.A(_04884_),
    .B(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__and3_1 _12125_ (.A(_04865_),
    .B(_04869_),
    .C(_04872_),
    .X(_04887_));
 sky130_fd_sc_hd__nor2_1 _12126_ (.A(_04873_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__and2b_1 _12127_ (.A_N(_04863_),
    .B(_04858_),
    .X(_04889_));
 sky130_fd_sc_hd__xor2_1 _12128_ (.A(_04889_),
    .B(_04862_),
    .X(_04890_));
 sky130_fd_sc_hd__nand2_1 _12129_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_04891_));
 sky130_fd_sc_hd__nand2_1 _12130_ (.A(_04857_),
    .B(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21oi_1 _12131_ (.A1(_04858_),
    .A2(_04862_),
    .B1(_04863_),
    .Y(_04893_));
 sky130_fd_sc_hd__xnor2_1 _12132_ (.A(_04892_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__or2_1 _12133_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_04895_));
 sky130_fd_sc_hd__nand2_1 _12134_ (.A(_04859_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__or4bb_1 _12135_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C_N(_04894_),
    .D_N(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__xnor2_2 _12136_ (.A(_04859_),
    .B(_04860_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand3_1 _12137_ (.A(_04857_),
    .B(_04864_),
    .C(_04852_),
    .Y(_04899_));
 sky130_fd_sc_hd__a21o_1 _12138_ (.A1(_04857_),
    .A2(_04864_),
    .B1(_04852_),
    .X(_04900_));
 sky130_fd_sc_hd__nand2_1 _12139_ (.A(_04899_),
    .B(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__or4bb_1 _12140_ (.A(_04890_),
    .B(_04897_),
    .C_N(_04898_),
    .D_N(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__a31o_1 _12141_ (.A1(_04857_),
    .A2(_04864_),
    .A3(_04852_),
    .B1(_04850_),
    .X(_04903_));
 sky130_fd_sc_hd__xor2_2 _12142_ (.A(_04855_),
    .B(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__a211o_1 _12143_ (.A1(_04899_),
    .A2(_04866_),
    .B1(_04853_),
    .C1(_04848_),
    .X(_04905_));
 sky130_fd_sc_hd__o211ai_1 _12144_ (.A1(_04899_),
    .A2(_04853_),
    .B1(_04867_),
    .C1(_04848_),
    .Y(_04906_));
 sky130_fd_sc_hd__nand2_1 _12145_ (.A(_04905_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__or4b_1 _12146_ (.A(_04888_),
    .B(_04902_),
    .C(_04904_),
    .D_N(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__a21o_1 _12147_ (.A1(_04846_),
    .A2(_04905_),
    .B1(_04845_),
    .X(_04909_));
 sky130_fd_sc_hd__nand3_1 _12148_ (.A(_04845_),
    .B(_04846_),
    .C(_04905_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand2_1 _12149_ (.A(_04909_),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__nand2_1 _12150_ (.A(_04876_),
    .B(_04874_),
    .Y(_04912_));
 sky130_fd_sc_hd__o21bai_1 _12151_ (.A1(_04870_),
    .A2(_04873_),
    .B1_N(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__or3b_1 _12152_ (.A(_04870_),
    .B(_04873_),
    .C_N(_04912_),
    .X(_04914_));
 sky130_fd_sc_hd__nand2_1 _12153_ (.A(_04913_),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__nand2_1 _12154_ (.A(_04911_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__o21a_1 _12155_ (.A1(_04873_),
    .A2(_04875_),
    .B1(_04876_),
    .X(_04917_));
 sky130_fd_sc_hd__nor2_1 _12156_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_04918_));
 sky130_fd_sc_hd__nor2_1 _12157_ (.A(_04918_),
    .B(_04878_),
    .Y(_04919_));
 sky130_fd_sc_hd__xnor2_1 _12158_ (.A(_04917_),
    .B(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__or4b_1 _12159_ (.A(_04886_),
    .B(_04908_),
    .C(_04916_),
    .D_N(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__nand2_1 _12160_ (.A(_04881_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__clkbuf_4 _12161_ (.A(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__nand2_1 _12162_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__or2_1 _12163_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_04923_),
    .X(_04925_));
 sky130_fd_sc_hd__and2_1 _12164_ (.A(_04924_),
    .B(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__and2_2 _12165_ (.A(_04881_),
    .B(_04921_),
    .X(_04927_));
 sky130_fd_sc_hd__clkbuf_4 _12166_ (.A(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__clkbuf_4 _12167_ (.A(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__a21oi_1 _12168_ (.A1(_03359_),
    .A2(_03351_),
    .B1(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__xnor2_1 _12169_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .B(_04929_),
    .Y(_04931_));
 sky130_fd_sc_hd__xnor2_1 _12170_ (.A(\rbzero.map_rom.i_row[4] ),
    .B(_04929_),
    .Y(_04932_));
 sky130_fd_sc_hd__nor2_1 _12171_ (.A(_03375_),
    .B(_04929_),
    .Y(_04933_));
 sky130_fd_sc_hd__xnor2_1 _12172_ (.A(_03358_),
    .B(_04928_),
    .Y(_04934_));
 sky130_fd_sc_hd__nand2_1 _12173_ (.A(_03390_),
    .B(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__o21ai_1 _12174_ (.A1(_03374_),
    .A2(_04928_),
    .B1(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__nor2_1 _12175_ (.A(_03346_),
    .B(_04928_),
    .Y(_04937_));
 sky130_fd_sc_hd__nor2_1 _12176_ (.A(_03345_),
    .B(_04923_),
    .Y(_04938_));
 sky130_fd_sc_hd__nor2_1 _12177_ (.A(_04937_),
    .B(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__a21o_1 _12178_ (.A1(_04936_),
    .A2(_04939_),
    .B1(_04937_),
    .X(_04940_));
 sky130_fd_sc_hd__nand2_1 _12179_ (.A(_03375_),
    .B(_04929_),
    .Y(_04941_));
 sky130_fd_sc_hd__o21a_1 _12180_ (.A1(_04933_),
    .A2(_04940_),
    .B1(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__and2_1 _12181_ (.A(_04932_),
    .B(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__and2_1 _12182_ (.A(_04931_),
    .B(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__or3_1 _12183_ (.A(_04926_),
    .B(_04930_),
    .C(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__buf_4 _12184_ (.A(_03341_),
    .X(_04946_));
 sky130_fd_sc_hd__buf_4 _12185_ (.A(\rbzero.wall_tracer.state[6] ),
    .X(_04947_));
 sky130_fd_sc_hd__buf_4 _12186_ (.A(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__buf_4 _12187_ (.A(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__clkbuf_4 _12188_ (.A(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__nor2_1 _12189_ (.A(\rbzero.wall_tracer.state[1] ),
    .B(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__nand2_1 _12190_ (.A(_03483_),
    .B(_03458_),
    .Y(_04952_));
 sky130_fd_sc_hd__inv_2 _12191_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .Y(_04953_));
 sky130_fd_sc_hd__inv_2 _12192_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(_04954_),
    .B(\rbzero.wall_tracer.trackDistX[9] ),
    .Y(_04955_));
 sky130_fd_sc_hd__inv_2 _12194_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .Y(_04956_));
 sky130_fd_sc_hd__inv_2 _12195_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .Y(_04957_));
 sky130_fd_sc_hd__inv_2 _12196_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .Y(_04958_));
 sky130_fd_sc_hd__inv_2 _12197_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .Y(_04959_));
 sky130_fd_sc_hd__inv_2 _12198_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .Y(_04960_));
 sky130_fd_sc_hd__inv_2 _12199_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .Y(_04961_));
 sky130_fd_sc_hd__inv_2 _12200_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .Y(_04962_));
 sky130_fd_sc_hd__inv_2 _12201_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .Y(_04963_));
 sky130_fd_sc_hd__inv_2 _12202_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .Y(_04964_));
 sky130_fd_sc_hd__a22o_1 _12203_ (.A1(_04963_),
    .A2(\rbzero.wall_tracer.trackDistX[0] ),
    .B1(_04964_),
    .B2(\rbzero.wall_tracer.trackDistX[-1] ),
    .X(_04965_));
 sky130_fd_sc_hd__inv_2 _12204_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .Y(_04966_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__o21ai_1 _12206_ (.A1(_04964_),
    .A2(\rbzero.wall_tracer.trackDistX[-1] ),
    .B1(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__nor2_1 _12207_ (.A(_04965_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__inv_2 _12208_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .Y(_04970_));
 sky130_fd_sc_hd__inv_2 _12209_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .Y(_04971_));
 sky130_fd_sc_hd__inv_2 _12210_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .Y(_04972_));
 sky130_fd_sc_hd__inv_2 _12211_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .Y(_04973_));
 sky130_fd_sc_hd__inv_2 _12212_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .Y(_04974_));
 sky130_fd_sc_hd__inv_2 _12213_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .Y(_04975_));
 sky130_fd_sc_hd__inv_2 _12214_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .Y(_04976_));
 sky130_fd_sc_hd__inv_2 _12215_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .Y(_04977_));
 sky130_fd_sc_hd__a211o_1 _12216_ (.A1(_04976_),
    .A2(\rbzero.wall_tracer.trackDistX[-10] ),
    .B1(_04977_),
    .C1(\rbzero.wall_tracer.trackDistX[-11] ),
    .X(_04978_));
 sky130_fd_sc_hd__o221a_1 _12217_ (.A1(_04975_),
    .A2(\rbzero.wall_tracer.trackDistX[-9] ),
    .B1(_04976_),
    .B2(\rbzero.wall_tracer.trackDistX[-10] ),
    .C1(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__a221o_1 _12218_ (.A1(_04974_),
    .A2(\rbzero.wall_tracer.trackDistX[-8] ),
    .B1(_04975_),
    .B2(\rbzero.wall_tracer.trackDistX[-9] ),
    .C1(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__o221a_1 _12219_ (.A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .A2(_04973_),
    .B1(_04974_),
    .B2(\rbzero.wall_tracer.trackDistX[-8] ),
    .C1(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__a221o_1 _12220_ (.A1(_04972_),
    .A2(\rbzero.wall_tracer.trackDistX[-6] ),
    .B1(\rbzero.wall_tracer.trackDistX[-7] ),
    .B2(_04973_),
    .C1(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__o221a_1 _12221_ (.A1(_04971_),
    .A2(\rbzero.wall_tracer.trackDistX[-5] ),
    .B1(_04972_),
    .B2(\rbzero.wall_tracer.trackDistX[-6] ),
    .C1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__a221o_1 _12222_ (.A1(_04970_),
    .A2(\rbzero.wall_tracer.trackDistX[-4] ),
    .B1(_04971_),
    .B2(\rbzero.wall_tracer.trackDistX[-5] ),
    .C1(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__inv_2 _12223_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .Y(_04985_));
 sky130_fd_sc_hd__inv_2 _12224_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .Y(_04986_));
 sky130_fd_sc_hd__a22o_1 _12225_ (.A1(_04985_),
    .A2(\rbzero.wall_tracer.trackDistX[-2] ),
    .B1(\rbzero.wall_tracer.trackDistX[-3] ),
    .B2(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__or2_1 _12226_ (.A(_04985_),
    .B(\rbzero.wall_tracer.trackDistX[-2] ),
    .X(_04988_));
 sky130_fd_sc_hd__o22a_1 _12227_ (.A1(\rbzero.wall_tracer.trackDistX[-3] ),
    .A2(_04986_),
    .B1(_04970_),
    .B2(\rbzero.wall_tracer.trackDistX[-4] ),
    .X(_04989_));
 sky130_fd_sc_hd__or2b_1 _12228_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B_N(\rbzero.wall_tracer.trackDistY[1] ),
    .X(_04990_));
 sky130_fd_sc_hd__and4b_1 _12229_ (.A_N(_04987_),
    .B(_04988_),
    .C(_04989_),
    .D(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__a32o_1 _12230_ (.A1(_04969_),
    .A2(_04987_),
    .A3(_04988_),
    .B1(_04967_),
    .B2(_04965_),
    .X(_04992_));
 sky130_fd_sc_hd__and2b_1 _12231_ (.A_N(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.trackDistX[1] ),
    .X(_04993_));
 sky130_fd_sc_hd__a221o_1 _12232_ (.A1(_04962_),
    .A2(\rbzero.wall_tracer.trackDistX[2] ),
    .B1(_04990_),
    .B2(_04992_),
    .C1(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__a31o_1 _12233_ (.A1(_04969_),
    .A2(_04984_),
    .A3(_04991_),
    .B1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__o221a_1 _12234_ (.A1(_04961_),
    .A2(\rbzero.wall_tracer.trackDistX[3] ),
    .B1(_04962_),
    .B2(\rbzero.wall_tracer.trackDistX[2] ),
    .C1(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__a221o_1 _12235_ (.A1(_04960_),
    .A2(\rbzero.wall_tracer.trackDistX[4] ),
    .B1(_04961_),
    .B2(\rbzero.wall_tracer.trackDistX[3] ),
    .C1(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__o221a_1 _12236_ (.A1(\rbzero.wall_tracer.trackDistX[5] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\rbzero.wall_tracer.trackDistX[4] ),
    .C1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__a221o_1 _12237_ (.A1(_04958_),
    .A2(\rbzero.wall_tracer.trackDistX[6] ),
    .B1(\rbzero.wall_tracer.trackDistX[5] ),
    .B2(_04959_),
    .C1(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__o221a_1 _12238_ (.A1(_04957_),
    .A2(\rbzero.wall_tracer.trackDistX[7] ),
    .B1(_04958_),
    .B2(\rbzero.wall_tracer.trackDistX[6] ),
    .C1(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__a221o_1 _12239_ (.A1(_04956_),
    .A2(\rbzero.wall_tracer.trackDistX[8] ),
    .B1(_04957_),
    .B2(\rbzero.wall_tracer.trackDistX[7] ),
    .C1(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__o22a_1 _12240_ (.A1(_04954_),
    .A2(\rbzero.wall_tracer.trackDistX[9] ),
    .B1(_04956_),
    .B2(\rbzero.wall_tracer.trackDistX[8] ),
    .X(_05002_));
 sky130_fd_sc_hd__a32oi_2 _12241_ (.A1(_04955_),
    .A2(_05001_),
    .A3(_05002_),
    .B1(_04953_),
    .B2(\rbzero.wall_tracer.trackDistX[10] ),
    .Y(_05003_));
 sky130_fd_sc_hd__a2bb2o_1 _12242_ (.A1_N(\rbzero.wall_tracer.trackDistX[10] ),
    .A2_N(_04953_),
    .B1(_04955_),
    .B2(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__nand2_1 _12243_ (.A(_03495_),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__or3b_4 _12244_ (.A(_04951_),
    .B(_04952_),
    .C_N(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__nor2_2 _12245_ (.A(_04946_),
    .B(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__o21ai_1 _12246_ (.A1(_04930_),
    .A2(_04944_),
    .B1(_04926_),
    .Y(_05008_));
 sky130_fd_sc_hd__clkbuf_4 _12247_ (.A(_05006_),
    .X(_05009_));
 sky130_fd_sc_hd__a32o_1 _12248_ (.A1(_04945_),
    .A2(_05007_),
    .A3(_05008_),
    .B1(_05009_),
    .B2(\rbzero.wall_tracer.mapY[6] ),
    .X(_00401_));
 sky130_fd_sc_hd__xnor2_1 _12249_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .B(_04923_),
    .Y(_05010_));
 sky130_fd_sc_hd__nand3_1 _12250_ (.A(_04924_),
    .B(_05008_),
    .C(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__a21o_1 _12251_ (.A1(_04924_),
    .A2(_05008_),
    .B1(_05010_),
    .X(_05012_));
 sky130_fd_sc_hd__a32o_1 _12252_ (.A1(_05007_),
    .A2(_05011_),
    .A3(_05012_),
    .B1(_05009_),
    .B2(\rbzero.wall_tracer.mapY[7] ),
    .X(_00402_));
 sky130_fd_sc_hd__clkinv_2 _12253_ (.A(_05010_),
    .Y(_05013_));
 sky130_fd_sc_hd__and3_1 _12254_ (.A(_04926_),
    .B(_04944_),
    .C(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__o41a_1 _12255_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(\rbzero.wall_tracer.mapY[5] ),
    .A3(\rbzero.wall_tracer.mapY[7] ),
    .A4(\rbzero.wall_tracer.mapY[6] ),
    .B1(_04923_),
    .X(_05015_));
 sky130_fd_sc_hd__xnor2_1 _12256_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_04929_),
    .Y(_05016_));
 sky130_fd_sc_hd__o21a_1 _12257_ (.A1(_05014_),
    .A2(_05015_),
    .B1(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__o31ai_1 _12258_ (.A1(_05016_),
    .A2(_05014_),
    .A3(_05015_),
    .B1(_05007_),
    .Y(_05018_));
 sky130_fd_sc_hd__a2bb2o_1 _12259_ (.A1_N(_05017_),
    .A2_N(_05018_),
    .B1(\rbzero.wall_tracer.mapY[8] ),
    .B2(_05009_),
    .X(_00403_));
 sky130_fd_sc_hd__a21o_1 _12260_ (.A1(\rbzero.wall_tracer.mapY[8] ),
    .A2(_04923_),
    .B1(_05017_),
    .X(_05019_));
 sky130_fd_sc_hd__xnor2_1 _12261_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(_04929_),
    .Y(_05020_));
 sky130_fd_sc_hd__or2_1 _12262_ (.A(_05019_),
    .B(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__nand2_1 _12263_ (.A(_05019_),
    .B(_05020_),
    .Y(_05022_));
 sky130_fd_sc_hd__a32o_1 _12264_ (.A1(_05007_),
    .A2(_05021_),
    .A3(_05022_),
    .B1(_05009_),
    .B2(\rbzero.wall_tracer.mapY[9] ),
    .X(_00404_));
 sky130_fd_sc_hd__o21a_1 _12265_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_04923_),
    .B1(_05019_),
    .X(_05023_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_04923_),
    .B1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__xnor2_1 _12267_ (.A(\rbzero.wall_tracer.mapY[10] ),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__or2_1 _12268_ (.A(_04929_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__nand2_1 _12269_ (.A(_04929_),
    .B(_05025_),
    .Y(_05027_));
 sky130_fd_sc_hd__a32o_1 _12270_ (.A1(_05007_),
    .A2(_05026_),
    .A3(_05027_),
    .B1(_05009_),
    .B2(\rbzero.wall_tracer.mapY[10] ),
    .X(_00405_));
 sky130_fd_sc_hd__or2_1 _12271_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_05028_));
 sky130_fd_sc_hd__or2_1 _12272_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_05029_));
 sky130_fd_sc_hd__or2_1 _12273_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_05030_));
 sky130_fd_sc_hd__nand2_1 _12274_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_05031_));
 sky130_fd_sc_hd__inv_2 _12275_ (.A(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__nor2_1 _12276_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_05033_));
 sky130_fd_sc_hd__nor2_1 _12277_ (.A(_05032_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_1 _12278_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_05035_));
 sky130_fd_sc_hd__or2_1 _12279_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_05036_));
 sky130_fd_sc_hd__and2_1 _12280_ (.A(_05035_),
    .B(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__nor2_1 _12281_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_05038_));
 sky130_fd_sc_hd__nor2_1 _12282_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_2 _12283_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_05040_));
 sky130_fd_sc_hd__nor2_1 _12284_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_05041_));
 sky130_fd_sc_hd__nand2_1 _12285_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_05042_));
 sky130_fd_sc_hd__nand2_1 _12286_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_05043_));
 sky130_fd_sc_hd__o211a_1 _12287_ (.A1(_05040_),
    .A2(_05041_),
    .B1(_05042_),
    .C1(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__nand2_1 _12288_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_05045_));
 sky130_fd_sc_hd__o31ai_4 _12289_ (.A1(_05038_),
    .A2(_05039_),
    .A3(_05044_),
    .B1(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__o211a_1 _12290_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(\rbzero.wall_tracer.rayAddendX[5] ),
    .C1(\rbzero.debug_overlay.facingX[-3] ),
    .X(_05047_));
 sky130_fd_sc_hd__a21o_1 _12291_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__a21o_1 _12292_ (.A1(_05031_),
    .A2(_05035_),
    .B1(_05033_),
    .X(_05049_));
 sky130_fd_sc_hd__inv_2 _12293_ (.A(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__a311o_1 _12294_ (.A1(_05034_),
    .A2(_05037_),
    .A3(_05046_),
    .B1(_05048_),
    .C1(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__or2_1 _12295_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_05052_));
 sky130_fd_sc_hd__a21o_1 _12296_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__o21a_1 _12297_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__and2_1 _12298_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_05055_));
 sky130_fd_sc_hd__and2_1 _12299_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_05056_));
 sky130_fd_sc_hd__a311o_1 _12300_ (.A1(_05030_),
    .A2(_05051_),
    .A3(_05054_),
    .B1(_05055_),
    .C1(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__nand2_1 _12301_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_05058_));
 sky130_fd_sc_hd__inv_2 _12302_ (.A(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__a31o_2 _12303_ (.A1(_05028_),
    .A2(_05029_),
    .A3(_05057_),
    .B1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__nor2_1 _12304_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_05061_));
 sky130_fd_sc_hd__nand2_1 _12305_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_05062_));
 sky130_fd_sc_hd__or2b_1 _12306_ (.A(_05061_),
    .B_N(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__xor2_2 _12307_ (.A(_05060_),
    .B(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__nand2_1 _12308_ (.A(_03489_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__inv_2 _12309_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .Y(_05066_));
 sky130_fd_sc_hd__buf_2 _12310_ (.A(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__a21o_1 _12311_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_05067_),
    .B1(_03488_),
    .X(_05068_));
 sky130_fd_sc_hd__a31o_1 _12312_ (.A1(_03480_),
    .A2(_04884_),
    .A3(_04885_),
    .B1(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__nor2_1 _12313_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_03480_),
    .Y(_05070_));
 sky130_fd_sc_hd__a211oi_2 _12314_ (.A1(_03480_),
    .A2(_04920_),
    .B1(_05070_),
    .C1(_03489_),
    .Y(_05071_));
 sky130_fd_sc_hd__inv_2 _12315_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_1 _12316_ (.A(_05029_),
    .B(_05057_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_1 _12317_ (.A(_05028_),
    .B(_05058_),
    .Y(_05074_));
 sky130_fd_sc_hd__xnor2_2 _12318_ (.A(_05073_),
    .B(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__nor2_1 _12319_ (.A(_05072_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__a211oi_4 _12320_ (.A1(_05065_),
    .A2(_05069_),
    .B1(_05071_),
    .C1(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__o311a_4 _12321_ (.A1(_04877_),
    .A2(_04878_),
    .A3(_04879_),
    .B1(_04880_),
    .C1(_03479_),
    .X(_05078_));
 sky130_fd_sc_hd__nor2_1 _12322_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_03480_),
    .Y(_05079_));
 sky130_fd_sc_hd__a211o_4 _12323_ (.A1(_05062_),
    .A2(_05060_),
    .B1(_05072_),
    .C1(_05061_),
    .X(_05080_));
 sky130_fd_sc_hd__o31ai_4 _12324_ (.A1(_03489_),
    .A2(_05078_),
    .A3(_05079_),
    .B1(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__xor2_1 _12325_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_05082_));
 sky130_fd_sc_hd__a31o_1 _12326_ (.A1(_05034_),
    .A2(_05037_),
    .A3(_05046_),
    .B1(_05050_),
    .X(_05083_));
 sky130_fd_sc_hd__nand2_1 _12327_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_05084_));
 sky130_fd_sc_hd__a21bo_1 _12328_ (.A1(_05052_),
    .A2(_05083_),
    .B1_N(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__xnor2_2 _12329_ (.A(_05082_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__nand2_1 _12330_ (.A(_03488_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__a21o_1 _12331_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_05067_),
    .B1(_03487_),
    .X(_05088_));
 sky130_fd_sc_hd__a31o_1 _12332_ (.A1(_03479_),
    .A2(_04909_),
    .A3(_04910_),
    .B1(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__nand2_1 _12333_ (.A(_05084_),
    .B(_05052_),
    .Y(_05090_));
 sky130_fd_sc_hd__xor2_2 _12334_ (.A(_05090_),
    .B(_05083_),
    .X(_05091_));
 sky130_fd_sc_hd__and3_1 _12335_ (.A(_03479_),
    .B(_04905_),
    .C(_04906_),
    .X(_05092_));
 sky130_fd_sc_hd__a21o_1 _12336_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_05067_),
    .B1(_03487_),
    .X(_05093_));
 sky130_fd_sc_hd__o2bb2a_2 _12337_ (.A1_N(_03488_),
    .A2_N(_05091_),
    .B1(_05092_),
    .B2(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__a21bo_1 _12338_ (.A1(_05037_),
    .A2(_05046_),
    .B1_N(_05035_),
    .X(_05095_));
 sky130_fd_sc_hd__xnor2_2 _12339_ (.A(_05034_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__nand2_1 _12340_ (.A(_03487_),
    .B(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__a21o_1 _12341_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_05067_),
    .B1(_03487_),
    .X(_05098_));
 sky130_fd_sc_hd__a21o_1 _12342_ (.A1(_03479_),
    .A2(_04904_),
    .B1(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__nor2_1 _12343_ (.A(_05038_),
    .B(_05044_),
    .Y(_05100_));
 sky130_fd_sc_hd__or2b_1 _12344_ (.A(_05039_),
    .B_N(_05045_),
    .X(_05101_));
 sky130_fd_sc_hd__xnor2_2 _12345_ (.A(_05100_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__nand2_1 _12346_ (.A(_03479_),
    .B(_04894_),
    .Y(_05103_));
 sky130_fd_sc_hd__o21a_1 _12347_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_03479_),
    .B1(_05072_),
    .X(_05104_));
 sky130_fd_sc_hd__a22o_2 _12348_ (.A1(_03487_),
    .A2(_05102_),
    .B1(_05103_),
    .B2(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__and2b_1 _12349_ (.A_N(_05041_),
    .B(_05042_),
    .X(_05106_));
 sky130_fd_sc_hd__xnor2_4 _12350_ (.A(_05040_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__nand2_1 _12351_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .B(_04898_),
    .Y(_05108_));
 sky130_fd_sc_hd__o211a_1 _12352_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(\rbzero.wall_tracer.rcp_sel[2] ),
    .B1(_05072_),
    .C1(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__nor2_1 _12353_ (.A(_05067_),
    .B(_04896_),
    .Y(_05110_));
 sky130_fd_sc_hd__a21o_1 _12354_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_05066_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_05111_));
 sky130_fd_sc_hd__or2_1 _12355_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_05112_));
 sky130_fd_sc_hd__and2_1 _12356_ (.A(_05040_),
    .B(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__o22a_2 _12357_ (.A1(_05110_),
    .A2(_05111_),
    .B1(_05113_),
    .B2(_05072_),
    .X(_05114_));
 sky130_fd_sc_hd__mux2_1 _12358_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05115_));
 sky130_fd_sc_hd__mux2_2 _12359_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_05115_),
    .S(_05072_),
    .X(_05116_));
 sky130_fd_sc_hd__mux2_1 _12360_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05117_));
 sky130_fd_sc_hd__mux2_2 _12361_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_05117_),
    .S(_05072_),
    .X(_05118_));
 sky130_fd_sc_hd__or2_1 _12362_ (.A(_05116_),
    .B(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a2111o_4 _12363_ (.A1(_03487_),
    .A2(_05107_),
    .B1(_05109_),
    .C1(_05114_),
    .D1(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__o21a_1 _12364_ (.A1(_05040_),
    .A2(_05041_),
    .B1(_05042_),
    .X(_05121_));
 sky130_fd_sc_hd__and2_1 _12365_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_05122_));
 sky130_fd_sc_hd__nor2_1 _12366_ (.A(_05122_),
    .B(_05038_),
    .Y(_05123_));
 sky130_fd_sc_hd__xnor2_2 _12367_ (.A(_05121_),
    .B(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A1(_04890_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05125_));
 sky130_fd_sc_hd__mux2_2 _12369_ (.A0(_05124_),
    .A1(_05125_),
    .S(_05072_),
    .X(_05126_));
 sky130_fd_sc_hd__or2_1 _12370_ (.A(_05120_),
    .B(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__xnor2_2 _12371_ (.A(_05037_),
    .B(_05046_),
    .Y(_05128_));
 sky130_fd_sc_hd__a21o_1 _12372_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_05067_),
    .B1(_03487_),
    .X(_05129_));
 sky130_fd_sc_hd__and3_1 _12373_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .B(_04899_),
    .C(_04900_),
    .X(_05130_));
 sky130_fd_sc_hd__o2bb2a_2 _12374_ (.A1_N(_03487_),
    .A2_N(_05128_),
    .B1(_05129_),
    .B2(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__a2111o_1 _12375_ (.A1(_05097_),
    .A2(_05099_),
    .B1(_05105_),
    .C1(_05127_),
    .D1(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__a211o_2 _12376_ (.A1(_05087_),
    .A2(_05089_),
    .B1(_05094_),
    .C1(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__nand2_1 _12377_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_1 _12378_ (.A(_05029_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__a31o_1 _12379_ (.A1(_05030_),
    .A2(_05051_),
    .A3(_05054_),
    .B1(_05056_),
    .X(_05136_));
 sky130_fd_sc_hd__xnor2_2 _12380_ (.A(_05135_),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__or2_1 _12381_ (.A(_05072_),
    .B(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__a21o_1 _12382_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_05067_),
    .B1(_03488_),
    .X(_05139_));
 sky130_fd_sc_hd__a31o_1 _12383_ (.A1(_03479_),
    .A2(_04913_),
    .A3(_04914_),
    .B1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__or2b_2 _12384_ (.A(_05056_),
    .B_N(_05030_),
    .X(_05141_));
 sky130_fd_sc_hd__nand2_2 _12385_ (.A(_05051_),
    .B(_05054_),
    .Y(_05142_));
 sky130_fd_sc_hd__xnor2_4 _12386_ (.A(_05141_),
    .B(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__a21oi_1 _12387_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_05067_),
    .B1(_03487_),
    .Y(_05144_));
 sky130_fd_sc_hd__o31a_1 _12388_ (.A1(_05067_),
    .A2(_04873_),
    .A3(_04887_),
    .B1(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__a21oi_4 _12389_ (.A1(_03488_),
    .A2(_05143_),
    .B1(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__a21o_1 _12390_ (.A1(_05138_),
    .A2(_05140_),
    .B1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__nor2_1 _12391_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_03479_),
    .Y(_05148_));
 sky130_fd_sc_hd__o31a_1 _12392_ (.A1(_03488_),
    .A2(_05078_),
    .A3(_05148_),
    .B1(_05080_),
    .X(_05149_));
 sky130_fd_sc_hd__nor4b_2 _12393_ (.A(_05081_),
    .B(_05133_),
    .C(_05147_),
    .D_N(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__nor2_1 _12394_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_03480_),
    .Y(_05151_));
 sky130_fd_sc_hd__o31a_1 _12395_ (.A1(_03489_),
    .A2(_05078_),
    .A3(_05151_),
    .B1(_05080_),
    .X(_05152_));
 sky130_fd_sc_hd__clkbuf_4 _12396_ (.A(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__a21oi_1 _12397_ (.A1(_05077_),
    .A2(_05150_),
    .B1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__or2_1 _12398_ (.A(_03488_),
    .B(_05078_),
    .X(_05155_));
 sky130_fd_sc_hd__nor2_1 _12399_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_03480_),
    .Y(_05156_));
 sky130_fd_sc_hd__o21a_1 _12400_ (.A1(_05155_),
    .A2(_05156_),
    .B1(_05080_),
    .X(_05157_));
 sky130_fd_sc_hd__xnor2_2 _12401_ (.A(_05154_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__and2_1 _12402_ (.A(_05077_),
    .B(_05150_),
    .X(_05159_));
 sky130_fd_sc_hd__nor2_1 _12403_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_03479_),
    .Y(_05160_));
 sky130_fd_sc_hd__o31a_2 _12404_ (.A1(_03488_),
    .A2(_05078_),
    .A3(_05160_),
    .B1(_05080_),
    .X(_05161_));
 sky130_fd_sc_hd__nor2_1 _12405_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_03480_),
    .Y(_05162_));
 sky130_fd_sc_hd__o31a_2 _12406_ (.A1(_03488_),
    .A2(_05078_),
    .A3(_05162_),
    .B1(_05080_),
    .X(_05163_));
 sky130_fd_sc_hd__inv_2 _12407_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .Y(_05164_));
 sky130_fd_sc_hd__a211o_1 _12408_ (.A1(_05164_),
    .A2(_05067_),
    .B1(_03489_),
    .C1(_05078_),
    .X(_05165_));
 sky130_fd_sc_hd__o2111a_1 _12409_ (.A1(_05155_),
    .A2(_05156_),
    .B1(_05161_),
    .C1(_05163_),
    .D1(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__nand2_1 _12410_ (.A(_05159_),
    .B(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__or4_1 _12411_ (.A(_03388_),
    .B(\rbzero.wall_tracer.visualWallDist[9] ),
    .C(_03480_),
    .D(_03489_),
    .X(_05168_));
 sky130_fd_sc_hd__nor2_1 _12412_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_03480_),
    .Y(_05169_));
 sky130_fd_sc_hd__o21a_1 _12413_ (.A1(_05078_),
    .A2(_05169_),
    .B1(_05072_),
    .X(_05170_));
 sky130_fd_sc_hd__a21o_1 _12414_ (.A1(_05062_),
    .A2(_05060_),
    .B1(_05061_),
    .X(_05171_));
 sky130_fd_sc_hd__a21oi_1 _12415_ (.A1(_03489_),
    .A2(_05171_),
    .B1(_05170_),
    .Y(_05172_));
 sky130_fd_sc_hd__a31o_1 _12416_ (.A1(_05077_),
    .A2(_05150_),
    .A3(_05166_),
    .B1(_05152_),
    .X(_05173_));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(_05170_),
    .A1(_05172_),
    .S(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__o21ba_1 _12418_ (.A1(_05167_),
    .A2(_05168_),
    .B1_N(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__o21a_1 _12419_ (.A1(_05155_),
    .A2(_05156_),
    .B1(_05161_),
    .X(_05176_));
 sky130_fd_sc_hd__a31o_1 _12420_ (.A1(_05077_),
    .A2(_05150_),
    .A3(_05176_),
    .B1(_05152_),
    .X(_05177_));
 sky130_fd_sc_hd__xor2_2 _12421_ (.A(_05163_),
    .B(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__nand2_1 _12422_ (.A(_05080_),
    .B(_05165_),
    .Y(_05179_));
 sky130_fd_sc_hd__a311o_1 _12423_ (.A1(_05159_),
    .A2(_05176_),
    .A3(_05163_),
    .B1(_05179_),
    .C1(_05153_),
    .X(_05180_));
 sky130_fd_sc_hd__o211ai_2 _12424_ (.A1(_05153_),
    .A2(_05163_),
    .B1(_05177_),
    .C1(_05179_),
    .Y(_05181_));
 sky130_fd_sc_hd__and3b_1 _12425_ (.A_N(_05178_),
    .B(_05180_),
    .C(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__a21oi_2 _12426_ (.A1(_05159_),
    .A2(_05157_),
    .B1(_05153_),
    .Y(_05183_));
 sky130_fd_sc_hd__xor2_1 _12427_ (.A(_05161_),
    .B(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__and4b_1 _12428_ (.A_N(_05158_),
    .B(_05175_),
    .C(_05182_),
    .D(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__nor2_1 _12429_ (.A(_05071_),
    .B(_05076_),
    .Y(_05186_));
 sky130_fd_sc_hd__o31ai_2 _12430_ (.A1(_03489_),
    .A2(_05078_),
    .A3(_05151_),
    .B1(_05080_),
    .Y(_05187_));
 sky130_fd_sc_hd__o21ai_2 _12431_ (.A1(_05133_),
    .A2(_05147_),
    .B1(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__xor2_2 _12432_ (.A(_05186_),
    .B(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__nand2_1 _12433_ (.A(_05138_),
    .B(_05140_),
    .Y(_05190_));
 sky130_fd_sc_hd__o21ai_1 _12434_ (.A1(_05133_),
    .A2(_05146_),
    .B1(_05187_),
    .Y(_05191_));
 sky130_fd_sc_hd__xnor2_2 _12435_ (.A(_05190_),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__or2b_1 _12436_ (.A(_05189_),
    .B_N(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__nand2_1 _12437_ (.A(_05065_),
    .B(_05069_),
    .Y(_05194_));
 sky130_fd_sc_hd__nor2_1 _12438_ (.A(_05133_),
    .B(_05147_),
    .Y(_05195_));
 sky130_fd_sc_hd__a21oi_1 _12439_ (.A1(_05186_),
    .A2(_05195_),
    .B1(_05153_),
    .Y(_05196_));
 sky130_fd_sc_hd__xnor2_2 _12440_ (.A(_05194_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__or2_1 _12441_ (.A(_05193_),
    .B(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__buf_2 _12442_ (.A(_05187_),
    .X(_05199_));
 sky130_fd_sc_hd__nand2_2 _12443_ (.A(_05199_),
    .B(_05133_),
    .Y(_05200_));
 sky130_fd_sc_hd__xor2_2 _12444_ (.A(_05146_),
    .B(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__a211o_1 _12445_ (.A1(_05077_),
    .A2(_05195_),
    .B1(_05149_),
    .C1(_05153_),
    .X(_05202_));
 sky130_fd_sc_hd__o211ai_2 _12446_ (.A1(_05153_),
    .A2(_05077_),
    .B1(_05149_),
    .C1(_05188_),
    .Y(_05203_));
 sky130_fd_sc_hd__a311oi_2 _12447_ (.A1(_05077_),
    .A2(_05195_),
    .A3(_05149_),
    .B1(_05081_),
    .C1(_05153_),
    .Y(_05204_));
 sky130_fd_sc_hd__or2_1 _12448_ (.A(_05153_),
    .B(_05149_),
    .X(_05205_));
 sky130_fd_sc_hd__o2111a_1 _12449_ (.A1(_05153_),
    .A2(_05077_),
    .B1(_05081_),
    .C1(_05188_),
    .D1(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__a211oi_2 _12450_ (.A1(_05202_),
    .A2(_05203_),
    .B1(_05204_),
    .C1(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__and3b_1 _12451_ (.A_N(_05198_),
    .B(_05201_),
    .C(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__nand2_4 _12452_ (.A(_05185_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__buf_4 _12453_ (.A(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__nand2_1 _12454_ (.A(_05120_),
    .B(_05199_),
    .Y(_05211_));
 sky130_fd_sc_hd__xnor2_4 _12455_ (.A(_05126_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__and2_1 _12456_ (.A(_05097_),
    .B(_05099_),
    .X(_05213_));
 sky130_fd_sc_hd__o31a_1 _12457_ (.A1(_05105_),
    .A2(_05127_),
    .A3(_05131_),
    .B1(_05199_),
    .X(_05214_));
 sky130_fd_sc_hd__xor2_2 _12458_ (.A(_05213_),
    .B(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__nand2_1 _12459_ (.A(_05199_),
    .B(_05127_),
    .Y(_05216_));
 sky130_fd_sc_hd__xnor2_4 _12460_ (.A(_05105_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__o21a_1 _12461_ (.A1(_05105_),
    .A2(_05127_),
    .B1(_05199_),
    .X(_05218_));
 sky130_fd_sc_hd__xnor2_4 _12462_ (.A(_05131_),
    .B(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__or4b_1 _12463_ (.A(_05212_),
    .B(_05215_),
    .C(_05217_),
    .D_N(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__o21bai_2 _12464_ (.A1(_05167_),
    .A2(_05168_),
    .B1_N(_05174_),
    .Y(_05221_));
 sky130_fd_sc_hd__nand3b_1 _12465_ (.A_N(_05178_),
    .B(_05180_),
    .C(_05181_),
    .Y(_05222_));
 sky130_fd_sc_hd__xnor2_2 _12466_ (.A(_05161_),
    .B(_05183_),
    .Y(_05223_));
 sky130_fd_sc_hd__or4_4 _12467_ (.A(_05158_),
    .B(_05221_),
    .C(_05222_),
    .D(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__xnor2_2 _12468_ (.A(_05146_),
    .B(_05200_),
    .Y(_05225_));
 sky130_fd_sc_hd__or3b_2 _12469_ (.A(_05198_),
    .B(_05225_),
    .C_N(_05207_),
    .X(_05226_));
 sky130_fd_sc_hd__nand2_2 _12470_ (.A(_05199_),
    .B(_05132_),
    .Y(_05227_));
 sky130_fd_sc_hd__xor2_2 _12471_ (.A(_05094_),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__nand2_2 _12472_ (.A(_05087_),
    .B(_05089_),
    .Y(_05229_));
 sky130_fd_sc_hd__o21a_1 _12473_ (.A1(_05094_),
    .A2(_05132_),
    .B1(_05199_),
    .X(_05230_));
 sky130_fd_sc_hd__xor2_2 _12474_ (.A(_05229_),
    .B(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__nand2_1 _12475_ (.A(_05228_),
    .B(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__or4_1 _12476_ (.A(_05220_),
    .B(_05224_),
    .C(_05226_),
    .D(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__buf_2 _12477_ (.A(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__or2_2 _12478_ (.A(_05120_),
    .B(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__a21oi_2 _12479_ (.A1(_03489_),
    .A2(_05107_),
    .B1(_05109_),
    .Y(_05236_));
 sky130_fd_sc_hd__o21a_1 _12480_ (.A1(_05114_),
    .A2(_05119_),
    .B1(_05199_),
    .X(_05237_));
 sky130_fd_sc_hd__xnor2_4 _12481_ (.A(_05236_),
    .B(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__nand2_1 _12482_ (.A(_05116_),
    .B(_05199_),
    .Y(_05239_));
 sky130_fd_sc_hd__xnor2_1 _12483_ (.A(_05118_),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2_1 _12484_ (.A(_05119_),
    .B(_05199_),
    .Y(_05241_));
 sky130_fd_sc_hd__xnor2_4 _12485_ (.A(_05114_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__or4b_2 _12486_ (.A(_05238_),
    .B(_05240_),
    .C(_05242_),
    .D_N(_05116_),
    .X(_05243_));
 sky130_fd_sc_hd__or2_2 _12487_ (.A(_05234_),
    .B(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__or2_1 _12488_ (.A(_05215_),
    .B(_05219_),
    .X(_05245_));
 sky130_fd_sc_hd__or4_2 _12489_ (.A(_05224_),
    .B(_05226_),
    .C(_05232_),
    .D(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__xnor2_2 _12490_ (.A(_05229_),
    .B(_05230_),
    .Y(_05247_));
 sky130_fd_sc_hd__or4b_1 _12491_ (.A(_05189_),
    .B(_05225_),
    .C(_05231_),
    .D_N(_05192_),
    .X(_05248_));
 sky130_fd_sc_hd__or4b_1 _12492_ (.A(_05158_),
    .B(_05248_),
    .C(_05197_),
    .D_N(_05207_),
    .X(_05249_));
 sky130_fd_sc_hd__or4_1 _12493_ (.A(_05221_),
    .B(_05222_),
    .C(_05223_),
    .D(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__o41a_1 _12494_ (.A1(_05224_),
    .A2(_05226_),
    .A3(_05228_),
    .A4(_05247_),
    .B1(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__nand2_1 _12495_ (.A(_05202_),
    .B(_05203_),
    .Y(_05252_));
 sky130_fd_sc_hd__or2_1 _12496_ (.A(_05204_),
    .B(_05206_),
    .X(_05253_));
 sky130_fd_sc_hd__or2_1 _12497_ (.A(_05158_),
    .B(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__nor2_1 _12498_ (.A(_05223_),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__xnor2_1 _12499_ (.A(_05213_),
    .B(_05214_),
    .Y(_05256_));
 sky130_fd_sc_hd__and2_1 _12500_ (.A(_05202_),
    .B(_05203_),
    .X(_05257_));
 sky130_fd_sc_hd__xnor2_2 _12501_ (.A(_05094_),
    .B(_05227_),
    .Y(_05258_));
 sky130_fd_sc_hd__or3_1 _12502_ (.A(_05225_),
    .B(_05258_),
    .C(_05247_),
    .X(_05259_));
 sky130_fd_sc_hd__or4_1 _12503_ (.A(_05256_),
    .B(_05198_),
    .C(_05257_),
    .D(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__xor2_2 _12504_ (.A(_05118_),
    .B(_05239_),
    .X(_05261_));
 sky130_fd_sc_hd__or3_1 _12505_ (.A(_05238_),
    .B(_05242_),
    .C(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__or4_1 _12506_ (.A(_05220_),
    .B(_05193_),
    .C(_05259_),
    .D(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__or4_1 _12507_ (.A(_05197_),
    .B(_05257_),
    .C(_05254_),
    .D(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_1 _12508_ (.A(_05175_),
    .B(_05182_),
    .Y(_05265_));
 sky130_fd_sc_hd__a41o_1 _12509_ (.A1(_05252_),
    .A2(_05255_),
    .A3(_05260_),
    .A4(_05264_),
    .B1(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__and3_1 _12510_ (.A(_05246_),
    .B(_05251_),
    .C(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__and3_1 _12511_ (.A(_05235_),
    .B(_05244_),
    .C(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__buf_2 _12512_ (.A(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__clkbuf_4 _12513_ (.A(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__buf_2 _12514_ (.A(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__a21oi_1 _12515_ (.A1(_05120_),
    .A2(_05243_),
    .B1(_05234_),
    .Y(_05272_));
 sky130_fd_sc_hd__or2b_1 _12516_ (.A(_05272_),
    .B_N(_05267_),
    .X(_05273_));
 sky130_fd_sc_hd__buf_4 _12517_ (.A(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__inv_2 _12518_ (.A(_05242_),
    .Y(_05275_));
 sky130_fd_sc_hd__o31a_2 _12519_ (.A1(_05234_),
    .A2(_05238_),
    .A3(_05275_),
    .B1(_05246_),
    .X(_05276_));
 sky130_fd_sc_hd__or4_1 _12520_ (.A(_05221_),
    .B(_05222_),
    .C(_05223_),
    .D(_05254_),
    .X(_05277_));
 sky130_fd_sc_hd__or4_2 _12521_ (.A(_05198_),
    .B(_05201_),
    .C(_05257_),
    .D(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__inv_2 _12522_ (.A(_05238_),
    .Y(_05279_));
 sky130_fd_sc_hd__or2_1 _12523_ (.A(_05189_),
    .B(_05192_),
    .X(_05280_));
 sky130_fd_sc_hd__o41a_1 _12524_ (.A1(_05220_),
    .A2(_05193_),
    .A3(_05279_),
    .A4(_05259_),
    .B1(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__o21a_1 _12525_ (.A1(_05197_),
    .A2(_05281_),
    .B1(_05207_),
    .X(_05282_));
 sky130_fd_sc_hd__o22a_1 _12526_ (.A1(_05221_),
    .A2(_05182_),
    .B1(_05224_),
    .B2(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__o211a_1 _12527_ (.A1(_05277_),
    .A2(_05260_),
    .B1(_05278_),
    .C1(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__and3_1 _12528_ (.A(_05235_),
    .B(_05276_),
    .C(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__and4_1 _12529_ (.A(_05185_),
    .B(_05208_),
    .C(_05258_),
    .D(_05231_),
    .X(_05286_));
 sky130_fd_sc_hd__nor4_1 _12530_ (.A(_05221_),
    .B(_05222_),
    .C(_05223_),
    .D(_05254_),
    .Y(_05287_));
 sky130_fd_sc_hd__a31o_1 _12531_ (.A1(_05178_),
    .A2(_05180_),
    .A3(_05181_),
    .B1(_05174_),
    .X(_05288_));
 sky130_fd_sc_hd__a41o_1 _12532_ (.A1(_05158_),
    .A2(_05175_),
    .A3(_05182_),
    .A4(_05184_),
    .B1(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a21o_1 _12533_ (.A1(_05257_),
    .A2(_05287_),
    .B1(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__or2b_1 _12534_ (.A(_05197_),
    .B_N(_05189_),
    .X(_05291_));
 sky130_fd_sc_hd__o21ai_1 _12535_ (.A1(_05198_),
    .A2(_05201_),
    .B1(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__and3_1 _12536_ (.A(_05252_),
    .B(_05287_),
    .C(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__inv_2 _12537_ (.A(_05217_),
    .Y(_05294_));
 sky130_fd_sc_hd__and4_1 _12538_ (.A(_05212_),
    .B(_05256_),
    .C(_05219_),
    .D(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__or4b_1 _12539_ (.A(_05224_),
    .B(_05226_),
    .C(_05232_),
    .D_N(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__nor4b_4 _12540_ (.A(_05286_),
    .B(_05290_),
    .C(_05293_),
    .D_N(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__and3_1 _12541_ (.A(_05244_),
    .B(_05276_),
    .C(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_2 _12542_ (.A(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__or3_2 _12543_ (.A(_05274_),
    .B(_05285_),
    .C(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__nor2_4 _12544_ (.A(_05120_),
    .B(_05234_),
    .Y(_05301_));
 sky130_fd_sc_hd__o31ai_4 _12545_ (.A1(_05234_),
    .A2(_05238_),
    .A3(_05275_),
    .B1(_05246_),
    .Y(_05302_));
 sky130_fd_sc_hd__or3b_1 _12546_ (.A(_05301_),
    .B(_05302_),
    .C_N(_05284_),
    .X(_05303_));
 sky130_fd_sc_hd__buf_2 _12547_ (.A(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__nor2_2 _12548_ (.A(_05234_),
    .B(_05243_),
    .Y(_05305_));
 sky130_fd_sc_hd__or4b_2 _12549_ (.A(_05286_),
    .B(_05290_),
    .C(_05293_),
    .D_N(_05296_),
    .X(_05306_));
 sky130_fd_sc_hd__or3_1 _12550_ (.A(_05305_),
    .B(_05302_),
    .C(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__a21o_1 _12551_ (.A1(_05304_),
    .A2(_05307_),
    .B1(_05269_),
    .X(_05308_));
 sky130_fd_sc_hd__nand2_1 _12552_ (.A(_05300_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__clkbuf_4 _12553_ (.A(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__clkbuf_4 _12554_ (.A(_05307_),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _12555_ (.A0(_05212_),
    .A1(_05217_),
    .S(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__clkbuf_4 _12556_ (.A(_05299_),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _12557_ (.A0(_05238_),
    .A1(_05242_),
    .S(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__xnor2_4 _12558_ (.A(_05304_),
    .B(_05299_),
    .Y(_05315_));
 sky130_fd_sc_hd__mux2_1 _12559_ (.A0(_05312_),
    .A1(_05314_),
    .S(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__o211a_1 _12560_ (.A1(_05198_),
    .A2(_05225_),
    .B1(_05252_),
    .C1(_05287_),
    .X(_05317_));
 sky130_fd_sc_hd__o21bai_1 _12561_ (.A1(_05277_),
    .A2(_05260_),
    .B1_N(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__and3b_1 _12562_ (.A_N(_05318_),
    .B(_05246_),
    .C(_05251_),
    .X(_05319_));
 sky130_fd_sc_hd__clkbuf_4 _12563_ (.A(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__xnor2_1 _12564_ (.A(_05269_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__a21boi_4 _12565_ (.A1(_05321_),
    .A2(_05300_),
    .B1_N(_05278_),
    .Y(_05322_));
 sky130_fd_sc_hd__nor2_4 _12566_ (.A(_05209_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__clkbuf_4 _12567_ (.A(_05313_),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_4 _12568_ (.A(_05304_),
    .X(_05325_));
 sky130_fd_sc_hd__mux4_1 _12569_ (.A0(_05256_),
    .A1(_05228_),
    .A2(_05231_),
    .A3(_05219_),
    .S0(_05324_),
    .S1(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__nand2_1 _12570_ (.A(_05310_),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__o211a_1 _12571_ (.A1(_05310_),
    .A2(_05316_),
    .B1(_05323_),
    .C1(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__clkbuf_4 _12572_ (.A(_05285_),
    .X(_05329_));
 sky130_fd_sc_hd__xnor2_1 _12573_ (.A(_05329_),
    .B(_05299_),
    .Y(_05330_));
 sky130_fd_sc_hd__mux2_1 _12574_ (.A0(_05116_),
    .A1(_05240_),
    .S(_05311_),
    .X(_05331_));
 sky130_fd_sc_hd__and2_1 _12575_ (.A(_05330_),
    .B(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__clkbuf_4 _12576_ (.A(_05321_),
    .X(_05333_));
 sky130_fd_sc_hd__a21bo_2 _12577_ (.A1(_05333_),
    .A2(_05300_),
    .B1_N(_05278_),
    .X(_05334_));
 sky130_fd_sc_hd__nor2_1 _12578_ (.A(_05210_),
    .B(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__or4b_1 _12579_ (.A(_05305_),
    .B(_05302_),
    .C(_05306_),
    .D_N(_05189_),
    .X(_05336_));
 sky130_fd_sc_hd__a31o_1 _12580_ (.A1(_05244_),
    .A2(_05276_),
    .A3(_05297_),
    .B1(_05192_),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_4 _12581_ (.A(_05304_),
    .X(_05338_));
 sky130_fd_sc_hd__a21oi_1 _12582_ (.A1(_05336_),
    .A2(_05337_),
    .B1(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__a31o_1 _12583_ (.A1(_05244_),
    .A2(_05276_),
    .A3(_05297_),
    .B1(_05231_),
    .X(_05340_));
 sky130_fd_sc_hd__or4_1 _12584_ (.A(_05201_),
    .B(_05305_),
    .C(_05302_),
    .D(_05306_),
    .X(_05341_));
 sky130_fd_sc_hd__a21oi_1 _12585_ (.A1(_05340_),
    .A2(_05341_),
    .B1(_05329_),
    .Y(_05342_));
 sky130_fd_sc_hd__or2_1 _12586_ (.A(_05339_),
    .B(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(_05158_),
    .A1(_05253_),
    .S(_05311_),
    .X(_05344_));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(_05197_),
    .A1(_05257_),
    .S(_05313_),
    .X(_05345_));
 sky130_fd_sc_hd__mux2_1 _12589_ (.A0(_05344_),
    .A1(_05345_),
    .S(_05338_),
    .X(_05346_));
 sky130_fd_sc_hd__clkbuf_4 _12590_ (.A(_05274_),
    .X(_05347_));
 sky130_fd_sc_hd__nand2_1 _12591_ (.A(_05180_),
    .B(_05181_),
    .Y(_05348_));
 sky130_fd_sc_hd__clkbuf_4 _12592_ (.A(_05311_),
    .X(_05349_));
 sky130_fd_sc_hd__mux2_1 _12593_ (.A0(_05178_),
    .A1(_05223_),
    .S(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(_05348_),
    .A1(_05350_),
    .S(_05325_),
    .X(_05351_));
 sky130_fd_sc_hd__a221o_1 _12595_ (.A1(_05317_),
    .A2(_05343_),
    .B1(_05346_),
    .B2(_05347_),
    .C1(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__a31o_1 _12596_ (.A1(_05310_),
    .A2(_05332_),
    .A3(_05335_),
    .B1(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__nor2_1 _12597_ (.A(_05328_),
    .B(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__clkbuf_4 _12598_ (.A(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__xnor2_4 _12599_ (.A(_05274_),
    .B(_05320_),
    .Y(_05356_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(_05253_),
    .A1(_05257_),
    .S(_05311_),
    .X(_05357_));
 sky130_fd_sc_hd__mux2_1 _12601_ (.A0(_05189_),
    .A1(_05197_),
    .S(_05313_),
    .X(_05358_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(_05357_),
    .A1(_05358_),
    .S(_05325_),
    .X(_05359_));
 sky130_fd_sc_hd__clkinv_2 _12603_ (.A(_05192_),
    .Y(_05360_));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(_05360_),
    .A1(_05225_),
    .S(_05311_),
    .X(_05361_));
 sky130_fd_sc_hd__mux2_1 _12605_ (.A0(_05258_),
    .A1(_05247_),
    .S(_05313_),
    .X(_05362_));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(_05361_),
    .A1(_05362_),
    .S(_05338_),
    .X(_05363_));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(_05359_),
    .A1(_05363_),
    .S(_05270_),
    .X(_05364_));
 sky130_fd_sc_hd__mux2_1 _12608_ (.A0(_05158_),
    .A1(_05223_),
    .S(_05313_),
    .X(_05365_));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(_05178_),
    .A1(_05348_),
    .S(_05324_),
    .X(_05366_));
 sky130_fd_sc_hd__clkbuf_4 _12610_ (.A(_05329_),
    .X(_05367_));
 sky130_fd_sc_hd__mux2_1 _12611_ (.A0(_05365_),
    .A1(_05366_),
    .S(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__nor2_4 _12612_ (.A(_05224_),
    .B(_05226_),
    .Y(_05369_));
 sky130_fd_sc_hd__a211o_1 _12613_ (.A1(_05356_),
    .A2(_05364_),
    .B1(_05368_),
    .C1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__nand2_1 _12614_ (.A(_05116_),
    .B(_05311_),
    .Y(_05371_));
 sky130_fd_sc_hd__nand2_2 _12615_ (.A(_05269_),
    .B(_05338_),
    .Y(_05372_));
 sky130_fd_sc_hd__clkbuf_4 _12616_ (.A(_05335_),
    .X(_05373_));
 sky130_fd_sc_hd__o21ai_2 _12617_ (.A1(_05371_),
    .A2(_05372_),
    .B1(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__and2_1 _12618_ (.A(_05300_),
    .B(_05308_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_4 _12619_ (.A(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__mux2_1 _12620_ (.A0(_05242_),
    .A1(_05240_),
    .S(_05313_),
    .X(_05377_));
 sky130_fd_sc_hd__a31o_1 _12621_ (.A1(_05244_),
    .A2(_05276_),
    .A3(_05297_),
    .B1(_05212_),
    .X(_05378_));
 sky130_fd_sc_hd__o21a_1 _12622_ (.A1(_05238_),
    .A2(_05349_),
    .B1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_4 _12623_ (.A(_05330_),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _12624_ (.A0(_05377_),
    .A1(_05379_),
    .S(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__inv_2 _12625_ (.A(_05219_),
    .Y(_05382_));
 sky130_fd_sc_hd__a31o_1 _12626_ (.A1(_05244_),
    .A2(_05276_),
    .A3(_05297_),
    .B1(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__or4_1 _12627_ (.A(_05217_),
    .B(_05305_),
    .C(_05302_),
    .D(_05306_),
    .X(_05384_));
 sky130_fd_sc_hd__nand2_1 _12628_ (.A(_05383_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__or4_1 _12629_ (.A(_05215_),
    .B(_05305_),
    .C(_05302_),
    .D(_05306_),
    .X(_05386_));
 sky130_fd_sc_hd__o21ai_1 _12630_ (.A1(_05258_),
    .A2(_05324_),
    .B1(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(_05385_),
    .A1(_05387_),
    .S(_05380_),
    .X(_05388_));
 sky130_fd_sc_hd__nor2_1 _12632_ (.A(_05376_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_4 _12633_ (.A(_05369_),
    .B(_05334_),
    .Y(_05390_));
 sky130_fd_sc_hd__a211o_1 _12634_ (.A1(_05376_),
    .A2(_05381_),
    .B1(_05389_),
    .C1(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__nand3_4 _12635_ (.A(_05370_),
    .B(_05374_),
    .C(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__and3_1 _12636_ (.A(_05338_),
    .B(_05383_),
    .C(_05386_),
    .X(_05393_));
 sky130_fd_sc_hd__a21o_1 _12637_ (.A1(_05367_),
    .A2(_05362_),
    .B1(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__nor2_4 _12638_ (.A(_05274_),
    .B(_05329_),
    .Y(_05395_));
 sky130_fd_sc_hd__mux2_1 _12639_ (.A0(_05238_),
    .A1(_05242_),
    .S(_05311_),
    .X(_05396_));
 sky130_fd_sc_hd__and4_1 _12640_ (.A(_05269_),
    .B(_05329_),
    .C(_05378_),
    .D(_05384_),
    .X(_05397_));
 sky130_fd_sc_hd__a211o_1 _12641_ (.A1(_05395_),
    .A2(_05396_),
    .B1(_05397_),
    .C1(_05333_),
    .X(_05398_));
 sky130_fd_sc_hd__a21oi_1 _12642_ (.A1(_05347_),
    .A2(_05394_),
    .B1(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__mux2_1 _12643_ (.A0(_05358_),
    .A1(_05361_),
    .S(_05338_),
    .X(_05400_));
 sky130_fd_sc_hd__nor2_1 _12644_ (.A(_05347_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__o2bb2a_1 _12645_ (.A1_N(_05330_),
    .A2_N(_05377_),
    .B1(_05371_),
    .B2(_05325_),
    .X(_05402_));
 sky130_fd_sc_hd__or4_1 _12646_ (.A(_05209_),
    .B(_05376_),
    .C(_05322_),
    .D(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__o31a_4 _12647_ (.A1(_05369_),
    .A2(_05399_),
    .A3(_05401_),
    .B1(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__mux2_1 _12648_ (.A0(_05256_),
    .A1(_05228_),
    .S(_05313_),
    .X(_05405_));
 sky130_fd_sc_hd__or4_1 _12649_ (.A(_05219_),
    .B(_05305_),
    .C(_05302_),
    .D(_05306_),
    .X(_05406_));
 sky130_fd_sc_hd__o211a_1 _12650_ (.A1(_05294_),
    .A2(_05313_),
    .B1(_05406_),
    .C1(_05304_),
    .X(_05407_));
 sky130_fd_sc_hd__a211o_1 _12651_ (.A1(_05329_),
    .A2(_05405_),
    .B1(_05407_),
    .C1(_05269_),
    .X(_05408_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(_05212_),
    .A1(_05238_),
    .S(_05311_),
    .X(_05409_));
 sky130_fd_sc_hd__nor2_2 _12653_ (.A(_05274_),
    .B(_05338_),
    .Y(_05410_));
 sky130_fd_sc_hd__o211a_1 _12654_ (.A1(_05242_),
    .A2(_05311_),
    .B1(_05338_),
    .C1(_05269_),
    .X(_05411_));
 sky130_fd_sc_hd__nand2_1 _12655_ (.A(_05261_),
    .B(_05349_),
    .Y(_05412_));
 sky130_fd_sc_hd__a221oi_1 _12656_ (.A1(_05409_),
    .A2(_05410_),
    .B1(_05411_),
    .B2(_05412_),
    .C1(_05333_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand2_2 _12657_ (.A(_05269_),
    .B(_05320_),
    .Y(_05414_));
 sky130_fd_sc_hd__o31a_1 _12658_ (.A1(_05414_),
    .A2(_05339_),
    .A3(_05342_),
    .B1(_05209_),
    .X(_05415_));
 sky130_fd_sc_hd__a21bo_1 _12659_ (.A1(_05408_),
    .A2(_05413_),
    .B1_N(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__or2_2 _12660_ (.A(_05414_),
    .B(_05363_),
    .X(_05417_));
 sky130_fd_sc_hd__a21o_1 _12661_ (.A1(_05378_),
    .A2(_05384_),
    .B1(_05329_),
    .X(_05418_));
 sky130_fd_sc_hd__a21o_1 _12662_ (.A1(_05383_),
    .A2(_05386_),
    .B1(_05338_),
    .X(_05419_));
 sky130_fd_sc_hd__a21o_1 _12663_ (.A1(_05418_),
    .A2(_05419_),
    .B1(_05270_),
    .X(_05420_));
 sky130_fd_sc_hd__nand2_1 _12664_ (.A(_05269_),
    .B(_05329_),
    .Y(_05421_));
 sky130_fd_sc_hd__or2_1 _12665_ (.A(_05421_),
    .B(_05396_),
    .X(_05422_));
 sky130_fd_sc_hd__o211ai_1 _12666_ (.A1(_05261_),
    .A2(_05349_),
    .B1(_05371_),
    .C1(_05395_),
    .Y(_05423_));
 sky130_fd_sc_hd__a31o_2 _12667_ (.A1(_05420_),
    .A2(_05422_),
    .A3(_05423_),
    .B1(_05333_),
    .X(_05424_));
 sky130_fd_sc_hd__nand4b_4 _12668_ (.A_N(_05416_),
    .B(_05417_),
    .C(_05424_),
    .D(_05209_),
    .Y(_05425_));
 sky130_fd_sc_hd__a211o_1 _12669_ (.A1(_05367_),
    .A2(_05405_),
    .B1(_05407_),
    .C1(_05274_),
    .X(_05426_));
 sky130_fd_sc_hd__and3_1 _12670_ (.A(_05338_),
    .B(_05340_),
    .C(_05341_),
    .X(_05427_));
 sky130_fd_sc_hd__and3_1 _12671_ (.A(_05329_),
    .B(_05336_),
    .C(_05337_),
    .X(_05428_));
 sky130_fd_sc_hd__o31a_1 _12672_ (.A1(_05270_),
    .A2(_05427_),
    .A3(_05428_),
    .B1(_05356_),
    .X(_05429_));
 sky130_fd_sc_hd__nand2_1 _12673_ (.A(_05426_),
    .B(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__or2_1 _12674_ (.A(_05414_),
    .B(_05346_),
    .X(_05431_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(_05316_),
    .A1(_05332_),
    .S(_05375_),
    .X(_05432_));
 sky130_fd_sc_hd__a32oi_4 _12676_ (.A1(_05209_),
    .A2(_05430_),
    .A3(_05431_),
    .B1(_05323_),
    .B2(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__mux2_1 _12677_ (.A0(_05314_),
    .A1(_05331_),
    .S(_05315_),
    .X(_05434_));
 sky130_fd_sc_hd__a21o_1 _12678_ (.A1(_05340_),
    .A2(_05341_),
    .B1(_05325_),
    .X(_05435_));
 sky130_fd_sc_hd__o211ai_1 _12679_ (.A1(_05367_),
    .A2(_05405_),
    .B1(_05435_),
    .C1(_05274_),
    .Y(_05436_));
 sky130_fd_sc_hd__o21ai_1 _12680_ (.A1(_05294_),
    .A2(_05313_),
    .B1(_05406_),
    .Y(_05437_));
 sky130_fd_sc_hd__o22a_1 _12681_ (.A1(_05372_),
    .A2(_05409_),
    .B1(_05421_),
    .B2(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__a21o_1 _12682_ (.A1(_05436_),
    .A2(_05438_),
    .B1(_05333_),
    .X(_05439_));
 sky130_fd_sc_hd__nand2_1 _12683_ (.A(_05336_),
    .B(_05337_),
    .Y(_05440_));
 sky130_fd_sc_hd__mux2_1 _12684_ (.A0(_05440_),
    .A1(_05345_),
    .S(_05329_),
    .X(_05441_));
 sky130_fd_sc_hd__o21a_1 _12685_ (.A1(_05414_),
    .A2(_05441_),
    .B1(_05209_),
    .X(_05442_));
 sky130_fd_sc_hd__a32oi_4 _12686_ (.A1(_05310_),
    .A2(_05323_),
    .A3(_05434_),
    .B1(_05439_),
    .B2(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__a31o_1 _12687_ (.A1(_05270_),
    .A2(_05418_),
    .A3(_05419_),
    .B1(_05333_),
    .X(_05444_));
 sky130_fd_sc_hd__a21o_1 _12688_ (.A1(_05347_),
    .A2(_05363_),
    .B1(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__or2_1 _12689_ (.A(_05414_),
    .B(_05359_),
    .X(_05446_));
 sky130_fd_sc_hd__nor2_2 _12690_ (.A(_05270_),
    .B(_05367_),
    .Y(_05447_));
 sky130_fd_sc_hd__a32o_2 _12691_ (.A1(_05116_),
    .A2(_05447_),
    .A3(_05349_),
    .B1(_05310_),
    .B2(_05381_),
    .X(_05448_));
 sky130_fd_sc_hd__a32oi_4 _12692_ (.A1(_05210_),
    .A2(_05445_),
    .A3(_05446_),
    .B1(_05323_),
    .B2(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__a2111o_4 _12693_ (.A1(_05404_),
    .A2(_05425_),
    .B1(_05433_),
    .C1(_05443_),
    .D1(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__or2_1 _12694_ (.A(_05309_),
    .B(_05402_),
    .X(_05451_));
 sky130_fd_sc_hd__nor2_1 _12695_ (.A(_05380_),
    .B(_05379_),
    .Y(_05452_));
 sky130_fd_sc_hd__a211o_1 _12696_ (.A1(_05380_),
    .A2(_05385_),
    .B1(_05452_),
    .C1(_05376_),
    .X(_05453_));
 sky130_fd_sc_hd__a21oi_1 _12697_ (.A1(_05451_),
    .A2(_05453_),
    .B1(_05390_),
    .Y(_05454_));
 sky130_fd_sc_hd__a22o_1 _12698_ (.A1(_05357_),
    .A2(_05395_),
    .B1(_05410_),
    .B2(_05365_),
    .X(_05455_));
 sky130_fd_sc_hd__mux2_1 _12699_ (.A0(_05394_),
    .A1(_05400_),
    .S(_05274_),
    .X(_05456_));
 sky130_fd_sc_hd__nand2_1 _12700_ (.A(_05356_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__nor3b_2 _12701_ (.A(_05454_),
    .B(_05455_),
    .C_N(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__or2_1 _12702_ (.A(_05270_),
    .B(_05441_),
    .X(_05459_));
 sky130_fd_sc_hd__o211ai_1 _12703_ (.A1(_05367_),
    .A2(_05405_),
    .B1(_05435_),
    .C1(_05270_),
    .Y(_05460_));
 sky130_fd_sc_hd__mux4_1 _12704_ (.A0(_05212_),
    .A1(_05215_),
    .A2(_05382_),
    .A3(_05217_),
    .S0(_05349_),
    .S1(_05367_),
    .X(_05461_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(_05461_),
    .A1(_05434_),
    .S(_05376_),
    .X(_05462_));
 sky130_fd_sc_hd__and2_1 _12706_ (.A(_05325_),
    .B(_05344_),
    .X(_05463_));
 sky130_fd_sc_hd__a221o_1 _12707_ (.A1(_05367_),
    .A2(_05350_),
    .B1(_05462_),
    .B2(_05323_),
    .C1(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__a31o_2 _12708_ (.A1(_05356_),
    .A2(_05459_),
    .A3(_05460_),
    .B1(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__a21bo_1 _12709_ (.A1(_05450_),
    .A2(_05458_),
    .B1_N(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__buf_4 _12710_ (.A(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__or2_1 _12711_ (.A(_05392_),
    .B(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__clkbuf_4 _12712_ (.A(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__xor2_1 _12713_ (.A(_05355_),
    .B(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__buf_2 _12714_ (.A(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__buf_2 _12715_ (.A(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__buf_2 _12716_ (.A(_05443_),
    .X(_05473_));
 sky130_fd_sc_hd__xor2_4 _12717_ (.A(_05392_),
    .B(_05467_),
    .X(_05474_));
 sky130_fd_sc_hd__nor2_1 _12718_ (.A(_05473_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__clkbuf_4 _12719_ (.A(_05323_),
    .X(_05476_));
 sky130_fd_sc_hd__a32o_2 _12720_ (.A1(_05210_),
    .A2(_05430_),
    .A3(_05431_),
    .B1(_05476_),
    .B2(_05432_),
    .X(_05477_));
 sky130_fd_sc_hd__or3b_1 _12721_ (.A(_05454_),
    .B(_05455_),
    .C_N(_05457_),
    .X(_05478_));
 sky130_fd_sc_hd__clkbuf_4 _12722_ (.A(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__xnor2_4 _12723_ (.A(_05450_),
    .B(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2_1 _12724_ (.A(_05477_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__or3b_1 _12725_ (.A(_05465_),
    .B(_05479_),
    .C_N(_05450_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_2 _12726_ (.A(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__clkbuf_4 _12727_ (.A(_05449_),
    .X(_05484_));
 sky130_fd_sc_hd__a21oi_2 _12728_ (.A1(_05467_),
    .A2(_05483_),
    .B1(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__xnor2_1 _12729_ (.A(_05481_),
    .B(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__xnor2_1 _12730_ (.A(_05475_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__nor2_4 _12731_ (.A(_05443_),
    .B(_05404_),
    .Y(_05488_));
 sky130_fd_sc_hd__nor2_4 _12732_ (.A(_05443_),
    .B(_05425_),
    .Y(_05489_));
 sky130_fd_sc_hd__and3_1 _12733_ (.A(_05443_),
    .B(_05404_),
    .C(_05425_),
    .X(_05490_));
 sky130_fd_sc_hd__buf_2 _12734_ (.A(_05465_),
    .X(_05491_));
 sky130_fd_sc_hd__o31a_2 _12735_ (.A1(_05488_),
    .A2(_05489_),
    .A3(_05490_),
    .B1(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__clkbuf_4 _12736_ (.A(_05458_),
    .X(_05493_));
 sky130_fd_sc_hd__a32o_4 _12737_ (.A1(_05210_),
    .A2(_05445_),
    .A3(_05446_),
    .B1(_05323_),
    .B2(_05448_),
    .X(_05494_));
 sky130_fd_sc_hd__a211o_4 _12738_ (.A1(_05404_),
    .A2(_05425_),
    .B1(_05449_),
    .C1(_05443_),
    .X(_05495_));
 sky130_fd_sc_hd__o31a_2 _12739_ (.A1(_05494_),
    .A2(_05488_),
    .A3(_05489_),
    .B1(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__nor2_1 _12740_ (.A(_05493_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__xor2_1 _12741_ (.A(_05492_),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__nor2_2 _12742_ (.A(_05495_),
    .B(_05433_),
    .Y(_05499_));
 sky130_fd_sc_hd__a22o_1 _12743_ (.A1(_05492_),
    .A2(_05497_),
    .B1(_05498_),
    .B2(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__and2b_1 _12744_ (.A_N(_05487_),
    .B(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__xnor2_1 _12745_ (.A(_05450_),
    .B(_05458_),
    .Y(_05502_));
 sky130_fd_sc_hd__clkbuf_4 _12746_ (.A(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__nor2_1 _12747_ (.A(_05473_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__buf_2 _12748_ (.A(_05404_),
    .X(_05505_));
 sky130_fd_sc_hd__nor2_1 _12749_ (.A(_05505_),
    .B(_05474_),
    .Y(_05506_));
 sky130_fd_sc_hd__nand2_1 _12750_ (.A(_05494_),
    .B(_05480_),
    .Y(_05507_));
 sky130_fd_sc_hd__a21oi_1 _12751_ (.A1(_05467_),
    .A2(_05483_),
    .B1(_05473_),
    .Y(_05508_));
 sky130_fd_sc_hd__xnor2_1 _12752_ (.A(_05507_),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__a22oi_2 _12753_ (.A1(_05485_),
    .A2(_05504_),
    .B1(_05506_),
    .B2(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__xnor2_1 _12754_ (.A(_05500_),
    .B(_05487_),
    .Y(_05511_));
 sky130_fd_sc_hd__and2b_1 _12755_ (.A_N(_05510_),
    .B(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__or2_1 _12756_ (.A(_05505_),
    .B(_05471_),
    .X(_05513_));
 sky130_fd_sc_hd__nand2_1 _12757_ (.A(_05380_),
    .B(_05331_),
    .Y(_05514_));
 sky130_fd_sc_hd__o31a_4 _12758_ (.A1(_05376_),
    .A2(_05390_),
    .A3(_05514_),
    .B1(_05416_),
    .X(_05515_));
 sky130_fd_sc_hd__buf_2 _12759_ (.A(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__o21ai_4 _12760_ (.A1(_05355_),
    .A2(_05469_),
    .B1(_05235_),
    .Y(_05517_));
 sky130_fd_sc_hd__or2_1 _12761_ (.A(_05516_),
    .B(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__or2_1 _12762_ (.A(_05513_),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__or2_1 _12763_ (.A(_05505_),
    .B(_05517_),
    .X(_05520_));
 sky130_fd_sc_hd__or2_1 _12764_ (.A(_05473_),
    .B(_05471_),
    .X(_05521_));
 sky130_fd_sc_hd__xor2_1 _12765_ (.A(_05520_),
    .B(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__xnor2_1 _12766_ (.A(_05519_),
    .B(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__o21a_1 _12767_ (.A1(_05501_),
    .A2(_05512_),
    .B1(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__nor2_1 _12768_ (.A(_05505_),
    .B(_05470_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand3_4 _12769_ (.A(_05210_),
    .B(_05424_),
    .C(_05417_),
    .Y(_05526_));
 sky130_fd_sc_hd__clkbuf_4 _12770_ (.A(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__nor2_1 _12771_ (.A(_05527_),
    .B(_05471_),
    .Y(_05528_));
 sky130_fd_sc_hd__or3b_1 _12772_ (.A(_05525_),
    .B(_05518_),
    .C_N(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__nor3_1 _12773_ (.A(_05523_),
    .B(_05501_),
    .C(_05512_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_1 _12774_ (.A(_05524_),
    .B(_05530_),
    .Y(_05531_));
 sky130_fd_sc_hd__and2b_1 _12775_ (.A_N(_05529_),
    .B(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__or2_1 _12776_ (.A(_05524_),
    .B(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__and3_1 _12777_ (.A(_05210_),
    .B(_05424_),
    .C(_05417_),
    .X(_05534_));
 sky130_fd_sc_hd__xnor2_2 _12778_ (.A(_05534_),
    .B(_05515_),
    .Y(_05535_));
 sky130_fd_sc_hd__xnor2_4 _12779_ (.A(_05404_),
    .B(_05425_),
    .Y(_05536_));
 sky130_fd_sc_hd__or4_1 _12780_ (.A(_05301_),
    .B(_05354_),
    .C(_05535_),
    .D(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__xnor2_4 _12781_ (.A(_05526_),
    .B(_05515_),
    .Y(_05538_));
 sky130_fd_sc_hd__a2bb2o_1 _12782_ (.A1_N(_05355_),
    .A2_N(_05536_),
    .B1(_05538_),
    .B2(_05235_),
    .X(_05539_));
 sky130_fd_sc_hd__nand2_1 _12783_ (.A(_05537_),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__nor2_1 _12784_ (.A(_05392_),
    .B(_05536_),
    .Y(_05541_));
 sky130_fd_sc_hd__mux2_1 _12785_ (.A0(_05515_),
    .A1(_05534_),
    .S(_05354_),
    .X(_05542_));
 sky130_fd_sc_hd__o2bb2a_1 _12786_ (.A1_N(_05541_),
    .A2_N(_05542_),
    .B1(_05355_),
    .B2(_05425_),
    .X(_05543_));
 sky130_fd_sc_hd__xnor2_2 _12787_ (.A(_05540_),
    .B(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__nand2_1 _12788_ (.A(_05495_),
    .B(_05433_),
    .Y(_05545_));
 sky130_fd_sc_hd__and2_1 _12789_ (.A(_05450_),
    .B(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__nor2_1 _12790_ (.A(_05493_),
    .B(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__nor2_1 _12791_ (.A(_05392_),
    .B(_05496_),
    .Y(_05548_));
 sky130_fd_sc_hd__o31ai_4 _12792_ (.A1(_05494_),
    .A2(_05488_),
    .A3(_05489_),
    .B1(_05495_),
    .Y(_05549_));
 sky130_fd_sc_hd__nor3_1 _12793_ (.A(_05488_),
    .B(_05489_),
    .C(_05490_),
    .Y(_05550_));
 sky130_fd_sc_hd__clkbuf_4 _12794_ (.A(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__o2bb2a_1 _12795_ (.A1_N(_05491_),
    .A2_N(_05549_),
    .B1(_05551_),
    .B2(_05392_),
    .X(_05552_));
 sky130_fd_sc_hd__a21oi_1 _12796_ (.A1(_05492_),
    .A2(_05548_),
    .B1(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__xnor2_1 _12797_ (.A(_05547_),
    .B(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__xor2_2 _12798_ (.A(_05544_),
    .B(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__xnor2_1 _12799_ (.A(_05541_),
    .B(_05542_),
    .Y(_05556_));
 sky130_fd_sc_hd__and4b_2 _12800_ (.A_N(_05416_),
    .B(_05417_),
    .C(_05424_),
    .D(_05210_),
    .X(_05557_));
 sky130_fd_sc_hd__or2_1 _12801_ (.A(_05404_),
    .B(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(_05505_),
    .B(_05557_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_1 _12803_ (.A(_05558_),
    .B(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__and2_1 _12804_ (.A(_05491_),
    .B(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__or2_1 _12805_ (.A(_05354_),
    .B(_05526_),
    .X(_05562_));
 sky130_fd_sc_hd__or2_1 _12806_ (.A(_05392_),
    .B(_05535_),
    .X(_05563_));
 sky130_fd_sc_hd__xor2_1 _12807_ (.A(_05562_),
    .B(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__nor2_1 _12808_ (.A(_05562_),
    .B(_05563_),
    .Y(_05565_));
 sky130_fd_sc_hd__a21oi_1 _12809_ (.A1(_05561_),
    .A2(_05564_),
    .B1(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__xnor2_1 _12810_ (.A(_05556_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__xnor2_1 _12811_ (.A(_05499_),
    .B(_05498_),
    .Y(_05568_));
 sky130_fd_sc_hd__or2_1 _12812_ (.A(_05556_),
    .B(_05566_),
    .X(_05569_));
 sky130_fd_sc_hd__o21a_1 _12813_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__xnor2_1 _12814_ (.A(_05555_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__xnor2_1 _12815_ (.A(_05510_),
    .B(_05511_),
    .Y(_05572_));
 sky130_fd_sc_hd__or2b_1 _12816_ (.A(_05570_),
    .B_N(_05555_),
    .X(_05573_));
 sky130_fd_sc_hd__a21bo_1 _12817_ (.A1(_05571_),
    .A2(_05572_),
    .B1_N(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__nand2_1 _12818_ (.A(_05560_),
    .B(_05537_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand2_2 _12819_ (.A(_05450_),
    .B(_05545_),
    .Y(_05576_));
 sky130_fd_sc_hd__nand2_1 _12820_ (.A(_05491_),
    .B(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__nor2_1 _12821_ (.A(_05355_),
    .B(_05551_),
    .Y(_05578_));
 sky130_fd_sc_hd__xnor2_1 _12822_ (.A(_05548_),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__or2_1 _12823_ (.A(_05577_),
    .B(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__nand2_1 _12824_ (.A(_05577_),
    .B(_05579_),
    .Y(_05581_));
 sky130_fd_sc_hd__nand2_1 _12825_ (.A(_05580_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__xor2_1 _12826_ (.A(_05575_),
    .B(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__or2_1 _12827_ (.A(_05544_),
    .B(_05554_),
    .X(_05584_));
 sky130_fd_sc_hd__o21ai_2 _12828_ (.A1(_05540_),
    .A2(_05543_),
    .B1(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__xnor2_1 _12829_ (.A(_05583_),
    .B(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__and3_1 _12830_ (.A(_05477_),
    .B(_05480_),
    .C(_05485_),
    .X(_05587_));
 sky130_fd_sc_hd__a21o_1 _12831_ (.A1(_05475_),
    .A2(_05486_),
    .B1(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a22oi_2 _12832_ (.A1(_05492_),
    .A2(_05548_),
    .B1(_05553_),
    .B2(_05547_),
    .Y(_05589_));
 sky130_fd_sc_hd__or2_1 _12833_ (.A(_05484_),
    .B(_05474_),
    .X(_05590_));
 sky130_fd_sc_hd__and4_1 _12834_ (.A(_05491_),
    .B(_05477_),
    .C(_05450_),
    .D(_05479_),
    .X(_05591_));
 sky130_fd_sc_hd__and2_1 _12835_ (.A(_05467_),
    .B(_05483_),
    .X(_05592_));
 sky130_fd_sc_hd__buf_2 _12836_ (.A(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__o22a_1 _12837_ (.A1(_05499_),
    .A2(_05493_),
    .B1(_05593_),
    .B2(_05433_),
    .X(_05594_));
 sky130_fd_sc_hd__nor2_1 _12838_ (.A(_05591_),
    .B(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__xnor2_1 _12839_ (.A(_05590_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__xnor2_1 _12840_ (.A(_05589_),
    .B(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__xnor2_1 _12841_ (.A(_05588_),
    .B(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__xnor2_1 _12842_ (.A(_05586_),
    .B(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__xor2_1 _12843_ (.A(_05574_),
    .B(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__xor2_1 _12844_ (.A(_05529_),
    .B(_05531_),
    .X(_05601_));
 sky130_fd_sc_hd__and2b_1 _12845_ (.A_N(_05599_),
    .B(_05574_),
    .X(_05602_));
 sky130_fd_sc_hd__o21ba_1 _12846_ (.A1(_05600_),
    .A2(_05601_),
    .B1_N(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__and2_1 _12847_ (.A(_05583_),
    .B(_05585_),
    .X(_05604_));
 sky130_fd_sc_hd__nor2_1 _12848_ (.A(_05586_),
    .B(_05598_),
    .Y(_05605_));
 sky130_fd_sc_hd__nor2_2 _12849_ (.A(_05355_),
    .B(_05496_),
    .Y(_05606_));
 sky130_fd_sc_hd__nor2_1 _12850_ (.A(_05301_),
    .B(_05551_),
    .Y(_05607_));
 sky130_fd_sc_hd__xnor2_1 _12851_ (.A(_05606_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__buf_2 _12852_ (.A(_05392_),
    .X(_05609_));
 sky130_fd_sc_hd__clkbuf_4 _12853_ (.A(_05546_),
    .X(_05610_));
 sky130_fd_sc_hd__or2_1 _12854_ (.A(_05609_),
    .B(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__xnor2_1 _12855_ (.A(_05608_),
    .B(_05611_),
    .Y(_05612_));
 sky130_fd_sc_hd__o21ai_1 _12856_ (.A1(_05536_),
    .A2(_05582_),
    .B1(_05537_),
    .Y(_05613_));
 sky130_fd_sc_hd__xor2_1 _12857_ (.A(_05612_),
    .B(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__nand2_1 _12858_ (.A(_05609_),
    .B(_05467_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand2_2 _12859_ (.A(_05469_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__a31o_1 _12860_ (.A1(_05494_),
    .A2(_05616_),
    .A3(_05595_),
    .B1(_05591_),
    .X(_05617_));
 sky130_fd_sc_hd__nor2_1 _12861_ (.A(_05609_),
    .B(_05551_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _12862_ (.A(_05618_),
    .B(_05606_),
    .Y(_05619_));
 sky130_fd_sc_hd__or2_1 _12863_ (.A(_05433_),
    .B(_05474_),
    .X(_05620_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(_05491_),
    .B(_05499_),
    .Y(_05621_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(_05616_),
    .A1(_05620_),
    .S(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__a21oi_1 _12866_ (.A1(_05619_),
    .A2(_05580_),
    .B1(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__and3_1 _12867_ (.A(_05619_),
    .B(_05580_),
    .C(_05622_),
    .X(_05624_));
 sky130_fd_sc_hd__or2_1 _12868_ (.A(_05623_),
    .B(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__xnor2_1 _12869_ (.A(_05617_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__xnor2_1 _12870_ (.A(_05614_),
    .B(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21ai_1 _12871_ (.A1(_05604_),
    .A2(_05605_),
    .B1(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__or3_1 _12872_ (.A(_05604_),
    .B(_05605_),
    .C(_05627_),
    .X(_05629_));
 sky130_fd_sc_hd__nand2_1 _12873_ (.A(_05628_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__or2b_1 _12874_ (.A(_05519_),
    .B_N(_05522_),
    .X(_05631_));
 sky130_fd_sc_hd__and2b_1 _12875_ (.A_N(_05589_),
    .B(_05596_),
    .X(_05632_));
 sky130_fd_sc_hd__a21o_1 _12876_ (.A1(_05588_),
    .A2(_05597_),
    .B1(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__or2_1 _12877_ (.A(_05473_),
    .B(_05517_),
    .X(_05634_));
 sky130_fd_sc_hd__nor2_1 _12878_ (.A(_05484_),
    .B(_05471_),
    .Y(_05635_));
 sky130_fd_sc_hd__or3_1 _12879_ (.A(_05513_),
    .B(_05634_),
    .C(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__xor2_1 _12880_ (.A(_05634_),
    .B(_05635_),
    .X(_05637_));
 sky130_fd_sc_hd__o21ai_1 _12881_ (.A1(_05520_),
    .A2(_05521_),
    .B1(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__and2_1 _12882_ (.A(_05636_),
    .B(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__xnor2_1 _12883_ (.A(_05633_),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__nor2_1 _12884_ (.A(_05631_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__and2_1 _12885_ (.A(_05631_),
    .B(_05640_),
    .X(_05642_));
 sky130_fd_sc_hd__nor2_1 _12886_ (.A(_05641_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__xnor2_1 _12887_ (.A(_05630_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__xnor2_1 _12888_ (.A(_05603_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__xnor2_1 _12889_ (.A(_05533_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__xnor2_1 _12890_ (.A(_05506_),
    .B(_05509_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_2 _12891_ (.A(_05477_),
    .B(_05549_),
    .Y(_05648_));
 sky130_fd_sc_hd__or2_1 _12892_ (.A(_05493_),
    .B(_05550_),
    .X(_05649_));
 sky130_fd_sc_hd__xnor2_2 _12893_ (.A(_05649_),
    .B(_05648_),
    .Y(_05650_));
 sky130_fd_sc_hd__nand2_1 _12894_ (.A(_05494_),
    .B(_05576_),
    .Y(_05651_));
 sky130_fd_sc_hd__o32ai_4 _12895_ (.A1(_05493_),
    .A2(_05551_),
    .A3(_05648_),
    .B1(_05650_),
    .B2(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__and2b_1 _12896_ (.A_N(_05647_),
    .B(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__nor2_1 _12897_ (.A(_05505_),
    .B(_05502_),
    .Y(_05654_));
 sky130_fd_sc_hd__nor2_1 _12898_ (.A(_05516_),
    .B(_05474_),
    .Y(_05655_));
 sky130_fd_sc_hd__a21o_1 _12899_ (.A1(_05467_),
    .A2(_05483_),
    .B1(_05505_),
    .X(_05656_));
 sky130_fd_sc_hd__xnor2_1 _12900_ (.A(_05504_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__a22oi_2 _12901_ (.A1(_05508_),
    .A2(_05654_),
    .B1(_05655_),
    .B2(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__xnor2_1 _12902_ (.A(_05652_),
    .B(_05647_),
    .Y(_05659_));
 sky130_fd_sc_hd__and2b_1 _12903_ (.A_N(_05658_),
    .B(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__or3_1 _12904_ (.A(_05526_),
    .B(_05471_),
    .C(_05518_),
    .X(_05661_));
 sky130_fd_sc_hd__xnor2_1 _12905_ (.A(_05525_),
    .B(_05518_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_1 _12906_ (.A(_05661_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__o21a_1 _12907_ (.A1(_05653_),
    .A2(_05660_),
    .B1(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__xnor2_1 _12908_ (.A(_05567_),
    .B(_05568_),
    .Y(_05665_));
 sky130_fd_sc_hd__xor2_1 _12909_ (.A(_05561_),
    .B(_05564_),
    .X(_05666_));
 sky130_fd_sc_hd__nor2_1 _12910_ (.A(_05493_),
    .B(_05536_),
    .Y(_05667_));
 sky130_fd_sc_hd__a2bb2o_1 _12911_ (.A1_N(_05392_),
    .A2_N(_05526_),
    .B1(_05538_),
    .B2(_05465_),
    .X(_05668_));
 sky130_fd_sc_hd__and4b_1 _12912_ (.A_N(_05392_),
    .B(_05465_),
    .C(_05534_),
    .D(_05538_),
    .X(_05669_));
 sky130_fd_sc_hd__a21oi_1 _12913_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__xor2_1 _12914_ (.A(_05666_),
    .B(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__xnor2_1 _12915_ (.A(_05651_),
    .B(_05650_),
    .Y(_05672_));
 sky130_fd_sc_hd__or2b_1 _12916_ (.A(_05670_),
    .B_N(_05666_),
    .X(_05673_));
 sky130_fd_sc_hd__o21a_1 _12917_ (.A1(_05671_),
    .A2(_05672_),
    .B1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__xor2_1 _12918_ (.A(_05665_),
    .B(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__xnor2_1 _12919_ (.A(_05658_),
    .B(_05659_),
    .Y(_05676_));
 sky130_fd_sc_hd__nor2_1 _12920_ (.A(_05665_),
    .B(_05674_),
    .Y(_05677_));
 sky130_fd_sc_hd__a21oi_1 _12921_ (.A1(_05675_),
    .A2(_05676_),
    .B1(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__xnor2_1 _12922_ (.A(_05571_),
    .B(_05572_),
    .Y(_05679_));
 sky130_fd_sc_hd__xnor2_1 _12923_ (.A(_05678_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__nor3_1 _12924_ (.A(_05653_),
    .B(_05660_),
    .C(_05663_),
    .Y(_05681_));
 sky130_fd_sc_hd__o32a_1 _12925_ (.A1(_05680_),
    .A2(_05664_),
    .A3(_05681_),
    .B1(_05679_),
    .B2(_05678_),
    .X(_05682_));
 sky130_fd_sc_hd__xor2_1 _12926_ (.A(_05600_),
    .B(_05601_),
    .X(_05683_));
 sky130_fd_sc_hd__xnor2_1 _12927_ (.A(_05682_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__or2b_1 _12928_ (.A(_05682_),
    .B_N(_05683_),
    .X(_05685_));
 sky130_fd_sc_hd__a21boi_1 _12929_ (.A1(_05664_),
    .A2(_05684_),
    .B1_N(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__xnor2_1 _12930_ (.A(_05646_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__xnor2_1 _12931_ (.A(_05655_),
    .B(_05657_),
    .Y(_05688_));
 sky130_fd_sc_hd__nor2_1 _12932_ (.A(_05450_),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__a21oi_1 _12933_ (.A1(_05467_),
    .A2(_05483_),
    .B1(_05516_),
    .Y(_05690_));
 sky130_fd_sc_hd__or2_1 _12934_ (.A(_05526_),
    .B(_05474_),
    .X(_05691_));
 sky130_fd_sc_hd__xnor2_1 _12935_ (.A(_05654_),
    .B(_05690_),
    .Y(_05692_));
 sky130_fd_sc_hd__o2bb2a_1 _12936_ (.A1_N(_05654_),
    .A2_N(_05690_),
    .B1(_05691_),
    .B2(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__xnor2_1 _12937_ (.A(_05499_),
    .B(_05688_),
    .Y(_05694_));
 sky130_fd_sc_hd__and2b_1 _12938_ (.A_N(_05693_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__inv_2 _12939_ (.A(_05517_),
    .Y(_05696_));
 sky130_fd_sc_hd__clkbuf_4 _12940_ (.A(_05534_),
    .X(_05697_));
 sky130_fd_sc_hd__a2bb2o_1 _12941_ (.A1_N(_05516_),
    .A2_N(_05471_),
    .B1(_05696_),
    .B2(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__and2_1 _12942_ (.A(_05661_),
    .B(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__o21a_1 _12943_ (.A1(_05689_),
    .A2(_05695_),
    .B1(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__xnor2_1 _12944_ (.A(_05671_),
    .B(_05672_),
    .Y(_05701_));
 sky130_fd_sc_hd__and2b_1 _12945_ (.A_N(_05669_),
    .B(_05668_),
    .X(_05702_));
 sky130_fd_sc_hd__xnor2_1 _12946_ (.A(_05667_),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__or4b_1 _12947_ (.A(_05526_),
    .B(_05493_),
    .C(_05535_),
    .D_N(_05465_),
    .X(_05704_));
 sky130_fd_sc_hd__nor2_1 _12948_ (.A(_05433_),
    .B(_05536_),
    .Y(_05705_));
 sky130_fd_sc_hd__a22o_1 _12949_ (.A1(_05465_),
    .A2(_05697_),
    .B1(_05479_),
    .B2(_05538_),
    .X(_05706_));
 sky130_fd_sc_hd__nand3_1 _12950_ (.A(_05704_),
    .B(_05705_),
    .C(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand2_1 _12951_ (.A(_05704_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__xor2_1 _12952_ (.A(_05703_),
    .B(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__mux2_1 _12953_ (.A0(_05473_),
    .A1(_05551_),
    .S(_05610_),
    .X(_05710_));
 sky130_fd_sc_hd__or2b_1 _12954_ (.A(_05703_),
    .B_N(_05708_),
    .X(_05711_));
 sky130_fd_sc_hd__o21ai_2 _12955_ (.A1(_05709_),
    .A2(_05710_),
    .B1(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__xnor2_1 _12956_ (.A(_05701_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__xnor2_1 _12957_ (.A(_05693_),
    .B(_05694_),
    .Y(_05714_));
 sky130_fd_sc_hd__and2b_1 _12958_ (.A_N(_05701_),
    .B(_05712_),
    .X(_05715_));
 sky130_fd_sc_hd__a21oi_1 _12959_ (.A1(_05713_),
    .A2(_05714_),
    .B1(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__xnor2_1 _12960_ (.A(_05675_),
    .B(_05676_),
    .Y(_05717_));
 sky130_fd_sc_hd__xor2_1 _12961_ (.A(_05716_),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nor3_1 _12962_ (.A(_05689_),
    .B(_05695_),
    .C(_05699_),
    .Y(_05719_));
 sky130_fd_sc_hd__nor2_1 _12963_ (.A(_05700_),
    .B(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__nor2_1 _12964_ (.A(_05716_),
    .B(_05717_),
    .Y(_05721_));
 sky130_fd_sc_hd__a21o_1 _12965_ (.A1(_05718_),
    .A2(_05720_),
    .B1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__or2_1 _12966_ (.A(_05664_),
    .B(_05681_),
    .X(_05723_));
 sky130_fd_sc_hd__xor2_1 _12967_ (.A(_05680_),
    .B(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__xor2_1 _12968_ (.A(_05722_),
    .B(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__xnor2_1 _12969_ (.A(_05700_),
    .B(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__xnor2_1 _12970_ (.A(_05691_),
    .B(_05692_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand2_1 _12971_ (.A(_05697_),
    .B(_05480_),
    .Y(_05728_));
 sky130_fd_sc_hd__xor2_1 _12972_ (.A(_05495_),
    .B(_05727_),
    .X(_05729_));
 sky130_fd_sc_hd__or4b_1 _12973_ (.A(_05516_),
    .B(_05728_),
    .C(_05593_),
    .D_N(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__o21a_1 _12974_ (.A1(_05495_),
    .A2(_05727_),
    .B1(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__and2b_1 _12975_ (.A_N(_05731_),
    .B(_05528_),
    .X(_05732_));
 sky130_fd_sc_hd__xor2_1 _12976_ (.A(_05709_),
    .B(_05710_),
    .X(_05733_));
 sky130_fd_sc_hd__a21o_1 _12977_ (.A1(_05704_),
    .A2(_05706_),
    .B1(_05705_),
    .X(_05734_));
 sky130_fd_sc_hd__nor2_1 _12978_ (.A(_05484_),
    .B(_05536_),
    .Y(_05735_));
 sky130_fd_sc_hd__a22o_1 _12979_ (.A1(_05697_),
    .A2(_05479_),
    .B1(_05538_),
    .B2(_05477_),
    .X(_05736_));
 sky130_fd_sc_hd__nor2_1 _12980_ (.A(_05526_),
    .B(_05433_),
    .Y(_05737_));
 sky130_fd_sc_hd__or3b_1 _12981_ (.A(_05493_),
    .B(_05535_),
    .C_N(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__a21bo_1 _12982_ (.A1(_05735_),
    .A2(_05736_),
    .B1_N(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__a21o_1 _12983_ (.A1(_05707_),
    .A2(_05734_),
    .B1(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__nand2_1 _12984_ (.A(_05484_),
    .B(_05473_),
    .Y(_05741_));
 sky130_fd_sc_hd__o211a_1 _12985_ (.A1(_05484_),
    .A2(_05473_),
    .B1(_05505_),
    .C1(_05425_),
    .X(_05742_));
 sky130_fd_sc_hd__a2bb2o_1 _12986_ (.A1_N(_05505_),
    .A2_N(_05610_),
    .B1(_05741_),
    .B2(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__and3_1 _12987_ (.A(_05707_),
    .B(_05734_),
    .C(_05739_),
    .X(_05744_));
 sky130_fd_sc_hd__a21oi_1 _12988_ (.A1(_05740_),
    .A2(_05743_),
    .B1(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__xnor2_1 _12989_ (.A(_05733_),
    .B(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__or3_1 _12990_ (.A(_05516_),
    .B(_05593_),
    .C(_05728_),
    .X(_05747_));
 sky130_fd_sc_hd__xnor2_1 _12991_ (.A(_05729_),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__and2b_1 _12992_ (.A_N(_05745_),
    .B(_05733_),
    .X(_05749_));
 sky130_fd_sc_hd__a21o_1 _12993_ (.A1(_05746_),
    .A2(_05748_),
    .B1(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__xnor2_1 _12994_ (.A(_05713_),
    .B(_05714_),
    .Y(_05751_));
 sky130_fd_sc_hd__xnor2_1 _12995_ (.A(_05750_),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__xnor2_1 _12996_ (.A(_05528_),
    .B(_05731_),
    .Y(_05753_));
 sky130_fd_sc_hd__and2b_1 _12997_ (.A_N(_05751_),
    .B(_05750_),
    .X(_05754_));
 sky130_fd_sc_hd__a21oi_1 _12998_ (.A1(_05752_),
    .A2(_05753_),
    .B1(_05754_),
    .Y(_05755_));
 sky130_fd_sc_hd__xor2_1 _12999_ (.A(_05718_),
    .B(_05720_),
    .X(_05756_));
 sky130_fd_sc_hd__xnor2_1 _13000_ (.A(_05755_),
    .B(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__and2b_1 _13001_ (.A_N(_05755_),
    .B(_05756_),
    .X(_05758_));
 sky130_fd_sc_hd__a21oi_1 _13002_ (.A1(_05732_),
    .A2(_05757_),
    .B1(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__nor2_1 _13003_ (.A(_05726_),
    .B(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__xnor2_1 _13004_ (.A(_05664_),
    .B(_05684_),
    .Y(_05761_));
 sky130_fd_sc_hd__and2_1 _13005_ (.A(_05700_),
    .B(_05725_),
    .X(_05762_));
 sky130_fd_sc_hd__a21oi_1 _13006_ (.A1(_05722_),
    .A2(_05724_),
    .B1(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__xnor2_1 _13007_ (.A(_05761_),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__inv_2 _13008_ (.A(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__nand2_1 _13009_ (.A(_05760_),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__xnor2_1 _13010_ (.A(_05732_),
    .B(_05757_),
    .Y(_05767_));
 sky130_fd_sc_hd__nand2_2 _13011_ (.A(_05467_),
    .B(_05483_),
    .Y(_05768_));
 sky130_fd_sc_hd__a2bb2o_1 _13012_ (.A1_N(_05516_),
    .A2_N(_05503_),
    .B1(_05768_),
    .B2(_05697_),
    .X(_05769_));
 sky130_fd_sc_hd__nand2_1 _13013_ (.A(_05747_),
    .B(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__nor2_1 _13014_ (.A(_05516_),
    .B(_05610_),
    .Y(_05771_));
 sky130_fd_sc_hd__mux2_1 _13015_ (.A0(_05484_),
    .A1(_05489_),
    .S(_05505_),
    .X(_05772_));
 sky130_fd_sc_hd__a22o_1 _13016_ (.A1(_05494_),
    .A2(_05488_),
    .B1(_05771_),
    .B2(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__xnor2_1 _13017_ (.A(_05770_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__and2b_1 _13018_ (.A_N(_05744_),
    .B(_05740_),
    .X(_05775_));
 sky130_fd_sc_hd__xnor2_1 _13019_ (.A(_05775_),
    .B(_05743_),
    .Y(_05776_));
 sky130_fd_sc_hd__nand3_1 _13020_ (.A(_05738_),
    .B(_05735_),
    .C(_05736_),
    .Y(_05777_));
 sky130_fd_sc_hd__a21o_1 _13021_ (.A1(_05738_),
    .A2(_05736_),
    .B1(_05735_),
    .X(_05778_));
 sky130_fd_sc_hd__nor2_1 _13022_ (.A(_05473_),
    .B(_05536_),
    .Y(_05779_));
 sky130_fd_sc_hd__a21o_1 _13023_ (.A1(_05494_),
    .A2(_05538_),
    .B1(_05737_),
    .X(_05780_));
 sky130_fd_sc_hd__and3_1 _13024_ (.A(_05494_),
    .B(_05538_),
    .C(_05737_),
    .X(_05781_));
 sky130_fd_sc_hd__a21o_1 _13025_ (.A1(_05779_),
    .A2(_05780_),
    .B1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__xor2_1 _13026_ (.A(_05771_),
    .B(_05772_),
    .X(_05783_));
 sky130_fd_sc_hd__nand2_1 _13027_ (.A(_05777_),
    .B(_05778_),
    .Y(_05784_));
 sky130_fd_sc_hd__xnor2_1 _13028_ (.A(_05784_),
    .B(_05782_),
    .Y(_05785_));
 sky130_fd_sc_hd__a32o_1 _13029_ (.A1(_05777_),
    .A2(_05778_),
    .A3(_05782_),
    .B1(_05783_),
    .B2(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__xnor2_1 _13030_ (.A(_05776_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__or2b_1 _13031_ (.A(_05776_),
    .B_N(_05786_),
    .X(_05788_));
 sky130_fd_sc_hd__a21bo_1 _13032_ (.A1(_05774_),
    .A2(_05787_),
    .B1_N(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__xor2_1 _13033_ (.A(_05746_),
    .B(_05748_),
    .X(_05790_));
 sky130_fd_sc_hd__and2_1 _13034_ (.A(_05789_),
    .B(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__or2b_1 _13035_ (.A(_05770_),
    .B_N(_05773_),
    .X(_05792_));
 sky130_fd_sc_hd__nor2_1 _13036_ (.A(_05789_),
    .B(_05790_),
    .Y(_05793_));
 sky130_fd_sc_hd__or2_1 _13037_ (.A(_05791_),
    .B(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__nor2_1 _13038_ (.A(_05792_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__xor2_1 _13039_ (.A(_05752_),
    .B(_05753_),
    .X(_05796_));
 sky130_fd_sc_hd__o21ai_1 _13040_ (.A1(_05791_),
    .A2(_05795_),
    .B1(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__or2_1 _13041_ (.A(_05767_),
    .B(_05797_),
    .X(_05798_));
 sky130_fd_sc_hd__xor2_1 _13042_ (.A(_05726_),
    .B(_05759_),
    .X(_05799_));
 sky130_fd_sc_hd__or2b_1 _13043_ (.A(_05798_),
    .B_N(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__xnor2_1 _13044_ (.A(_05798_),
    .B(_05799_),
    .Y(_05801_));
 sky130_fd_sc_hd__xor2_1 _13045_ (.A(_05774_),
    .B(_05787_),
    .X(_05802_));
 sky130_fd_sc_hd__or2b_1 _13046_ (.A(_05781_),
    .B_N(_05780_),
    .X(_05803_));
 sky130_fd_sc_hd__xnor2_1 _13047_ (.A(_05779_),
    .B(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__clkbuf_4 _13048_ (.A(_05535_),
    .X(_05805_));
 sky130_fd_sc_hd__o22a_1 _13049_ (.A1(_05484_),
    .A2(_05526_),
    .B1(_05805_),
    .B2(_05473_),
    .X(_05806_));
 sky130_fd_sc_hd__nand2_1 _13050_ (.A(_05494_),
    .B(_05489_),
    .Y(_05807_));
 sky130_fd_sc_hd__o21ai_1 _13051_ (.A1(_05558_),
    .A2(_05806_),
    .B1(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__nand2_1 _13052_ (.A(_05804_),
    .B(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__nor2_1 _13053_ (.A(_05516_),
    .B(_05496_),
    .Y(_05810_));
 sky130_fd_sc_hd__xnor2_1 _13054_ (.A(_05488_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__or3_1 _13055_ (.A(_05527_),
    .B(_05610_),
    .C(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__o21ai_1 _13056_ (.A1(_05527_),
    .A2(_05610_),
    .B1(_05811_),
    .Y(_05813_));
 sky130_fd_sc_hd__and2_1 _13057_ (.A(_05812_),
    .B(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__or2_1 _13058_ (.A(_05804_),
    .B(_05808_),
    .X(_05815_));
 sky130_fd_sc_hd__and2_1 _13059_ (.A(_05809_),
    .B(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__nand2_1 _13060_ (.A(_05814_),
    .B(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__xnor2_1 _13061_ (.A(_05783_),
    .B(_05785_),
    .Y(_05818_));
 sky130_fd_sc_hd__a21oi_1 _13062_ (.A1(_05809_),
    .A2(_05817_),
    .B1(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__a21bo_1 _13063_ (.A1(_05488_),
    .A2(_05810_),
    .B1_N(_05812_),
    .X(_05820_));
 sky130_fd_sc_hd__xor2_1 _13064_ (.A(_05728_),
    .B(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__and3_1 _13065_ (.A(_05818_),
    .B(_05809_),
    .C(_05817_),
    .X(_05822_));
 sky130_fd_sc_hd__nor3_1 _13066_ (.A(_05819_),
    .B(_05821_),
    .C(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__or2_1 _13067_ (.A(_05819_),
    .B(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__and2_1 _13068_ (.A(_05802_),
    .B(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__and3_1 _13069_ (.A(_05697_),
    .B(_05480_),
    .C(_05820_),
    .X(_05826_));
 sky130_fd_sc_hd__inv_2 _13070_ (.A(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__xnor2_1 _13071_ (.A(_05802_),
    .B(_05824_),
    .Y(_05828_));
 sky130_fd_sc_hd__nor2_1 _13072_ (.A(_05827_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__and2_1 _13073_ (.A(_05792_),
    .B(_05794_),
    .X(_05830_));
 sky130_fd_sc_hd__nor2_1 _13074_ (.A(_05795_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__o21ai_1 _13075_ (.A1(_05825_),
    .A2(_05829_),
    .B1(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__or3_1 _13076_ (.A(_05796_),
    .B(_05791_),
    .C(_05795_),
    .X(_05833_));
 sky130_fd_sc_hd__nand2_1 _13077_ (.A(_05797_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__nor3_2 _13078_ (.A(_05767_),
    .B(_05832_),
    .C(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__xor2_2 _13079_ (.A(_05801_),
    .B(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__nand2_1 _13080_ (.A(_05767_),
    .B(_05797_),
    .Y(_05837_));
 sky130_fd_sc_hd__a21oi_1 _13081_ (.A1(_05558_),
    .A2(_05806_),
    .B1(_05808_),
    .Y(_05838_));
 sky130_fd_sc_hd__and2_1 _13082_ (.A(_05489_),
    .B(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__a2bb2o_1 _13083_ (.A1_N(_05516_),
    .A2_N(_05551_),
    .B1(_05549_),
    .B2(_05697_),
    .X(_05840_));
 sky130_fd_sc_hd__o2111a_1 _13084_ (.A1(_05489_),
    .A2(_05838_),
    .B1(_05840_),
    .C1(_05807_),
    .D1(_05817_),
    .X(_05841_));
 sky130_fd_sc_hd__o21ai_1 _13085_ (.A1(_05814_),
    .A2(_05816_),
    .B1(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__nor2_1 _13086_ (.A(_05823_),
    .B(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__o2bb2a_1 _13087_ (.A1_N(_05827_),
    .A2_N(_05828_),
    .B1(_05839_),
    .B2(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__or3_1 _13088_ (.A(_05831_),
    .B(_05825_),
    .C(_05829_),
    .X(_05845_));
 sky130_fd_sc_hd__and3b_1 _13089_ (.A_N(_05834_),
    .B(_05845_),
    .C(_05832_),
    .X(_05846_));
 sky130_fd_sc_hd__and3_1 _13090_ (.A(_05837_),
    .B(_05844_),
    .C(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__and2_1 _13091_ (.A(_05801_),
    .B(_05835_),
    .X(_05848_));
 sky130_fd_sc_hd__a21o_1 _13092_ (.A1(_05836_),
    .A2(_05847_),
    .B1(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__and2b_1 _13093_ (.A_N(_05760_),
    .B(_05800_),
    .X(_05850_));
 sky130_fd_sc_hd__xnor2_1 _13094_ (.A(_05765_),
    .B(_05850_),
    .Y(_05851_));
 sky130_fd_sc_hd__a2bb2o_1 _13095_ (.A1_N(_05764_),
    .A2_N(_05800_),
    .B1(_05849_),
    .B2(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__nor2_1 _13096_ (.A(_05761_),
    .B(_05763_),
    .Y(_05853_));
 sky130_fd_sc_hd__a21o_1 _13097_ (.A1(_05760_),
    .A2(_05765_),
    .B1(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__xnor2_1 _13098_ (.A(_05687_),
    .B(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__a2bb2o_1 _13099_ (.A1_N(_05687_),
    .A2_N(_05766_),
    .B1(_05852_),
    .B2(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__a21o_1 _13100_ (.A1(_05633_),
    .A2(_05639_),
    .B1(_05641_),
    .X(_05857_));
 sky130_fd_sc_hd__or2b_1 _13101_ (.A(_05630_),
    .B_N(_05643_),
    .X(_05858_));
 sky130_fd_sc_hd__or2b_1 _13102_ (.A(_05612_),
    .B_N(_05613_),
    .X(_05859_));
 sky130_fd_sc_hd__or2b_1 _13103_ (.A(_05614_),
    .B_N(_05626_),
    .X(_05860_));
 sky130_fd_sc_hd__nor2_1 _13104_ (.A(_05301_),
    .B(_05610_),
    .Y(_05861_));
 sky130_fd_sc_hd__clkbuf_4 _13105_ (.A(_05496_),
    .X(_05862_));
 sky130_fd_sc_hd__o22a_1 _13106_ (.A1(_05301_),
    .A2(_05862_),
    .B1(_05610_),
    .B2(_05355_),
    .X(_05863_));
 sky130_fd_sc_hd__a21o_1 _13107_ (.A1(_05606_),
    .A2(_05861_),
    .B1(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__o2bb2ai_1 _13108_ (.A1_N(_05606_),
    .A2_N(_05607_),
    .B1(_05608_),
    .B2(_05611_),
    .Y(_05865_));
 sky130_fd_sc_hd__o22a_1 _13109_ (.A1(_05479_),
    .A2(_05474_),
    .B1(_05480_),
    .B2(_05609_),
    .X(_05866_));
 sky130_fd_sc_hd__xnor2_1 _13110_ (.A(_05865_),
    .B(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__a21oi_1 _13111_ (.A1(_05609_),
    .A2(_05499_),
    .B1(_05467_),
    .Y(_05868_));
 sky130_fd_sc_hd__xor2_1 _13112_ (.A(_05867_),
    .B(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__or2_1 _13113_ (.A(_05864_),
    .B(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__nand2_1 _13114_ (.A(_05864_),
    .B(_05869_),
    .Y(_05871_));
 sky130_fd_sc_hd__nand2_1 _13115_ (.A(_05870_),
    .B(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__a21o_1 _13116_ (.A1(_05859_),
    .A2(_05860_),
    .B1(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__nand3_1 _13117_ (.A(_05859_),
    .B(_05860_),
    .C(_05872_),
    .Y(_05874_));
 sky130_fd_sc_hd__and2_1 _13118_ (.A(_05873_),
    .B(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__and2b_1 _13119_ (.A_N(_05625_),
    .B(_05617_),
    .X(_05876_));
 sky130_fd_sc_hd__or2_1 _13120_ (.A(_05623_),
    .B(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__or2_1 _13121_ (.A(_05484_),
    .B(_05517_),
    .X(_05878_));
 sky130_fd_sc_hd__or2_1 _13122_ (.A(_05433_),
    .B(_05471_),
    .X(_05879_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13123_ (.A(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__xnor2_1 _13124_ (.A(_05878_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__or3_1 _13125_ (.A(_05521_),
    .B(_05878_),
    .C(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__o21ai_1 _13126_ (.A1(_05521_),
    .A2(_05878_),
    .B1(_05881_),
    .Y(_05883_));
 sky130_fd_sc_hd__and2_1 _13127_ (.A(_05882_),
    .B(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__xnor2_1 _13128_ (.A(_05877_),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__xor2_1 _13129_ (.A(_05636_),
    .B(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__xnor2_1 _13130_ (.A(_05875_),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__a21o_1 _13131_ (.A1(_05628_),
    .A2(_05858_),
    .B1(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__nand3_1 _13132_ (.A(_05628_),
    .B(_05858_),
    .C(_05887_),
    .Y(_05889_));
 sky130_fd_sc_hd__and2_1 _13133_ (.A(_05888_),
    .B(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__xnor2_1 _13134_ (.A(_05857_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__or2b_1 _13135_ (.A(_05603_),
    .B_N(_05644_),
    .X(_05892_));
 sky130_fd_sc_hd__a21boi_1 _13136_ (.A1(_05533_),
    .A2(_05645_),
    .B1_N(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__xnor2_1 _13137_ (.A(_05891_),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__nor2_1 _13138_ (.A(_05646_),
    .B(_05686_),
    .Y(_05895_));
 sky130_fd_sc_hd__inv_2 _13139_ (.A(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__or3_1 _13140_ (.A(_05687_),
    .B(_05761_),
    .C(_05763_),
    .X(_05897_));
 sky130_fd_sc_hd__and2_1 _13141_ (.A(_05896_),
    .B(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__xor2_1 _13142_ (.A(_05894_),
    .B(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__xnor2_1 _13143_ (.A(_05856_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__xor2_2 _13144_ (.A(_05852_),
    .B(_05855_),
    .X(_05901_));
 sky130_fd_sc_hd__xnor2_2 _13145_ (.A(_05836_),
    .B(_05847_),
    .Y(_05902_));
 sky130_fd_sc_hd__xor2_2 _13146_ (.A(_05849_),
    .B(_05851_),
    .X(_05903_));
 sky130_fd_sc_hd__and2b_1 _13147_ (.A_N(_05902_),
    .B(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__nor2_1 _13148_ (.A(_05901_),
    .B(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__nand2_1 _13149_ (.A(_05900_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__a2bb2o_1 _13150_ (.A1_N(_05894_),
    .A2_N(_05897_),
    .B1(_05899_),
    .B2(_05856_),
    .X(_05907_));
 sky130_fd_sc_hd__nand2_1 _13151_ (.A(_05857_),
    .B(_05890_),
    .Y(_05908_));
 sky130_fd_sc_hd__nor2_1 _13152_ (.A(_05636_),
    .B(_05885_),
    .Y(_05909_));
 sky130_fd_sc_hd__a21oi_1 _13153_ (.A1(_05877_),
    .A2(_05884_),
    .B1(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__nand2_1 _13154_ (.A(_05875_),
    .B(_05886_),
    .Y(_05911_));
 sky130_fd_sc_hd__nand2_1 _13155_ (.A(_05606_),
    .B(_05861_),
    .Y(_05912_));
 sky130_fd_sc_hd__nand2_1 _13156_ (.A(_05491_),
    .B(_05616_),
    .Y(_05913_));
 sky130_fd_sc_hd__nor2_1 _13157_ (.A(_05355_),
    .B(_05503_),
    .Y(_05914_));
 sky130_fd_sc_hd__nor2_1 _13158_ (.A(_05609_),
    .B(_05593_),
    .Y(_05915_));
 sky130_fd_sc_hd__xnor2_1 _13159_ (.A(_05914_),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__xnor2_1 _13160_ (.A(_05913_),
    .B(_05916_),
    .Y(_05917_));
 sky130_fd_sc_hd__xnor2_1 _13161_ (.A(_05912_),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__xor2_1 _13162_ (.A(_05469_),
    .B(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__xnor2_1 _13163_ (.A(_05861_),
    .B(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__or2_1 _13164_ (.A(_05870_),
    .B(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__nand2_1 _13165_ (.A(_05870_),
    .B(_05920_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand2_1 _13166_ (.A(_05921_),
    .B(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__or2b_1 _13167_ (.A(_05867_),
    .B_N(_05868_),
    .X(_05924_));
 sky130_fd_sc_hd__a21bo_1 _13168_ (.A1(_05865_),
    .A2(_05866_),
    .B1_N(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__or2_1 _13169_ (.A(_05433_),
    .B(_05517_),
    .X(_05926_));
 sky130_fd_sc_hd__or4_2 _13170_ (.A(_05484_),
    .B(_05479_),
    .C(_05472_),
    .D(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__or2_1 _13171_ (.A(_05493_),
    .B(_05517_),
    .X(_05928_));
 sky130_fd_sc_hd__nor2_1 _13172_ (.A(_05880_),
    .B(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__o21a_1 _13173_ (.A1(_05493_),
    .A2(_05471_),
    .B1(_05926_),
    .X(_05930_));
 sky130_fd_sc_hd__o22ai_1 _13174_ (.A1(_05878_),
    .A2(_05880_),
    .B1(_05929_),
    .B2(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__and2_1 _13175_ (.A(_05927_),
    .B(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__xor2_1 _13176_ (.A(_05925_),
    .B(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__xnor2_1 _13177_ (.A(_05882_),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__xor2_1 _13178_ (.A(_05923_),
    .B(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__a21o_1 _13179_ (.A1(_05873_),
    .A2(_05911_),
    .B1(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__nand3_1 _13180_ (.A(_05873_),
    .B(_05911_),
    .C(_05935_),
    .Y(_05937_));
 sky130_fd_sc_hd__and2_1 _13181_ (.A(_05936_),
    .B(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__or2b_1 _13182_ (.A(_05910_),
    .B_N(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__or2b_1 _13183_ (.A(_05938_),
    .B_N(_05910_),
    .X(_05940_));
 sky130_fd_sc_hd__nand2_1 _13184_ (.A(_05939_),
    .B(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__a21oi_2 _13185_ (.A1(_05888_),
    .A2(_05908_),
    .B1(_05941_),
    .Y(_05942_));
 sky130_fd_sc_hd__and3_1 _13186_ (.A(_05888_),
    .B(_05908_),
    .C(_05941_),
    .X(_05943_));
 sky130_fd_sc_hd__nor2_1 _13187_ (.A(_05942_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__nor2_1 _13188_ (.A(_05891_),
    .B(_05893_),
    .Y(_05945_));
 sky130_fd_sc_hd__nor2_1 _13189_ (.A(_05896_),
    .B(_05894_),
    .Y(_05946_));
 sky130_fd_sc_hd__nor2_1 _13190_ (.A(_05945_),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__xnor2_1 _13191_ (.A(_05944_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__xor2_1 _13192_ (.A(_05907_),
    .B(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__or2_2 _13193_ (.A(_05906_),
    .B(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__or2b_1 _13194_ (.A(_05923_),
    .B_N(_05934_),
    .X(_05951_));
 sky130_fd_sc_hd__nand2_1 _13195_ (.A(_05861_),
    .B(_05919_),
    .Y(_05952_));
 sky130_fd_sc_hd__and2_1 _13196_ (.A(_05768_),
    .B(_05914_),
    .X(_05953_));
 sky130_fd_sc_hd__nor2_1 _13197_ (.A(_05355_),
    .B(_05593_),
    .Y(_05954_));
 sky130_fd_sc_hd__nor2_1 _13198_ (.A(_05480_),
    .B(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__or2_1 _13199_ (.A(_05953_),
    .B(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__nor2_1 _13200_ (.A(_05952_),
    .B(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__and2_1 _13201_ (.A(_05952_),
    .B(_05956_),
    .X(_05958_));
 sky130_fd_sc_hd__or2_1 _13202_ (.A(_05957_),
    .B(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__or2_1 _13203_ (.A(_05469_),
    .B(_05918_),
    .X(_05960_));
 sky130_fd_sc_hd__o21ai_1 _13204_ (.A1(_05912_),
    .A2(_05917_),
    .B1(_05960_),
    .Y(_05961_));
 sky130_fd_sc_hd__inv_2 _13205_ (.A(_05471_),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_1 _13206_ (.A(_05491_),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__nor2_1 _13207_ (.A(_05928_),
    .B(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__or3_1 _13208_ (.A(_05880_),
    .B(_05928_),
    .C(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__and2_1 _13209_ (.A(_05928_),
    .B(_05963_),
    .X(_05966_));
 sky130_fd_sc_hd__o22ai_1 _13210_ (.A1(_05880_),
    .A2(_05928_),
    .B1(_05964_),
    .B2(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__and2_1 _13211_ (.A(_05965_),
    .B(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__xnor2_1 _13212_ (.A(_05961_),
    .B(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__xnor2_1 _13213_ (.A(_05927_),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__xnor2_1 _13214_ (.A(_05959_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__a21oi_1 _13215_ (.A1(_05921_),
    .A2(_05951_),
    .B1(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__and3_1 _13216_ (.A(_05921_),
    .B(_05951_),
    .C(_05971_),
    .X(_05973_));
 sky130_fd_sc_hd__nor2_1 _13217_ (.A(_05972_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__and2b_1 _13218_ (.A_N(_05882_),
    .B(_05933_),
    .X(_05975_));
 sky130_fd_sc_hd__a21oi_2 _13219_ (.A1(_05925_),
    .A2(_05932_),
    .B1(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__xor2_2 _13220_ (.A(_05974_),
    .B(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__a21oi_4 _13221_ (.A1(_05936_),
    .A2(_05939_),
    .B1(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__and3_1 _13222_ (.A(_05936_),
    .B(_05939_),
    .C(_05977_),
    .X(_05979_));
 sky130_fd_sc_hd__nor2_1 _13223_ (.A(_05978_),
    .B(_05979_),
    .Y(_05980_));
 sky130_fd_sc_hd__xor2_1 _13224_ (.A(_05942_),
    .B(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__and3_1 _13225_ (.A(_05945_),
    .B(_05944_),
    .C(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__a21oi_1 _13226_ (.A1(_05945_),
    .A2(_05944_),
    .B1(_05981_),
    .Y(_05983_));
 sky130_fd_sc_hd__nor2_2 _13227_ (.A(_05982_),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__a22o_2 _13228_ (.A1(_05944_),
    .A2(_05946_),
    .B1(_05948_),
    .B2(_05907_),
    .X(_05985_));
 sky130_fd_sc_hd__xor2_4 _13229_ (.A(_05984_),
    .B(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__xnor2_4 _13230_ (.A(_05950_),
    .B(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__clkbuf_4 _13231_ (.A(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__or2_1 _13232_ (.A(_05472_),
    .B(_05988_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_4 _13233_ (.A(_05517_),
    .X(_05990_));
 sky130_fd_sc_hd__xnor2_1 _13234_ (.A(_05906_),
    .B(_05949_),
    .Y(_05991_));
 sky130_fd_sc_hd__clkbuf_4 _13235_ (.A(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__nor2_1 _13236_ (.A(_05990_),
    .B(_05992_),
    .Y(_05993_));
 sky130_fd_sc_hd__xnor2_1 _13237_ (.A(_05900_),
    .B(_05905_),
    .Y(_05994_));
 sky130_fd_sc_hd__clkbuf_4 _13238_ (.A(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__nor2_1 _13239_ (.A(_05472_),
    .B(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__and3_1 _13240_ (.A(_05989_),
    .B(_05993_),
    .C(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__xnor2_1 _13241_ (.A(_05989_),
    .B(_05993_),
    .Y(_05998_));
 sky130_fd_sc_hd__a21oi_1 _13242_ (.A1(_05993_),
    .A2(_05996_),
    .B1(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__or2_1 _13243_ (.A(_05997_),
    .B(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_4 _13244_ (.A(_05593_),
    .X(_06001_));
 sky130_fd_sc_hd__nor2_4 _13245_ (.A(_05950_),
    .B(_05986_),
    .Y(_06002_));
 sky130_fd_sc_hd__a21o_1 _13246_ (.A1(_05984_),
    .A2(_05985_),
    .B1(_05982_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2_2 _13247_ (.A(_05942_),
    .B(_05980_),
    .Y(_06004_));
 sky130_fd_sc_hd__and2b_1 _13248_ (.A_N(_05976_),
    .B(_05974_),
    .X(_06005_));
 sky130_fd_sc_hd__nor2_1 _13249_ (.A(_05959_),
    .B(_05970_),
    .Y(_06006_));
 sky130_fd_sc_hd__nor2_1 _13250_ (.A(_05469_),
    .B(_05956_),
    .Y(_06007_));
 sky130_fd_sc_hd__clkbuf_4 _13251_ (.A(_05474_),
    .X(_06008_));
 sky130_fd_sc_hd__o22a_1 _13252_ (.A1(_05355_),
    .A2(_06008_),
    .B1(_05593_),
    .B2(_05301_),
    .X(_06009_));
 sky130_fd_sc_hd__a31oi_1 _13253_ (.A1(_05235_),
    .A2(_05616_),
    .A3(_05954_),
    .B1(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__o21a_1 _13254_ (.A1(_05953_),
    .A2(_06007_),
    .B1(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__nor3_1 _13255_ (.A(_05953_),
    .B(_06007_),
    .C(_06010_),
    .Y(_06012_));
 sky130_fd_sc_hd__nor2_1 _13256_ (.A(_06011_),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__o2bb2a_1 _13257_ (.A1_N(_05491_),
    .A2_N(_05696_),
    .B1(_05472_),
    .B2(_05609_),
    .X(_06014_));
 sky130_fd_sc_hd__or4b_1 _13258_ (.A(_05609_),
    .B(_05990_),
    .C(_05472_),
    .D_N(_05491_),
    .X(_06015_));
 sky130_fd_sc_hd__inv_2 _13259_ (.A(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__nor2_1 _13260_ (.A(_05469_),
    .B(_06007_),
    .Y(_06017_));
 sky130_fd_sc_hd__or4_1 _13261_ (.A(_05964_),
    .B(_06014_),
    .C(_06016_),
    .D(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__xor2_1 _13262_ (.A(_05965_),
    .B(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__nand2_1 _13263_ (.A(_06013_),
    .B(_06019_),
    .Y(_06020_));
 sky130_fd_sc_hd__or2_1 _13264_ (.A(_06013_),
    .B(_06019_),
    .X(_06021_));
 sky130_fd_sc_hd__and2_1 _13265_ (.A(_06020_),
    .B(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__o21a_1 _13266_ (.A1(_05957_),
    .A2(_06006_),
    .B1(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__nor3_1 _13267_ (.A(_05957_),
    .B(_06006_),
    .C(_06022_),
    .Y(_06024_));
 sky130_fd_sc_hd__nor2_1 _13268_ (.A(_06023_),
    .B(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__nor2_1 _13269_ (.A(_05927_),
    .B(_05969_),
    .Y(_06026_));
 sky130_fd_sc_hd__a21oi_1 _13270_ (.A1(_05961_),
    .A2(_05968_),
    .B1(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__xnor2_1 _13271_ (.A(_06025_),
    .B(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__o21ai_1 _13272_ (.A1(_05972_),
    .A2(_06005_),
    .B1(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__or3_1 _13273_ (.A(_05972_),
    .B(_06005_),
    .C(_06028_),
    .X(_06030_));
 sky130_fd_sc_hd__and2_1 _13274_ (.A(_06029_),
    .B(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__xor2_4 _13275_ (.A(_05978_),
    .B(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__xnor2_4 _13276_ (.A(_06004_),
    .B(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__xnor2_4 _13277_ (.A(_06003_),
    .B(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__xnor2_4 _13278_ (.A(_06002_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__o22a_1 _13279_ (.A1(_06001_),
    .A2(_05987_),
    .B1(_06035_),
    .B2(_05503_),
    .X(_06036_));
 sky130_fd_sc_hd__nor2_1 _13280_ (.A(_06008_),
    .B(_05992_),
    .Y(_06037_));
 sky130_fd_sc_hd__and2b_1 _13281_ (.A_N(_06036_),
    .B(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__and2_1 _13282_ (.A(_05984_),
    .B(_05985_),
    .X(_06039_));
 sky130_fd_sc_hd__and2b_1 _13283_ (.A_N(_06027_),
    .B(_06025_),
    .X(_06040_));
 sky130_fd_sc_hd__or2_1 _13284_ (.A(_05609_),
    .B(_06016_),
    .X(_06041_));
 sky130_fd_sc_hd__xnor2_1 _13285_ (.A(_06011_),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__o21ba_1 _13286_ (.A1(_05965_),
    .A2(_06018_),
    .B1_N(_06017_),
    .X(_06043_));
 sky130_fd_sc_hd__o21a_1 _13287_ (.A1(_05964_),
    .A2(_06042_),
    .B1(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__or3_1 _13288_ (.A(_05301_),
    .B(_06008_),
    .C(_05954_),
    .X(_06045_));
 sky130_fd_sc_hd__xor2_1 _13289_ (.A(_06020_),
    .B(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__xnor2_1 _13290_ (.A(_06044_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__or3_1 _13291_ (.A(_06023_),
    .B(_06040_),
    .C(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__a21boi_1 _13292_ (.A1(_05914_),
    .A2(_05915_),
    .B1_N(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__nor2_1 _13293_ (.A(_06029_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__a221o_1 _13294_ (.A1(_05978_),
    .A2(_06031_),
    .B1(_06049_),
    .B2(_06029_),
    .C1(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__inv_2 _13295_ (.A(_05982_),
    .Y(_06052_));
 sky130_fd_sc_hd__a21boi_1 _13296_ (.A1(_06004_),
    .A2(_06052_),
    .B1_N(_06032_),
    .Y(_06053_));
 sky130_fd_sc_hd__a211oi_4 _13297_ (.A1(_06039_),
    .A2(_06033_),
    .B1(_06051_),
    .C1(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__a21oi_4 _13298_ (.A1(_06002_),
    .A2(_06034_),
    .B1(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__buf_2 _13299_ (.A(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__and3_1 _13300_ (.A(_05549_),
    .B(_05576_),
    .C(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13301_ (.A(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__or2_1 _13302_ (.A(_06008_),
    .B(_05988_),
    .X(_06059_));
 sky130_fd_sc_hd__nand2_2 _13303_ (.A(_05480_),
    .B(_06056_),
    .Y(_06060_));
 sky130_fd_sc_hd__clkbuf_4 _13304_ (.A(_06035_),
    .X(_06061_));
 sky130_fd_sc_hd__nor2_1 _13305_ (.A(_06001_),
    .B(_06061_),
    .Y(_06062_));
 sky130_fd_sc_hd__xnor2_1 _13306_ (.A(_06060_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__xnor2_1 _13307_ (.A(_06059_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__xor2_1 _13308_ (.A(_06058_),
    .B(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__and2_1 _13309_ (.A(_06058_),
    .B(_06064_),
    .X(_06066_));
 sky130_fd_sc_hd__a21oi_1 _13310_ (.A1(_06038_),
    .A2(_06065_),
    .B1(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__nor2_1 _13311_ (.A(_05990_),
    .B(_05995_),
    .Y(_06068_));
 sky130_fd_sc_hd__and2_1 _13312_ (.A(_05901_),
    .B(_05904_),
    .X(_06069_));
 sky130_fd_sc_hd__or2_1 _13313_ (.A(_05905_),
    .B(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__clkbuf_4 _13314_ (.A(_06070_),
    .X(_06071_));
 sky130_fd_sc_hd__nor2_1 _13315_ (.A(_05472_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__nand2_1 _13316_ (.A(_06068_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__or2_1 _13317_ (.A(_05472_),
    .B(_05992_),
    .X(_06074_));
 sky130_fd_sc_hd__xor2_1 _13318_ (.A(_06074_),
    .B(_06068_),
    .X(_06075_));
 sky130_fd_sc_hd__nor2_1 _13319_ (.A(_06073_),
    .B(_06075_),
    .Y(_06076_));
 sky130_fd_sc_hd__xor2_1 _13320_ (.A(_06000_),
    .B(_06067_),
    .X(_06077_));
 sky130_fd_sc_hd__nand2_1 _13321_ (.A(_06076_),
    .B(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__o21ai_1 _13322_ (.A1(_06000_),
    .A2(_06067_),
    .B1(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__or2_1 _13323_ (.A(_05990_),
    .B(_06061_),
    .X(_06080_));
 sky130_fd_sc_hd__and2_1 _13324_ (.A(_05962_),
    .B(_06056_),
    .X(_06081_));
 sky130_fd_sc_hd__nor2_1 _13325_ (.A(_05989_),
    .B(_06080_),
    .Y(_06082_));
 sky130_fd_sc_hd__o22a_1 _13326_ (.A1(_05990_),
    .A2(_05988_),
    .B1(_06061_),
    .B2(_05472_),
    .X(_06083_));
 sky130_fd_sc_hd__o32a_1 _13327_ (.A1(_05990_),
    .A2(_06074_),
    .A3(_05988_),
    .B1(_06082_),
    .B2(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__a21o_1 _13328_ (.A1(_06080_),
    .A2(_06081_),
    .B1(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__and2_1 _13329_ (.A(_05768_),
    .B(_06055_),
    .X(_06086_));
 sky130_fd_sc_hd__xnor2_2 _13330_ (.A(_06060_),
    .B(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__nor2_1 _13331_ (.A(_06008_),
    .B(_06061_),
    .Y(_06088_));
 sky130_fd_sc_hd__xor2_1 _13332_ (.A(_06087_),
    .B(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__xnor2_1 _13333_ (.A(_06058_),
    .B(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__or2b_1 _13334_ (.A(_06059_),
    .B_N(_06063_),
    .X(_06091_));
 sky130_fd_sc_hd__o31a_1 _13335_ (.A1(_06001_),
    .A2(_06061_),
    .A3(_06060_),
    .B1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__nand2_1 _13336_ (.A(_06058_),
    .B(_06089_),
    .Y(_06093_));
 sky130_fd_sc_hd__o21a_1 _13337_ (.A1(_06090_),
    .A2(_06092_),
    .B1(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__xor2_1 _13338_ (.A(_06085_),
    .B(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__xor2_1 _13339_ (.A(_05997_),
    .B(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__buf_4 _13340_ (.A(_05301_),
    .X(_06097_));
 sky130_fd_sc_hd__nor2_2 _13341_ (.A(_06097_),
    .B(_06055_),
    .Y(_06098_));
 sky130_fd_sc_hd__and2_1 _13342_ (.A(_05576_),
    .B(_06055_),
    .X(_06099_));
 sky130_fd_sc_hd__a211o_1 _13343_ (.A1(_05549_),
    .A2(_06098_),
    .B1(_06099_),
    .C1(_06097_),
    .X(_06100_));
 sky130_fd_sc_hd__xor2_1 _13344_ (.A(_06090_),
    .B(_06092_),
    .X(_06101_));
 sky130_fd_sc_hd__nand2_1 _13345_ (.A(_06100_),
    .B(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__clkbuf_4 _13346_ (.A(_05610_),
    .X(_06103_));
 sky130_fd_sc_hd__or2_1 _13347_ (.A(_06001_),
    .B(_06060_),
    .X(_06104_));
 sky130_fd_sc_hd__nand2_1 _13348_ (.A(_06087_),
    .B(_06088_),
    .Y(_06105_));
 sky130_fd_sc_hd__and2_1 _13349_ (.A(_05616_),
    .B(_06056_),
    .X(_06106_));
 sky130_fd_sc_hd__nand2_1 _13350_ (.A(_06087_),
    .B(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__or2_1 _13351_ (.A(_06087_),
    .B(_06106_),
    .X(_06108_));
 sky130_fd_sc_hd__nand2_1 _13352_ (.A(_06107_),
    .B(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__and3b_1 _13353_ (.A_N(_05609_),
    .B(_06011_),
    .C(_06015_),
    .X(_06110_));
 sky130_fd_sc_hd__a31o_1 _13354_ (.A1(_06104_),
    .A2(_06105_),
    .A3(_06109_),
    .B1(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__o21a_1 _13355_ (.A1(_06103_),
    .A2(_06056_),
    .B1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__xor2_1 _13356_ (.A(_06102_),
    .B(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__nand2_1 _13357_ (.A(_06096_),
    .B(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__or2_1 _13358_ (.A(_06096_),
    .B(_06113_),
    .X(_06115_));
 sky130_fd_sc_hd__nand2_1 _13359_ (.A(_06114_),
    .B(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__or2_1 _13360_ (.A(_06076_),
    .B(_06077_),
    .X(_06117_));
 sky130_fd_sc_hd__and2_1 _13361_ (.A(_06078_),
    .B(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__xnor2_1 _13362_ (.A(_06100_),
    .B(_06101_),
    .Y(_06119_));
 sky130_fd_sc_hd__xor2_1 _13363_ (.A(_06038_),
    .B(_06065_),
    .X(_06120_));
 sky130_fd_sc_hd__buf_2 _13364_ (.A(_05551_),
    .X(_06121_));
 sky130_fd_sc_hd__buf_2 _13365_ (.A(_05536_),
    .X(_06122_));
 sky130_fd_sc_hd__a211o_1 _13366_ (.A1(_06002_),
    .A2(_06034_),
    .B1(_06054_),
    .C1(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__or2_1 _13367_ (.A(_06121_),
    .B(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__and2_1 _13368_ (.A(_05549_),
    .B(_06055_),
    .X(_06125_));
 sky130_fd_sc_hd__xnor2_1 _13369_ (.A(_06125_),
    .B(_06099_),
    .Y(_06126_));
 sky130_fd_sc_hd__o31a_1 _13370_ (.A1(_06097_),
    .A2(_06121_),
    .A3(_06056_),
    .B1(_06126_),
    .X(_06127_));
 sky130_fd_sc_hd__a211o_1 _13371_ (.A1(_06002_),
    .A2(_06034_),
    .B1(_06054_),
    .C1(_06121_),
    .X(_06128_));
 sky130_fd_sc_hd__nand2_1 _13372_ (.A(_06122_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__a21oi_1 _13373_ (.A1(_06123_),
    .A2(_06129_),
    .B1(_06097_),
    .Y(_06130_));
 sky130_fd_sc_hd__o21a_1 _13374_ (.A1(_06126_),
    .A2(_06130_),
    .B1(_06124_),
    .X(_06131_));
 sky130_fd_sc_hd__nor2_1 _13375_ (.A(_06127_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__a21oi_1 _13376_ (.A1(_06124_),
    .A2(_06127_),
    .B1(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__a21oi_1 _13377_ (.A1(_06120_),
    .A2(_06133_),
    .B1(_06132_),
    .Y(_06134_));
 sky130_fd_sc_hd__nor2_1 _13378_ (.A(_06119_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__and2_1 _13379_ (.A(_06119_),
    .B(_06134_),
    .X(_06136_));
 sky130_fd_sc_hd__nor2_1 _13380_ (.A(_06135_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__a21oi_1 _13381_ (.A1(_06118_),
    .A2(_06137_),
    .B1(_06135_),
    .Y(_06138_));
 sky130_fd_sc_hd__xor2_1 _13382_ (.A(_06116_),
    .B(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__xnor2_1 _13383_ (.A(_06079_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__and2_1 _13384_ (.A(_06073_),
    .B(_06075_),
    .X(_06141_));
 sky130_fd_sc_hd__or2_1 _13385_ (.A(_06076_),
    .B(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__nor2_1 _13386_ (.A(_05862_),
    .B(_06035_),
    .Y(_06143_));
 sky130_fd_sc_hd__xnor2_1 _13387_ (.A(_06037_),
    .B(_06036_),
    .Y(_06144_));
 sky130_fd_sc_hd__and3_1 _13388_ (.A(_06099_),
    .B(_06143_),
    .C(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__a21oi_1 _13389_ (.A1(_06099_),
    .A2(_06143_),
    .B1(_06144_),
    .Y(_06146_));
 sky130_fd_sc_hd__or2_1 _13390_ (.A(_06145_),
    .B(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__or2_1 _13391_ (.A(_05503_),
    .B(_05992_),
    .X(_06148_));
 sky130_fd_sc_hd__nor2_1 _13392_ (.A(_06001_),
    .B(_05992_),
    .Y(_06149_));
 sky130_fd_sc_hd__or2_1 _13393_ (.A(_05503_),
    .B(_05987_),
    .X(_06150_));
 sky130_fd_sc_hd__xnor2_1 _13394_ (.A(_06149_),
    .B(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__or3b_1 _13395_ (.A(_06008_),
    .B(_05995_),
    .C_N(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__o31a_1 _13396_ (.A1(_06001_),
    .A2(_05988_),
    .A3(_06148_),
    .B1(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__o21ba_1 _13397_ (.A1(_06147_),
    .A2(_06153_),
    .B1_N(_06145_),
    .X(_06154_));
 sky130_fd_sc_hd__xnor2_1 _13398_ (.A(_05902_),
    .B(_05903_),
    .Y(_06155_));
 sky130_fd_sc_hd__clkbuf_4 _13399_ (.A(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__nor2_1 _13400_ (.A(_05990_),
    .B(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__nand2_1 _13401_ (.A(_06072_),
    .B(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__nor2_1 _13402_ (.A(_05990_),
    .B(_06071_),
    .Y(_06159_));
 sky130_fd_sc_hd__or2_1 _13403_ (.A(_05996_),
    .B(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__a21oi_1 _13404_ (.A1(_06073_),
    .A2(_06160_),
    .B1(_06097_),
    .Y(_06161_));
 sky130_fd_sc_hd__or2_1 _13405_ (.A(_06158_),
    .B(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__xor2_1 _13406_ (.A(_06142_),
    .B(_06154_),
    .X(_06163_));
 sky130_fd_sc_hd__or2b_1 _13407_ (.A(_06162_),
    .B_N(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__o21ai_1 _13408_ (.A1(_06142_),
    .A2(_06154_),
    .B1(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__xnor2_1 _13409_ (.A(_06126_),
    .B(_06130_),
    .Y(_06166_));
 sky130_fd_sc_hd__o2bb2a_1 _13410_ (.A1_N(_05549_),
    .A2_N(_06055_),
    .B1(_05610_),
    .B2(_06061_),
    .X(_06167_));
 sky130_fd_sc_hd__a21oi_1 _13411_ (.A1(_06099_),
    .A2(_06143_),
    .B1(_06167_),
    .Y(_06168_));
 sky130_fd_sc_hd__nand2_1 _13412_ (.A(_06123_),
    .B(_06128_),
    .Y(_06169_));
 sky130_fd_sc_hd__a21o_1 _13413_ (.A1(_05538_),
    .A2(_06098_),
    .B1(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__xor2_1 _13414_ (.A(_06123_),
    .B(_06128_),
    .X(_06171_));
 sky130_fd_sc_hd__and2_1 _13415_ (.A(_05538_),
    .B(_06055_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_2 _13416_ (.A(_06172_),
    .X(_06173_));
 sky130_fd_sc_hd__and2_1 _13417_ (.A(_06171_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__a21oi_1 _13418_ (.A1(_06168_),
    .A2(_06170_),
    .B1(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__or2_1 _13419_ (.A(_06166_),
    .B(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__xor2_1 _13420_ (.A(_06147_),
    .B(_06153_),
    .X(_06177_));
 sky130_fd_sc_hd__nand2_1 _13421_ (.A(_06166_),
    .B(_06175_),
    .Y(_06178_));
 sky130_fd_sc_hd__and2_1 _13422_ (.A(_06176_),
    .B(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__nand2_1 _13423_ (.A(_06177_),
    .B(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__xnor2_1 _13424_ (.A(_06120_),
    .B(_06133_),
    .Y(_06181_));
 sky130_fd_sc_hd__a21o_1 _13425_ (.A1(_06176_),
    .A2(_06180_),
    .B1(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__xnor2_1 _13426_ (.A(_06162_),
    .B(_06163_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand3_1 _13427_ (.A(_06181_),
    .B(_06176_),
    .C(_06180_),
    .Y(_06184_));
 sky130_fd_sc_hd__and2_1 _13428_ (.A(_06182_),
    .B(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__nand2_1 _13429_ (.A(_06183_),
    .B(_06185_),
    .Y(_06186_));
 sky130_fd_sc_hd__xnor2_1 _13430_ (.A(_06118_),
    .B(_06137_),
    .Y(_06187_));
 sky130_fd_sc_hd__a21oi_1 _13431_ (.A1(_06182_),
    .A2(_06186_),
    .B1(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__and3_1 _13432_ (.A(_06187_),
    .B(_06182_),
    .C(_06186_),
    .X(_06189_));
 sky130_fd_sc_hd__nor2_1 _13433_ (.A(_06188_),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__a21oi_1 _13434_ (.A1(_06165_),
    .A2(_06190_),
    .B1(_06188_),
    .Y(_06191_));
 sky130_fd_sc_hd__nor2_1 _13435_ (.A(_06140_),
    .B(_06191_),
    .Y(_06192_));
 sky130_fd_sc_hd__nand2_1 _13436_ (.A(_05997_),
    .B(_06095_),
    .Y(_06193_));
 sky130_fd_sc_hd__o21ai_1 _13437_ (.A1(_06085_),
    .A2(_06094_),
    .B1(_06193_),
    .Y(_06194_));
 sky130_fd_sc_hd__a211o_1 _13438_ (.A1(_05480_),
    .A2(_06098_),
    .B1(_06106_),
    .C1(_06086_),
    .X(_06195_));
 sky130_fd_sc_hd__and3_1 _13439_ (.A(_05616_),
    .B(_05768_),
    .C(_06056_),
    .X(_06196_));
 sky130_fd_sc_hd__a21o_1 _13440_ (.A1(_06104_),
    .A2(_06107_),
    .B1(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__a21o_1 _13441_ (.A1(_06195_),
    .A2(_06197_),
    .B1(_06097_),
    .X(_06198_));
 sky130_fd_sc_hd__nor2_1 _13442_ (.A(_06080_),
    .B(_06081_),
    .Y(_06199_));
 sky130_fd_sc_hd__nand2_1 _13443_ (.A(_06080_),
    .B(_06081_),
    .Y(_06200_));
 sky130_fd_sc_hd__o31a_1 _13444_ (.A1(_06082_),
    .A2(_06110_),
    .A3(_06199_),
    .B1(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__xnor2_1 _13445_ (.A(_06198_),
    .B(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__o21a_1 _13446_ (.A1(_06102_),
    .A2(_06112_),
    .B1(_06114_),
    .X(_06203_));
 sky130_fd_sc_hd__xor2_1 _13447_ (.A(_06202_),
    .B(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__xnor2_1 _13448_ (.A(_06194_),
    .B(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__nor2_1 _13449_ (.A(_06116_),
    .B(_06138_),
    .Y(_06206_));
 sky130_fd_sc_hd__a21oi_1 _13450_ (.A1(_06079_),
    .A2(_06139_),
    .B1(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__nor2_1 _13451_ (.A(_06205_),
    .B(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__and2_1 _13452_ (.A(_06205_),
    .B(_06207_),
    .X(_06209_));
 sky130_fd_sc_hd__nor2_1 _13453_ (.A(_06208_),
    .B(_06209_),
    .Y(_06210_));
 sky130_fd_sc_hd__and2_1 _13454_ (.A(_06192_),
    .B(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__and3_1 _13455_ (.A(_06056_),
    .B(_06200_),
    .C(_06197_),
    .X(_06212_));
 sky130_fd_sc_hd__a21oi_1 _13456_ (.A1(_05768_),
    .A2(_06098_),
    .B1(_06106_),
    .Y(_06213_));
 sky130_fd_sc_hd__nor2_1 _13457_ (.A(_06196_),
    .B(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__nor2_1 _13458_ (.A(_06212_),
    .B(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__nand2_1 _13459_ (.A(_06212_),
    .B(_06214_),
    .Y(_06216_));
 sky130_fd_sc_hd__nand3_1 _13460_ (.A(_06198_),
    .B(_06201_),
    .C(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__inv_2 _13461_ (.A(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__o21a_1 _13462_ (.A1(_06215_),
    .A2(_06218_),
    .B1(_06200_),
    .X(_06219_));
 sky130_fd_sc_hd__nor2_1 _13463_ (.A(_06202_),
    .B(_06203_),
    .Y(_06220_));
 sky130_fd_sc_hd__a21oi_1 _13464_ (.A1(_06194_),
    .A2(_06204_),
    .B1(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__or2_1 _13465_ (.A(_06219_),
    .B(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__nand2_1 _13466_ (.A(_06219_),
    .B(_06221_),
    .Y(_06223_));
 sky130_fd_sc_hd__and3_1 _13467_ (.A(_06208_),
    .B(_06222_),
    .C(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__and2_1 _13468_ (.A(_06222_),
    .B(_06223_),
    .X(_06225_));
 sky130_fd_sc_hd__nor2_1 _13469_ (.A(_06208_),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__nor2_1 _13470_ (.A(_06224_),
    .B(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__xnor2_1 _13471_ (.A(_06165_),
    .B(_06190_),
    .Y(_06228_));
 sky130_fd_sc_hd__xnor2_1 _13472_ (.A(_06183_),
    .B(_06185_),
    .Y(_06229_));
 sky130_fd_sc_hd__buf_2 _13473_ (.A(_05902_),
    .X(_06230_));
 sky130_fd_sc_hd__or2_1 _13474_ (.A(_05472_),
    .B(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__nor3_2 _13475_ (.A(_05990_),
    .B(_06156_),
    .C(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__or2_1 _13476_ (.A(_06072_),
    .B(_06157_),
    .X(_06233_));
 sky130_fd_sc_hd__and2_1 _13477_ (.A(_06158_),
    .B(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__nand2_1 _13478_ (.A(_06232_),
    .B(_06234_),
    .Y(_06235_));
 sky130_fd_sc_hd__nand2_1 _13479_ (.A(_06158_),
    .B(_06161_),
    .Y(_06236_));
 sky130_fd_sc_hd__nand2_1 _13480_ (.A(_06162_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__or3_1 _13481_ (.A(_05301_),
    .B(_05527_),
    .C(_06055_),
    .X(_06238_));
 sky130_fd_sc_hd__xor2_1 _13482_ (.A(_06143_),
    .B(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__or3_1 _13483_ (.A(_05862_),
    .B(_06061_),
    .C(_06238_),
    .X(_06240_));
 sky130_fd_sc_hd__o31ai_2 _13484_ (.A1(_06103_),
    .A2(_05988_),
    .A3(_06239_),
    .B1(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__o21bai_1 _13485_ (.A1(_06008_),
    .A2(_05995_),
    .B1_N(_06151_),
    .Y(_06242_));
 sky130_fd_sc_hd__and2_1 _13486_ (.A(_06152_),
    .B(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__xnor2_1 _13487_ (.A(_06241_),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__nor2_1 _13488_ (.A(_05503_),
    .B(_05995_),
    .Y(_06245_));
 sky130_fd_sc_hd__nor2_1 _13489_ (.A(_06008_),
    .B(_06071_),
    .Y(_06246_));
 sky130_fd_sc_hd__nor2_1 _13490_ (.A(_06001_),
    .B(_05995_),
    .Y(_06247_));
 sky130_fd_sc_hd__xnor2_1 _13491_ (.A(_06148_),
    .B(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__a22oi_2 _13492_ (.A1(_06149_),
    .A2(_06245_),
    .B1(_06246_),
    .B2(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand2_1 _13493_ (.A(_06241_),
    .B(_06243_),
    .Y(_06250_));
 sky130_fd_sc_hd__o21a_1 _13494_ (.A1(_06244_),
    .A2(_06249_),
    .B1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__xor2_1 _13495_ (.A(_06237_),
    .B(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__xnor2_1 _13496_ (.A(_06235_),
    .B(_06252_),
    .Y(_06253_));
 sky130_fd_sc_hd__xnor2_1 _13497_ (.A(_06177_),
    .B(_06179_),
    .Y(_06254_));
 sky130_fd_sc_hd__xor2_1 _13498_ (.A(_06244_),
    .B(_06249_),
    .X(_06255_));
 sky130_fd_sc_hd__and2b_1 _13499_ (.A_N(_06174_),
    .B(_06170_),
    .X(_06256_));
 sky130_fd_sc_hd__xnor2_1 _13500_ (.A(_06168_),
    .B(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__nor2_1 _13501_ (.A(_06103_),
    .B(_05988_),
    .Y(_06258_));
 sky130_fd_sc_hd__xnor2_1 _13502_ (.A(_06239_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__xnor2_1 _13503_ (.A(_06171_),
    .B(_06173_),
    .Y(_06260_));
 sky130_fd_sc_hd__o21ai_1 _13504_ (.A1(_06121_),
    .A2(_06035_),
    .B1(_06123_),
    .Y(_06261_));
 sky130_fd_sc_hd__or3_1 _13505_ (.A(_06122_),
    .B(_06035_),
    .C(_06128_),
    .X(_06262_));
 sky130_fd_sc_hd__a21boi_1 _13506_ (.A1(_06173_),
    .A2(_06261_),
    .B1_N(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__xor2_1 _13507_ (.A(_06260_),
    .B(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__nor2_1 _13508_ (.A(_06260_),
    .B(_06263_),
    .Y(_06265_));
 sky130_fd_sc_hd__a21oi_1 _13509_ (.A1(_06259_),
    .A2(_06264_),
    .B1(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__xor2_1 _13510_ (.A(_06257_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__nor2_1 _13511_ (.A(_06257_),
    .B(_06266_),
    .Y(_06268_));
 sky130_fd_sc_hd__a21oi_1 _13512_ (.A1(_06255_),
    .A2(_06267_),
    .B1(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__xor2_1 _13513_ (.A(_06254_),
    .B(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__nor2_1 _13514_ (.A(_06254_),
    .B(_06269_),
    .Y(_06271_));
 sky130_fd_sc_hd__a21oi_1 _13515_ (.A1(_06253_),
    .A2(_06270_),
    .B1(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__xnor2_1 _13516_ (.A(_06229_),
    .B(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nor2_1 _13517_ (.A(_06237_),
    .B(_06251_),
    .Y(_06274_));
 sky130_fd_sc_hd__a31o_1 _13518_ (.A1(_06232_),
    .A2(_06234_),
    .A3(_06252_),
    .B1(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__or2b_1 _13519_ (.A(_06273_),
    .B_N(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__o21a_1 _13520_ (.A1(_06229_),
    .A2(_06272_),
    .B1(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__nor2_1 _13521_ (.A(_06228_),
    .B(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__and2_1 _13522_ (.A(_06140_),
    .B(_06191_),
    .X(_06279_));
 sky130_fd_sc_hd__nor2_1 _13523_ (.A(_06192_),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__nand2_1 _13524_ (.A(_06278_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nor2_1 _13525_ (.A(_06192_),
    .B(_06210_),
    .Y(_06282_));
 sky130_fd_sc_hd__or2_1 _13526_ (.A(_06211_),
    .B(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__nand2_1 _13527_ (.A(_06281_),
    .B(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__or2_1 _13528_ (.A(_06278_),
    .B(_06280_),
    .X(_06285_));
 sky130_fd_sc_hd__xor2_1 _13529_ (.A(_06275_),
    .B(_06273_),
    .X(_06286_));
 sky130_fd_sc_hd__xnor2_1 _13530_ (.A(_06246_),
    .B(_06248_),
    .Y(_06287_));
 sky130_fd_sc_hd__and2_1 _13531_ (.A(_05697_),
    .B(_06055_),
    .X(_06288_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13532_ (.A(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__nor2_1 _13533_ (.A(_05862_),
    .B(_05988_),
    .Y(_06290_));
 sky130_fd_sc_hd__xnor2_1 _13534_ (.A(_06289_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__nand2_1 _13535_ (.A(_06289_),
    .B(_06290_),
    .Y(_06292_));
 sky130_fd_sc_hd__o31ai_2 _13536_ (.A1(_06103_),
    .A2(_05992_),
    .A3(_06291_),
    .B1(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__or2b_1 _13537_ (.A(_06287_),
    .B_N(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__xor2_1 _13538_ (.A(_06293_),
    .B(_06287_),
    .X(_06295_));
 sky130_fd_sc_hd__nor2_1 _13539_ (.A(_05503_),
    .B(_06071_),
    .Y(_06296_));
 sky130_fd_sc_hd__or2_1 _13540_ (.A(_06008_),
    .B(_06156_),
    .X(_06297_));
 sky130_fd_sc_hd__nor2_1 _13541_ (.A(_06001_),
    .B(_06071_),
    .Y(_06298_));
 sky130_fd_sc_hd__nor2_1 _13542_ (.A(_06245_),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__a21o_1 _13543_ (.A1(_06247_),
    .A2(_06296_),
    .B1(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__o2bb2a_1 _13544_ (.A1_N(_06247_),
    .A2_N(_06296_),
    .B1(_06297_),
    .B2(_06300_),
    .X(_06301_));
 sky130_fd_sc_hd__or2_1 _13545_ (.A(_06295_),
    .B(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__xnor2_1 _13546_ (.A(_06232_),
    .B(_06234_),
    .Y(_06303_));
 sky130_fd_sc_hd__a21oi_2 _13547_ (.A1(_06294_),
    .A2(_06302_),
    .B1(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__xnor2_1 _13548_ (.A(_06253_),
    .B(_06270_),
    .Y(_06305_));
 sky130_fd_sc_hd__and3_1 _13549_ (.A(_06294_),
    .B(_06302_),
    .C(_06303_),
    .X(_06306_));
 sky130_fd_sc_hd__nor2_1 _13550_ (.A(_06304_),
    .B(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__xnor2_1 _13551_ (.A(_06255_),
    .B(_06267_),
    .Y(_06308_));
 sky130_fd_sc_hd__xor2_1 _13552_ (.A(_06295_),
    .B(_06301_),
    .X(_06309_));
 sky130_fd_sc_hd__xnor2_1 _13553_ (.A(_06259_),
    .B(_06264_),
    .Y(_06310_));
 sky130_fd_sc_hd__nor2_1 _13554_ (.A(_06103_),
    .B(_05992_),
    .Y(_06311_));
 sky130_fd_sc_hd__xnor2_1 _13555_ (.A(_06291_),
    .B(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__nand3_1 _13556_ (.A(_06173_),
    .B(_06262_),
    .C(_06261_),
    .Y(_06313_));
 sky130_fd_sc_hd__a21o_1 _13557_ (.A1(_06262_),
    .A2(_06261_),
    .B1(_06173_),
    .X(_06314_));
 sky130_fd_sc_hd__o22ai_2 _13558_ (.A1(_06121_),
    .A2(_05988_),
    .B1(_06061_),
    .B2(_06122_),
    .Y(_06315_));
 sky130_fd_sc_hd__or4_1 _13559_ (.A(_06121_),
    .B(_06122_),
    .C(_05987_),
    .D(_06035_),
    .X(_06316_));
 sky130_fd_sc_hd__a21bo_1 _13560_ (.A1(_06173_),
    .A2(_06315_),
    .B1_N(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__a21o_1 _13561_ (.A1(_06313_),
    .A2(_06314_),
    .B1(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__nand3_1 _13562_ (.A(_06313_),
    .B(_06314_),
    .C(_06317_),
    .Y(_06319_));
 sky130_fd_sc_hd__a21boi_1 _13563_ (.A1(_06312_),
    .A2(_06318_),
    .B1_N(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__xor2_1 _13564_ (.A(_06310_),
    .B(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__nor2_1 _13565_ (.A(_06310_),
    .B(_06320_),
    .Y(_06322_));
 sky130_fd_sc_hd__a21oi_1 _13566_ (.A1(_06309_),
    .A2(_06321_),
    .B1(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__xor2_1 _13567_ (.A(_06308_),
    .B(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__nor2_1 _13568_ (.A(_06308_),
    .B(_06323_),
    .Y(_06325_));
 sky130_fd_sc_hd__a21oi_1 _13569_ (.A1(_06307_),
    .A2(_06324_),
    .B1(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__xor2_1 _13570_ (.A(_06305_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__nor2_1 _13571_ (.A(_06305_),
    .B(_06326_),
    .Y(_06328_));
 sky130_fd_sc_hd__a21oi_1 _13572_ (.A1(_06304_),
    .A2(_06327_),
    .B1(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__nor2_1 _13573_ (.A(_06286_),
    .B(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__xor2_1 _13574_ (.A(_06228_),
    .B(_06277_),
    .X(_06331_));
 sky130_fd_sc_hd__nand2_1 _13575_ (.A(_06330_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__a21bo_1 _13576_ (.A1(_06281_),
    .A2(_06285_),
    .B1_N(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__and2_1 _13577_ (.A(_06286_),
    .B(_06329_),
    .X(_06334_));
 sky130_fd_sc_hd__nor2_1 _13578_ (.A(_06330_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__xnor2_1 _13579_ (.A(_06297_),
    .B(_06300_),
    .Y(_06336_));
 sky130_fd_sc_hd__nor2_1 _13580_ (.A(_05527_),
    .B(_05992_),
    .Y(_06337_));
 sky130_fd_sc_hd__nor2_1 _13581_ (.A(_05862_),
    .B(_05992_),
    .Y(_06338_));
 sky130_fd_sc_hd__or2_1 _13582_ (.A(_06289_),
    .B(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__nor2_1 _13583_ (.A(_06103_),
    .B(_05995_),
    .Y(_06340_));
 sky130_fd_sc_hd__a22o_1 _13584_ (.A1(_06125_),
    .A2(_06337_),
    .B1(_06339_),
    .B2(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__or2b_1 _13585_ (.A(_06336_),
    .B_N(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__xor2_1 _13586_ (.A(_06341_),
    .B(_06336_),
    .X(_06343_));
 sky130_fd_sc_hd__nor2_1 _13587_ (.A(_06001_),
    .B(_06156_),
    .Y(_06344_));
 sky130_fd_sc_hd__or2_1 _13588_ (.A(_06008_),
    .B(_06230_),
    .X(_06345_));
 sky130_fd_sc_hd__nor2_1 _13589_ (.A(_05503_),
    .B(_06156_),
    .Y(_06346_));
 sky130_fd_sc_hd__nor2_1 _13590_ (.A(_06296_),
    .B(_06344_),
    .Y(_06347_));
 sky130_fd_sc_hd__a21o_1 _13591_ (.A1(_06298_),
    .A2(_06346_),
    .B1(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__nor2_1 _13592_ (.A(_06345_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__a21oi_1 _13593_ (.A1(_06296_),
    .A2(_06344_),
    .B1(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__or2_1 _13594_ (.A(_06343_),
    .B(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__o22a_1 _13595_ (.A1(_05990_),
    .A2(_06230_),
    .B1(_06156_),
    .B2(_05472_),
    .X(_06352_));
 sky130_fd_sc_hd__or2_1 _13596_ (.A(_06232_),
    .B(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__a21oi_2 _13597_ (.A1(_06342_),
    .A2(_06351_),
    .B1(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__xnor2_1 _13598_ (.A(_06307_),
    .B(_06324_),
    .Y(_06355_));
 sky130_fd_sc_hd__and3_1 _13599_ (.A(_06342_),
    .B(_06351_),
    .C(_06353_),
    .X(_06356_));
 sky130_fd_sc_hd__nor2_1 _13600_ (.A(_06354_),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__xnor2_1 _13601_ (.A(_06309_),
    .B(_06321_),
    .Y(_06358_));
 sky130_fd_sc_hd__xor2_1 _13602_ (.A(_06343_),
    .B(_06350_),
    .X(_06359_));
 sky130_fd_sc_hd__nand3_1 _13603_ (.A(_06319_),
    .B(_06312_),
    .C(_06318_),
    .Y(_06360_));
 sky130_fd_sc_hd__a21o_1 _13604_ (.A1(_06319_),
    .A2(_06318_),
    .B1(_06312_),
    .X(_06361_));
 sky130_fd_sc_hd__xnor2_1 _13605_ (.A(_06289_),
    .B(_06338_),
    .Y(_06362_));
 sky130_fd_sc_hd__xnor2_1 _13606_ (.A(_06362_),
    .B(_06340_),
    .Y(_06363_));
 sky130_fd_sc_hd__nand3_1 _13607_ (.A(_06173_),
    .B(_06316_),
    .C(_06315_),
    .Y(_06364_));
 sky130_fd_sc_hd__a21o_1 _13608_ (.A1(_06316_),
    .A2(_06315_),
    .B1(_06173_),
    .X(_06365_));
 sky130_fd_sc_hd__or2_1 _13609_ (.A(_06122_),
    .B(_05991_),
    .X(_06366_));
 sky130_fd_sc_hd__nor3_1 _13610_ (.A(_06121_),
    .B(_05987_),
    .C(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__nor2_1 _13611_ (.A(_06121_),
    .B(_05991_),
    .Y(_06368_));
 sky130_fd_sc_hd__o21ba_1 _13612_ (.A1(_06122_),
    .A2(_05987_),
    .B1_N(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__or4_1 _13613_ (.A(_05805_),
    .B(_06035_),
    .C(_06367_),
    .D(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__or2b_1 _13614_ (.A(_06367_),
    .B_N(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__a21o_1 _13615_ (.A1(_06364_),
    .A2(_06365_),
    .B1(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__nand3_1 _13616_ (.A(_06364_),
    .B(_06365_),
    .C(_06371_),
    .Y(_06373_));
 sky130_fd_sc_hd__a21bo_1 _13617_ (.A1(_06363_),
    .A2(_06372_),
    .B1_N(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__a21o_1 _13618_ (.A1(_06360_),
    .A2(_06361_),
    .B1(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__nand3_1 _13619_ (.A(_06360_),
    .B(_06361_),
    .C(_06374_),
    .Y(_06376_));
 sky130_fd_sc_hd__a21boi_1 _13620_ (.A1(_06359_),
    .A2(_06375_),
    .B1_N(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__xor2_1 _13621_ (.A(_06358_),
    .B(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__nor2_1 _13622_ (.A(_06358_),
    .B(_06377_),
    .Y(_06379_));
 sky130_fd_sc_hd__a21oi_1 _13623_ (.A1(_06357_),
    .A2(_06378_),
    .B1(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__xor2_1 _13624_ (.A(_06355_),
    .B(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__xnor2_1 _13625_ (.A(_06354_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__nor2_1 _13626_ (.A(_05527_),
    .B(_05995_),
    .Y(_06383_));
 sky130_fd_sc_hd__nor2_1 _13627_ (.A(_05862_),
    .B(_05995_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand3_1 _13628_ (.A(_05697_),
    .B(_06056_),
    .C(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__a21o_1 _13629_ (.A1(_05697_),
    .A2(_06055_),
    .B1(_06384_),
    .X(_06386_));
 sky130_fd_sc_hd__nor2_1 _13630_ (.A(_06103_),
    .B(_06071_),
    .Y(_06387_));
 sky130_fd_sc_hd__and3_1 _13631_ (.A(_06385_),
    .B(_06386_),
    .C(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__a21oi_1 _13632_ (.A1(_06125_),
    .A2(_06383_),
    .B1(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__and2_1 _13633_ (.A(_06345_),
    .B(_06348_),
    .X(_06390_));
 sky130_fd_sc_hd__nor2_1 _13634_ (.A(_06001_),
    .B(_06230_),
    .Y(_06391_));
 sky130_fd_sc_hd__and2_1 _13635_ (.A(_06346_),
    .B(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__nor2_1 _13636_ (.A(_06349_),
    .B(_06390_),
    .Y(_06393_));
 sky130_fd_sc_hd__xnor2_1 _13637_ (.A(_06389_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2_1 _13638_ (.A(_06392_),
    .B(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__o31a_1 _13639_ (.A1(_06349_),
    .A2(_06389_),
    .A3(_06390_),
    .B1(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__nor2_1 _13640_ (.A(_06231_),
    .B(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__xnor2_1 _13641_ (.A(_06357_),
    .B(_06378_),
    .Y(_06398_));
 sky130_fd_sc_hd__xor2_1 _13642_ (.A(_06231_),
    .B(_06396_),
    .X(_06399_));
 sky130_fd_sc_hd__nand3_1 _13643_ (.A(_06376_),
    .B(_06359_),
    .C(_06375_),
    .Y(_06400_));
 sky130_fd_sc_hd__a21o_1 _13644_ (.A1(_06376_),
    .A2(_06375_),
    .B1(_06359_),
    .X(_06401_));
 sky130_fd_sc_hd__xnor2_1 _13645_ (.A(_06392_),
    .B(_06394_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand3_1 _13646_ (.A(_06373_),
    .B(_06363_),
    .C(_06372_),
    .Y(_06403_));
 sky130_fd_sc_hd__a21o_1 _13647_ (.A1(_06373_),
    .A2(_06372_),
    .B1(_06363_),
    .X(_06404_));
 sky130_fd_sc_hd__a21oi_1 _13648_ (.A1(_06385_),
    .A2(_06386_),
    .B1(_06387_),
    .Y(_06405_));
 sky130_fd_sc_hd__nor2_1 _13649_ (.A(_06388_),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__o22ai_1 _13650_ (.A1(_05805_),
    .A2(_06061_),
    .B1(_06367_),
    .B2(_06369_),
    .Y(_06407_));
 sky130_fd_sc_hd__nor2_1 _13651_ (.A(_06122_),
    .B(_05994_),
    .Y(_06408_));
 sky130_fd_sc_hd__nor2_1 _13652_ (.A(_05805_),
    .B(_05987_),
    .Y(_06409_));
 sky130_fd_sc_hd__nor2_1 _13653_ (.A(_06121_),
    .B(_05994_),
    .Y(_06410_));
 sky130_fd_sc_hd__xnor2_1 _13654_ (.A(_06366_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__a22o_1 _13655_ (.A1(_06368_),
    .A2(_06408_),
    .B1(_06409_),
    .B2(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__and3_1 _13656_ (.A(_06370_),
    .B(_06407_),
    .C(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__a21oi_1 _13657_ (.A1(_06370_),
    .A2(_06407_),
    .B1(_06412_),
    .Y(_06414_));
 sky130_fd_sc_hd__nor2_1 _13658_ (.A(_06413_),
    .B(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__a21o_1 _13659_ (.A1(_06406_),
    .A2(_06415_),
    .B1(_06413_),
    .X(_06416_));
 sky130_fd_sc_hd__a21oi_1 _13660_ (.A1(_06403_),
    .A2(_06404_),
    .B1(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__and3_1 _13661_ (.A(_06403_),
    .B(_06404_),
    .C(_06416_),
    .X(_06418_));
 sky130_fd_sc_hd__o21bai_1 _13662_ (.A1(_06402_),
    .A2(_06417_),
    .B1_N(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__a21o_1 _13663_ (.A1(_06400_),
    .A2(_06401_),
    .B1(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__and3_1 _13664_ (.A(_06400_),
    .B(_06401_),
    .C(_06419_),
    .X(_06421_));
 sky130_fd_sc_hd__a21o_1 _13665_ (.A1(_06399_),
    .A2(_06420_),
    .B1(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__xnor2_1 _13666_ (.A(_06398_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__and2b_1 _13667_ (.A_N(_06398_),
    .B(_06422_),
    .X(_06424_));
 sky130_fd_sc_hd__a21o_1 _13668_ (.A1(_06397_),
    .A2(_06423_),
    .B1(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__and2b_1 _13669_ (.A_N(_06382_),
    .B(_06425_),
    .X(_06426_));
 sky130_fd_sc_hd__xnor2_1 _13670_ (.A(_06304_),
    .B(_06327_),
    .Y(_06427_));
 sky130_fd_sc_hd__nor2_1 _13671_ (.A(_06355_),
    .B(_06380_),
    .Y(_06428_));
 sky130_fd_sc_hd__a21oi_1 _13672_ (.A1(_06354_),
    .A2(_06381_),
    .B1(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__xor2_1 _13673_ (.A(_06427_),
    .B(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__and2_1 _13674_ (.A(_06426_),
    .B(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__nor2_1 _13675_ (.A(_06427_),
    .B(_06429_),
    .Y(_06432_));
 sky130_fd_sc_hd__nor2_1 _13676_ (.A(_06432_),
    .B(_06431_),
    .Y(_06433_));
 sky130_fd_sc_hd__xnor2_1 _13677_ (.A(_06335_),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__xnor2_2 _13678_ (.A(_06382_),
    .B(_06425_),
    .Y(_06435_));
 sky130_fd_sc_hd__xor2_1 _13679_ (.A(_06397_),
    .B(_06423_),
    .X(_06436_));
 sky130_fd_sc_hd__and2b_1 _13680_ (.A_N(_06421_),
    .B(_06420_),
    .X(_06437_));
 sky130_fd_sc_hd__xnor2_1 _13681_ (.A(_06399_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__nor2_1 _13682_ (.A(_05527_),
    .B(_06071_),
    .Y(_06439_));
 sky130_fd_sc_hd__or3b_1 _13683_ (.A(_05862_),
    .B(_06035_),
    .C_N(_06439_),
    .X(_06440_));
 sky130_fd_sc_hd__o22ai_1 _13684_ (.A1(_05527_),
    .A2(_06061_),
    .B1(_06071_),
    .B2(_05862_),
    .Y(_06441_));
 sky130_fd_sc_hd__nor2_1 _13685_ (.A(_06103_),
    .B(_06156_),
    .Y(_06442_));
 sky130_fd_sc_hd__nand3_1 _13686_ (.A(_06440_),
    .B(_06441_),
    .C(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__or2_1 _13687_ (.A(_06346_),
    .B(_06391_),
    .X(_06444_));
 sky130_fd_sc_hd__or2b_1 _13688_ (.A(_06392_),
    .B_N(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__a21oi_1 _13689_ (.A1(_06440_),
    .A2(_06443_),
    .B1(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__or3_1 _13690_ (.A(_06418_),
    .B(_06402_),
    .C(_06417_),
    .X(_06447_));
 sky130_fd_sc_hd__o21ai_1 _13691_ (.A1(_06418_),
    .A2(_06417_),
    .B1(_06402_),
    .Y(_06448_));
 sky130_fd_sc_hd__and3_1 _13692_ (.A(_06440_),
    .B(_06443_),
    .C(_06445_),
    .X(_06449_));
 sky130_fd_sc_hd__nor2_1 _13693_ (.A(_06446_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__xor2_1 _13694_ (.A(_06406_),
    .B(_06415_),
    .X(_06451_));
 sky130_fd_sc_hd__xnor2_1 _13695_ (.A(_06409_),
    .B(_06411_),
    .Y(_06452_));
 sky130_fd_sc_hd__nor2_1 _13696_ (.A(_06122_),
    .B(_06070_),
    .Y(_06453_));
 sky130_fd_sc_hd__nor2_1 _13697_ (.A(_05805_),
    .B(_05992_),
    .Y(_06454_));
 sky130_fd_sc_hd__nor2_1 _13698_ (.A(_06121_),
    .B(_06070_),
    .Y(_06455_));
 sky130_fd_sc_hd__xor2_1 _13699_ (.A(_06408_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__a22o_1 _13700_ (.A1(_06410_),
    .A2(_06453_),
    .B1(_06454_),
    .B2(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__or2b_1 _13701_ (.A(_06452_),
    .B_N(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__a21o_1 _13702_ (.A1(_06440_),
    .A2(_06441_),
    .B1(_06442_),
    .X(_06459_));
 sky130_fd_sc_hd__xnor2_1 _13703_ (.A(_06452_),
    .B(_06457_),
    .Y(_06460_));
 sky130_fd_sc_hd__nand3_1 _13704_ (.A(_06443_),
    .B(_06459_),
    .C(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__nand2_1 _13705_ (.A(_06458_),
    .B(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__xor2_1 _13706_ (.A(_06451_),
    .B(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__and2_1 _13707_ (.A(_06451_),
    .B(_06462_),
    .X(_06464_));
 sky130_fd_sc_hd__a21o_1 _13708_ (.A1(_06450_),
    .A2(_06463_),
    .B1(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__a21o_1 _13709_ (.A1(_06447_),
    .A2(_06448_),
    .B1(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__nand3_1 _13710_ (.A(_06447_),
    .B(_06448_),
    .C(_06465_),
    .Y(_06467_));
 sky130_fd_sc_hd__a21boi_1 _13711_ (.A1(_06446_),
    .A2(_06466_),
    .B1_N(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__nor2_1 _13712_ (.A(_06438_),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__and2_1 _13713_ (.A(_06436_),
    .B(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__a21oi_1 _13714_ (.A1(_06435_),
    .A2(_06470_),
    .B1(_06426_),
    .Y(_06471_));
 sky130_fd_sc_hd__xnor2_1 _13715_ (.A(_06430_),
    .B(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__nand2_1 _13716_ (.A(_06438_),
    .B(_06468_),
    .Y(_06473_));
 sky130_fd_sc_hd__and2_1 _13717_ (.A(_06436_),
    .B(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__and3_1 _13718_ (.A(_06446_),
    .B(_06467_),
    .C(_06466_),
    .X(_06475_));
 sky130_fd_sc_hd__a21oi_1 _13719_ (.A1(_06467_),
    .A2(_06466_),
    .B1(_06446_),
    .Y(_06476_));
 sky130_fd_sc_hd__nor2_1 _13720_ (.A(_06475_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__xor2_1 _13721_ (.A(_06450_),
    .B(_06463_),
    .X(_06478_));
 sky130_fd_sc_hd__a21o_1 _13722_ (.A1(_06443_),
    .A2(_06459_),
    .B1(_06460_),
    .X(_06479_));
 sky130_fd_sc_hd__nor2_1 _13723_ (.A(_05862_),
    .B(_06156_),
    .Y(_06480_));
 sky130_fd_sc_hd__or3b_1 _13724_ (.A(_05527_),
    .B(_05987_),
    .C_N(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__o21bai_1 _13725_ (.A1(_05527_),
    .A2(_05988_),
    .B1_N(_06480_),
    .Y(_06482_));
 sky130_fd_sc_hd__nand2_1 _13726_ (.A(_06481_),
    .B(_06482_),
    .Y(_06483_));
 sky130_fd_sc_hd__nor2_1 _13727_ (.A(_06103_),
    .B(_06230_),
    .Y(_06484_));
 sky130_fd_sc_hd__xnor2_1 _13728_ (.A(_06483_),
    .B(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__xnor2_1 _13729_ (.A(_06454_),
    .B(_06456_),
    .Y(_06486_));
 sky130_fd_sc_hd__nor2_1 _13730_ (.A(_05536_),
    .B(_06155_),
    .Y(_06487_));
 sky130_fd_sc_hd__nor2_1 _13731_ (.A(_05805_),
    .B(_05995_),
    .Y(_06488_));
 sky130_fd_sc_hd__or2_1 _13732_ (.A(_05551_),
    .B(_06155_),
    .X(_06489_));
 sky130_fd_sc_hd__xnor2_1 _13733_ (.A(_06453_),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__a22o_1 _13734_ (.A1(_06455_),
    .A2(_06487_),
    .B1(_06488_),
    .B2(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__and2b_1 _13735_ (.A_N(_06486_),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__and2b_1 _13736_ (.A_N(_06491_),
    .B(_06486_),
    .X(_06493_));
 sky130_fd_sc_hd__nor2_1 _13737_ (.A(_06492_),
    .B(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__a21o_1 _13738_ (.A1(_06485_),
    .A2(_06494_),
    .B1(_06492_),
    .X(_06495_));
 sky130_fd_sc_hd__and3_1 _13739_ (.A(_06461_),
    .B(_06479_),
    .C(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__inv_2 _13740_ (.A(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__or2_1 _13741_ (.A(_05503_),
    .B(_06230_),
    .X(_06498_));
 sky130_fd_sc_hd__o31a_1 _13742_ (.A1(_06103_),
    .A2(_06230_),
    .A3(_06483_),
    .B1(_06481_),
    .X(_06499_));
 sky130_fd_sc_hd__or2_1 _13743_ (.A(_06498_),
    .B(_06499_),
    .X(_06500_));
 sky130_fd_sc_hd__nand2_1 _13744_ (.A(_06498_),
    .B(_06499_),
    .Y(_06501_));
 sky130_fd_sc_hd__and2_1 _13745_ (.A(_06500_),
    .B(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__a21o_1 _13746_ (.A1(_06461_),
    .A2(_06479_),
    .B1(_06495_),
    .X(_06503_));
 sky130_fd_sc_hd__nand3b_1 _13747_ (.A_N(_06496_),
    .B(_06502_),
    .C(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__nand2_1 _13748_ (.A(_06497_),
    .B(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__xor2_1 _13749_ (.A(_06478_),
    .B(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__or2b_1 _13750_ (.A(_06500_),
    .B_N(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__a21bo_1 _13751_ (.A1(_06478_),
    .A2(_06505_),
    .B1_N(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__and2_1 _13752_ (.A(_06477_),
    .B(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__nand2_1 _13753_ (.A(_06436_),
    .B(_06469_),
    .Y(_06510_));
 sky130_fd_sc_hd__xnor2_1 _13754_ (.A(_06500_),
    .B(_06506_),
    .Y(_06511_));
 sky130_fd_sc_hd__a21o_1 _13755_ (.A1(_06497_),
    .A2(_06503_),
    .B1(_06502_),
    .X(_06512_));
 sky130_fd_sc_hd__nor2_1 _13756_ (.A(_05862_),
    .B(_06230_),
    .Y(_06513_));
 sky130_fd_sc_hd__xnor2_1 _13757_ (.A(_06485_),
    .B(_06494_),
    .Y(_06514_));
 sky130_fd_sc_hd__nand2_1 _13758_ (.A(_06337_),
    .B(_06513_),
    .Y(_06515_));
 sky130_fd_sc_hd__or2_1 _13759_ (.A(_06337_),
    .B(_06513_),
    .X(_06516_));
 sky130_fd_sc_hd__and2_1 _13760_ (.A(_06515_),
    .B(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__xnor2_1 _13761_ (.A(_06488_),
    .B(_06490_),
    .Y(_06518_));
 sky130_fd_sc_hd__nor2_1 _13762_ (.A(_05551_),
    .B(_06230_),
    .Y(_06519_));
 sky130_fd_sc_hd__xor2_1 _13763_ (.A(_06487_),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__or3b_1 _13764_ (.A(_05805_),
    .B(_06071_),
    .C_N(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__a21bo_1 _13765_ (.A1(_06487_),
    .A2(_06519_),
    .B1_N(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__xnor2_1 _13766_ (.A(_06518_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__and2b_1 _13767_ (.A_N(_06518_),
    .B(_06522_),
    .X(_06524_));
 sky130_fd_sc_hd__a21o_1 _13768_ (.A1(_06517_),
    .A2(_06523_),
    .B1(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__and2b_1 _13769_ (.A_N(_06514_),
    .B(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__and2b_1 _13770_ (.A_N(_06525_),
    .B(_06514_),
    .X(_06527_));
 sky130_fd_sc_hd__nor2_1 _13771_ (.A(_06526_),
    .B(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__a31o_1 _13772_ (.A1(_06337_),
    .A2(_06513_),
    .A3(_06528_),
    .B1(_06526_),
    .X(_06529_));
 sky130_fd_sc_hd__a21oi_1 _13773_ (.A1(_06504_),
    .A2(_06512_),
    .B1(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__xnor2_1 _13774_ (.A(_06517_),
    .B(_06523_),
    .Y(_06531_));
 sky130_fd_sc_hd__or2_1 _13775_ (.A(_06122_),
    .B(_06230_),
    .X(_06532_));
 sky130_fd_sc_hd__or3_1 _13776_ (.A(_05805_),
    .B(_06156_),
    .C(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__o21bai_1 _13777_ (.A1(_05805_),
    .A2(_06071_),
    .B1_N(_06520_),
    .Y(_06534_));
 sky130_fd_sc_hd__nand2_1 _13778_ (.A(_06521_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__xor2_1 _13779_ (.A(_06533_),
    .B(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__nand2_1 _13780_ (.A(_06383_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__o21a_1 _13781_ (.A1(_06533_),
    .A2(_06535_),
    .B1(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__or2_1 _13782_ (.A(_06531_),
    .B(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__xor2_1 _13783_ (.A(_06515_),
    .B(_06528_),
    .X(_06540_));
 sky130_fd_sc_hd__or2_1 _13784_ (.A(_06539_),
    .B(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__and3_1 _13785_ (.A(_06504_),
    .B(_06512_),
    .C(_06529_),
    .X(_06542_));
 sky130_fd_sc_hd__o21bai_1 _13786_ (.A1(_06530_),
    .A2(_06541_),
    .B1_N(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__o21ai_1 _13787_ (.A1(_05805_),
    .A2(_06156_),
    .B1(_06532_),
    .Y(_06544_));
 sky130_fd_sc_hd__and2_1 _13788_ (.A(_06533_),
    .B(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__nand2_1 _13789_ (.A(_06439_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__o211ai_1 _13790_ (.A1(_06439_),
    .A2(_06545_),
    .B1(_05557_),
    .C1(_05904_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand2_1 _13791_ (.A(_06531_),
    .B(_06538_),
    .Y(_06548_));
 sky130_fd_sc_hd__nand2_1 _13792_ (.A(_06539_),
    .B(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__or2_1 _13793_ (.A(_06383_),
    .B(_06536_),
    .X(_06550_));
 sky130_fd_sc_hd__nand2_1 _13794_ (.A(_06537_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__a211o_1 _13795_ (.A1(_06546_),
    .A2(_06547_),
    .B1(_06549_),
    .C1(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__a21oi_1 _13796_ (.A1(_06539_),
    .A2(_06540_),
    .B1(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__nor2_1 _13797_ (.A(_06530_),
    .B(_06542_),
    .Y(_06554_));
 sky130_fd_sc_hd__a22o_1 _13798_ (.A1(_06511_),
    .A2(_06543_),
    .B1(_06553_),
    .B2(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__o221a_1 _13799_ (.A1(_06477_),
    .A2(_06508_),
    .B1(_06511_),
    .B2(_06543_),
    .C1(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__and3_1 _13800_ (.A(_06436_),
    .B(_06473_),
    .C(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__a22o_1 _13801_ (.A1(_06474_),
    .A2(_06509_),
    .B1(_06510_),
    .B2(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__and2_1 _13802_ (.A(_06435_),
    .B(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__a32o_1 _13803_ (.A1(_06435_),
    .A2(_06470_),
    .A3(_06430_),
    .B1(_06472_),
    .B2(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__a22o_1 _13804_ (.A1(_06335_),
    .A2(_06431_),
    .B1(_06434_),
    .B2(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__or2_1 _13805_ (.A(_06330_),
    .B(_06331_),
    .X(_06562_));
 sky130_fd_sc_hd__and2_1 _13806_ (.A(_06432_),
    .B(_06335_),
    .X(_06563_));
 sky130_fd_sc_hd__a21o_1 _13807_ (.A1(_06332_),
    .A2(_06562_),
    .B1(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__and3_1 _13808_ (.A(_06331_),
    .B(_06432_),
    .C(_06335_),
    .X(_06565_));
 sky130_fd_sc_hd__a21o_1 _13809_ (.A1(_06561_),
    .A2(_06564_),
    .B1(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__and3_1 _13810_ (.A(_06280_),
    .B(_06330_),
    .C(_06331_),
    .X(_06567_));
 sky130_fd_sc_hd__a21o_1 _13811_ (.A1(_06333_),
    .A2(_06566_),
    .B1(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__nor2_1 _13812_ (.A(_06281_),
    .B(_06283_),
    .Y(_06569_));
 sky130_fd_sc_hd__a21o_1 _13813_ (.A1(_06284_),
    .A2(_06568_),
    .B1(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__xor2_1 _13814_ (.A(_06227_),
    .B(_06570_),
    .X(_06571_));
 sky130_fd_sc_hd__xor2_2 _13815_ (.A(_06211_),
    .B(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__and2b_1 _13816_ (.A_N(_06569_),
    .B(_06284_),
    .X(_06573_));
 sky130_fd_sc_hd__a21o_1 _13817_ (.A1(_06573_),
    .A2(_06568_),
    .B1(_06227_),
    .X(_06574_));
 sky130_fd_sc_hd__a22o_1 _13818_ (.A1(_06227_),
    .A2(_06570_),
    .B1(_06574_),
    .B2(_06211_),
    .X(_06575_));
 sky130_fd_sc_hd__nor2_1 _13819_ (.A(_05616_),
    .B(_06056_),
    .Y(_06576_));
 sky130_fd_sc_hd__and2_1 _13820_ (.A(_06197_),
    .B(_06216_),
    .X(_06577_));
 sky130_fd_sc_hd__nor3b_1 _13821_ (.A(_06196_),
    .B(_06576_),
    .C_N(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__nor2_1 _13822_ (.A(_06218_),
    .B(_06578_),
    .Y(_06579_));
 sky130_fd_sc_hd__a31o_1 _13823_ (.A1(_06198_),
    .A2(_06201_),
    .A3(_06578_),
    .B1(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__nor2_2 _13824_ (.A(_06222_),
    .B(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__and2_1 _13825_ (.A(_06222_),
    .B(_06580_),
    .X(_06582_));
 sky130_fd_sc_hd__nor2_1 _13826_ (.A(_06581_),
    .B(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__and2_1 _13827_ (.A(_06224_),
    .B(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__nor2_1 _13828_ (.A(_06224_),
    .B(_06583_),
    .Y(_06585_));
 sky130_fd_sc_hd__nor2_1 _13829_ (.A(_06584_),
    .B(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__xor2_1 _13830_ (.A(_06575_),
    .B(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__buf_2 _13831_ (.A(_05324_),
    .X(_06588_));
 sky130_fd_sc_hd__mux2_1 _13832_ (.A0(_06572_),
    .A1(_06587_),
    .S(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__or3_1 _13833_ (.A(_06081_),
    .B(_06196_),
    .C(_06576_),
    .X(_06590_));
 sky130_fd_sc_hd__a2bb2o_1 _13834_ (.A1_N(_06577_),
    .A2_N(_06590_),
    .B1(_06578_),
    .B2(_06218_),
    .X(_06591_));
 sky130_fd_sc_hd__a21oi_2 _13835_ (.A1(_06577_),
    .A2(_06590_),
    .B1(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__xor2_2 _13836_ (.A(_06581_),
    .B(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__o21a_1 _13837_ (.A1(_06581_),
    .A2(_06584_),
    .B1(_06592_),
    .X(_06594_));
 sky130_fd_sc_hd__a31o_1 _13838_ (.A1(_06575_),
    .A2(_06586_),
    .A3(_06593_),
    .B1(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__a211o_1 _13839_ (.A1(_05696_),
    .A2(_06098_),
    .B1(_06081_),
    .C1(_06097_),
    .X(_06596_));
 sky130_fd_sc_hd__or3_2 _13840_ (.A(_06196_),
    .B(_06591_),
    .C(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__xor2_2 _13841_ (.A(_06595_),
    .B(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__a21oi_1 _13842_ (.A1(_06575_),
    .A2(_06586_),
    .B1(_06584_),
    .Y(_06599_));
 sky130_fd_sc_hd__xnor2_2 _13843_ (.A(_06593_),
    .B(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__buf_2 _13844_ (.A(_05349_),
    .X(_06601_));
 sky130_fd_sc_hd__mux2_1 _13845_ (.A0(_06598_),
    .A1(_06600_),
    .S(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__buf_2 _13846_ (.A(_05367_),
    .X(_06603_));
 sky130_fd_sc_hd__mux2_1 _13847_ (.A0(_06589_),
    .A1(_06602_),
    .S(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__and3_1 _13848_ (.A(_06601_),
    .B(_06595_),
    .C(_06597_),
    .X(_06605_));
 sky130_fd_sc_hd__o21a_1 _13849_ (.A1(_06097_),
    .A2(_06605_),
    .B1(_05447_),
    .X(_06606_));
 sky130_fd_sc_hd__a211o_1 _13850_ (.A1(_05271_),
    .A2(_06604_),
    .B1(_06606_),
    .C1(_05356_),
    .X(_06607_));
 sky130_fd_sc_hd__a211o_1 _13851_ (.A1(_06474_),
    .A2(_06509_),
    .B1(_06470_),
    .C1(_06557_),
    .X(_06608_));
 sky130_fd_sc_hd__xor2_2 _13852_ (.A(_06435_),
    .B(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__and2_1 _13853_ (.A(_06601_),
    .B(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__xnor2_1 _13854_ (.A(_06559_),
    .B(_06472_),
    .Y(_06611_));
 sky130_fd_sc_hd__nor2_1 _13855_ (.A(_05349_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__or2_1 _13856_ (.A(_06610_),
    .B(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__xnor2_2 _13857_ (.A(_06560_),
    .B(_06434_),
    .Y(_06614_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(_05324_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__and2b_1 _13859_ (.A_N(_06565_),
    .B(_06564_),
    .X(_06616_));
 sky130_fd_sc_hd__xnor2_1 _13860_ (.A(_06561_),
    .B(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__nor2_1 _13861_ (.A(_06601_),
    .B(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__nor2_1 _13862_ (.A(_06615_),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__xnor2_1 _13863_ (.A(_06573_),
    .B(_06568_),
    .Y(_06620_));
 sky130_fd_sc_hd__nor2_1 _13864_ (.A(_06601_),
    .B(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__nor2_1 _13865_ (.A(_06333_),
    .B(_06566_),
    .Y(_06622_));
 sky130_fd_sc_hd__o2bb2a_1 _13866_ (.A1_N(_06567_),
    .A2_N(_06566_),
    .B1(_06568_),
    .B2(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__nor2_1 _13867_ (.A(_06588_),
    .B(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__nor2_1 _13868_ (.A(_06621_),
    .B(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__mux2_1 _13869_ (.A0(_06619_),
    .A1(_06625_),
    .S(_06603_),
    .X(_06626_));
 sky130_fd_sc_hd__nor2_1 _13870_ (.A(_05271_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__a211o_1 _13871_ (.A1(_05410_),
    .A2(_06613_),
    .B1(_06627_),
    .C1(_05333_),
    .X(_06628_));
 sky130_fd_sc_hd__clkbuf_4 _13872_ (.A(_05272_),
    .X(_06629_));
 sky130_fd_sc_hd__clkbuf_4 _13873_ (.A(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__a31o_1 _13874_ (.A1(_05210_),
    .A2(_06607_),
    .A3(_06628_),
    .B1(_06630_),
    .X(_06631_));
 sky130_fd_sc_hd__mux2_1 _13875_ (.A0(\rbzero.wall_tracer.stepDistY[-11] ),
    .A1(_06631_),
    .S(_00004_),
    .X(_06632_));
 sky130_fd_sc_hd__clkbuf_1 _13876_ (.A(_06632_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _13877_ (.A0(_06587_),
    .A1(_06600_),
    .S(_06588_),
    .X(_06633_));
 sky130_fd_sc_hd__and3_1 _13878_ (.A(_05324_),
    .B(_06595_),
    .C(_06597_),
    .X(_06634_));
 sky130_fd_sc_hd__a21o_1 _13879_ (.A1(_06601_),
    .A2(_06598_),
    .B1(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__mux2_1 _13880_ (.A0(_06633_),
    .A1(_06635_),
    .S(_06603_),
    .X(_06636_));
 sky130_fd_sc_hd__nor2_4 _13881_ (.A(_05369_),
    .B(_05333_),
    .Y(_06637_));
 sky130_fd_sc_hd__or2_1 _13882_ (.A(_05324_),
    .B(_06617_),
    .X(_06638_));
 sky130_fd_sc_hd__or2_1 _13883_ (.A(_05349_),
    .B(_06623_),
    .X(_06639_));
 sky130_fd_sc_hd__nand2_1 _13884_ (.A(_06638_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__nor2_1 _13885_ (.A(_06588_),
    .B(_06620_),
    .Y(_06641_));
 sky130_fd_sc_hd__a21o_1 _13886_ (.A1(_06588_),
    .A2(_06572_),
    .B1(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__mux2_1 _13887_ (.A0(_06640_),
    .A1(_06642_),
    .S(_06603_),
    .X(_06643_));
 sky130_fd_sc_hd__nor2_1 _13888_ (.A(_05324_),
    .B(_06611_),
    .Y(_06644_));
 sky130_fd_sc_hd__o21bai_1 _13889_ (.A1(_06601_),
    .A2(_06614_),
    .B1_N(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__and3_1 _13890_ (.A(_06588_),
    .B(_05395_),
    .C(_06609_),
    .X(_06646_));
 sky130_fd_sc_hd__a221o_1 _13891_ (.A1(_05347_),
    .A2(_06643_),
    .B1(_06645_),
    .B2(_05410_),
    .C1(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__a21o_1 _13892_ (.A1(_06637_),
    .A2(_06647_),
    .B1(_06630_),
    .X(_06648_));
 sky130_fd_sc_hd__a31o_1 _13893_ (.A1(_05265_),
    .A2(_05271_),
    .A3(_06636_),
    .B1(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__mux2_1 _13894_ (.A0(\rbzero.wall_tracer.stepDistY[-10] ),
    .A1(_06649_),
    .S(_00004_),
    .X(_06650_));
 sky130_fd_sc_hd__clkbuf_1 _13895_ (.A(_06650_),
    .X(_00407_));
 sky130_fd_sc_hd__and2_1 _13896_ (.A(_05367_),
    .B(_06605_),
    .X(_06651_));
 sky130_fd_sc_hd__a21o_1 _13897_ (.A1(_05325_),
    .A2(_06602_),
    .B1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__nor2_1 _13898_ (.A(_06603_),
    .B(_06625_),
    .Y(_06653_));
 sky130_fd_sc_hd__a211o_1 _13899_ (.A1(_06603_),
    .A2(_06589_),
    .B1(_06653_),
    .C1(_05271_),
    .X(_06654_));
 sky130_fd_sc_hd__inv_2 _13900_ (.A(_06619_),
    .Y(_06655_));
 sky130_fd_sc_hd__o221a_1 _13901_ (.A1(_05421_),
    .A2(_06655_),
    .B1(_06613_),
    .B2(_05372_),
    .C1(_06637_),
    .X(_06656_));
 sky130_fd_sc_hd__a21o_1 _13902_ (.A1(_06654_),
    .A2(_06656_),
    .B1(_06630_),
    .X(_06657_));
 sky130_fd_sc_hd__a31o_1 _13903_ (.A1(_05265_),
    .A2(_05271_),
    .A3(_06652_),
    .B1(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__mux2_1 _13904_ (.A0(\rbzero.wall_tracer.stepDistY[-9] ),
    .A1(_06658_),
    .S(_00004_),
    .X(_06659_));
 sky130_fd_sc_hd__clkbuf_1 _13905_ (.A(_06659_),
    .X(_00408_));
 sky130_fd_sc_hd__and2_1 _13906_ (.A(_05325_),
    .B(_06642_),
    .X(_06660_));
 sky130_fd_sc_hd__a211o_1 _13907_ (.A1(_06603_),
    .A2(_06633_),
    .B1(_06660_),
    .C1(_05271_),
    .X(_06661_));
 sky130_fd_sc_hd__o221a_1 _13908_ (.A1(_05421_),
    .A2(_06640_),
    .B1(_06645_),
    .B2(_05372_),
    .C1(_06637_),
    .X(_06662_));
 sky130_fd_sc_hd__and2_1 _13909_ (.A(_05395_),
    .B(_06635_),
    .X(_06663_));
 sky130_fd_sc_hd__clkbuf_4 _13910_ (.A(_05380_),
    .X(_06664_));
 sky130_fd_sc_hd__a21o_1 _13911_ (.A1(_05324_),
    .A2(_06609_),
    .B1(_06644_),
    .X(_06665_));
 sky130_fd_sc_hd__nand2_1 _13912_ (.A(_06664_),
    .B(_06665_),
    .Y(_06666_));
 sky130_fd_sc_hd__nor2_1 _13913_ (.A(_05376_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__a21o_1 _13914_ (.A1(_05476_),
    .A2(_06667_),
    .B1(_06630_),
    .X(_06668_));
 sky130_fd_sc_hd__a221o_2 _13915_ (.A1(_06661_),
    .A2(_06662_),
    .B1(_06663_),
    .B2(_05265_),
    .C1(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__mux2_1 _13916_ (.A0(\rbzero.wall_tracer.stepDistY[-8] ),
    .A1(_06669_),
    .S(_00004_),
    .X(_06670_));
 sky130_fd_sc_hd__clkbuf_1 _13917_ (.A(_06670_),
    .X(_00409_));
 sky130_fd_sc_hd__nor2_1 _13918_ (.A(_05347_),
    .B(_06626_),
    .Y(_06671_));
 sky130_fd_sc_hd__a211o_1 _13919_ (.A1(_05347_),
    .A2(_06604_),
    .B1(_06671_),
    .C1(_05333_),
    .X(_06672_));
 sky130_fd_sc_hd__o21ai_2 _13920_ (.A1(_06097_),
    .A2(_06605_),
    .B1(_05395_),
    .Y(_06673_));
 sky130_fd_sc_hd__a21oi_1 _13921_ (.A1(_05333_),
    .A2(_06673_),
    .B1(_05369_),
    .Y(_06674_));
 sky130_fd_sc_hd__buf_2 _13922_ (.A(_05310_),
    .X(_06675_));
 sky130_fd_sc_hd__or2_1 _13923_ (.A(_06615_),
    .B(_06612_),
    .X(_06676_));
 sky130_fd_sc_hd__mux2_1 _13924_ (.A0(_06610_),
    .A1(_06676_),
    .S(_06664_),
    .X(_06677_));
 sky130_fd_sc_hd__and2_1 _13925_ (.A(_06675_),
    .B(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__a221o_2 _13926_ (.A1(_06672_),
    .A2(_06674_),
    .B1(_06678_),
    .B2(_05476_),
    .C1(_06629_),
    .X(_06679_));
 sky130_fd_sc_hd__mux2_1 _13927_ (.A0(\rbzero.wall_tracer.stepDistY[-7] ),
    .A1(_06679_),
    .S(_00004_),
    .X(_06680_));
 sky130_fd_sc_hd__clkbuf_1 _13928_ (.A(_06680_),
    .X(_00410_));
 sky130_fd_sc_hd__o21a_1 _13929_ (.A1(_05347_),
    .A2(_06643_),
    .B1(_06637_),
    .X(_06681_));
 sky130_fd_sc_hd__o21a_1 _13930_ (.A1(_05271_),
    .A2(_06636_),
    .B1(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__o21ai_1 _13931_ (.A1(_06601_),
    .A2(_06614_),
    .B1(_06638_),
    .Y(_06683_));
 sky130_fd_sc_hd__mux2_1 _13932_ (.A0(_06665_),
    .A1(_06683_),
    .S(_06664_),
    .X(_06684_));
 sky130_fd_sc_hd__a31o_1 _13933_ (.A1(_06675_),
    .A2(_05476_),
    .A3(_06684_),
    .B1(_06629_),
    .X(_06685_));
 sky130_fd_sc_hd__or2_1 _13934_ (.A(_06682_),
    .B(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__mux2_1 _13935_ (.A0(\rbzero.wall_tracer.stepDistY[-6] ),
    .A1(_06686_),
    .S(_00004_),
    .X(_06687_));
 sky130_fd_sc_hd__clkbuf_1 _13936_ (.A(_06687_),
    .X(_00411_));
 sky130_fd_sc_hd__a211o_1 _13937_ (.A1(_05325_),
    .A2(_06602_),
    .B1(_06651_),
    .C1(_05271_),
    .X(_06688_));
 sky130_fd_sc_hd__a211o_1 _13938_ (.A1(_06603_),
    .A2(_06589_),
    .B1(_06653_),
    .C1(_05347_),
    .X(_06689_));
 sky130_fd_sc_hd__nor2_1 _13939_ (.A(_06618_),
    .B(_06624_),
    .Y(_06690_));
 sky130_fd_sc_hd__nor2_1 _13940_ (.A(_06664_),
    .B(_06676_),
    .Y(_06691_));
 sky130_fd_sc_hd__a21oi_1 _13941_ (.A1(_06664_),
    .A2(_06690_),
    .B1(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__a22o_1 _13942_ (.A1(_05447_),
    .A2(_06610_),
    .B1(_06692_),
    .B2(_06675_),
    .X(_06693_));
 sky130_fd_sc_hd__a21o_1 _13943_ (.A1(_05476_),
    .A2(_06693_),
    .B1(_06629_),
    .X(_06694_));
 sky130_fd_sc_hd__a31o_2 _13944_ (.A1(_06637_),
    .A2(_06688_),
    .A3(_06689_),
    .B1(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__mux2_1 _13945_ (.A0(\rbzero.wall_tracer.stepDistY[-5] ),
    .A1(_06695_),
    .S(_00004_),
    .X(_06696_));
 sky130_fd_sc_hd__clkbuf_1 _13946_ (.A(_06696_),
    .X(_00412_));
 sky130_fd_sc_hd__a21o_1 _13947_ (.A1(_05325_),
    .A2(_06635_),
    .B1(_05271_),
    .X(_06697_));
 sky130_fd_sc_hd__a211o_1 _13948_ (.A1(_06603_),
    .A2(_06633_),
    .B1(_06660_),
    .C1(_05347_),
    .X(_06698_));
 sky130_fd_sc_hd__o21ai_1 _13949_ (.A1(_05324_),
    .A2(_06620_),
    .B1(_06639_),
    .Y(_06699_));
 sky130_fd_sc_hd__or2_1 _13950_ (.A(_05380_),
    .B(_06683_),
    .X(_06700_));
 sky130_fd_sc_hd__o21ai_1 _13951_ (.A1(_05315_),
    .A2(_06699_),
    .B1(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__or2_1 _13952_ (.A(_05310_),
    .B(_06666_),
    .X(_06702_));
 sky130_fd_sc_hd__o21ai_1 _13953_ (.A1(_05376_),
    .A2(_06701_),
    .B1(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__a21o_1 _13954_ (.A1(_05476_),
    .A2(_06703_),
    .B1(_06629_),
    .X(_06704_));
 sky130_fd_sc_hd__a31o_2 _13955_ (.A1(_06637_),
    .A2(_06697_),
    .A3(_06698_),
    .B1(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__mux2_1 _13956_ (.A0(\rbzero.wall_tracer.stepDistY[-4] ),
    .A1(_06705_),
    .S(_00004_),
    .X(_06706_));
 sky130_fd_sc_hd__clkbuf_1 _13957_ (.A(_06706_),
    .X(_00413_));
 sky130_fd_sc_hd__a21o_1 _13958_ (.A1(_05271_),
    .A2(_06604_),
    .B1(_06606_),
    .X(_06707_));
 sky130_fd_sc_hd__a21oi_1 _13959_ (.A1(_06601_),
    .A2(_06572_),
    .B1(_06621_),
    .Y(_06708_));
 sky130_fd_sc_hd__mux2_1 _13960_ (.A0(_06690_),
    .A1(_06708_),
    .S(_06664_),
    .X(_06709_));
 sky130_fd_sc_hd__nor2_1 _13961_ (.A(_06675_),
    .B(_06677_),
    .Y(_06710_));
 sky130_fd_sc_hd__a21oi_2 _13962_ (.A1(_06675_),
    .A2(_06709_),
    .B1(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__a221o_2 _13963_ (.A1(_06707_),
    .A2(_06637_),
    .B1(_06711_),
    .B2(_05476_),
    .C1(_06629_),
    .X(_06712_));
 sky130_fd_sc_hd__mux2_1 _13964_ (.A0(\rbzero.wall_tracer.stepDistY[-3] ),
    .A1(_06712_),
    .S(_00004_),
    .X(_06713_));
 sky130_fd_sc_hd__clkbuf_1 _13965_ (.A(_06713_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _13966_ (.A0(_06572_),
    .A1(_06587_),
    .S(_05349_),
    .X(_06714_));
 sky130_fd_sc_hd__mux4_2 _13967_ (.A0(_06665_),
    .A1(_06683_),
    .A2(_06699_),
    .A3(_06714_),
    .S0(_05380_),
    .S1(_05310_),
    .X(_06715_));
 sky130_fd_sc_hd__a21o_1 _13968_ (.A1(_05476_),
    .A2(_06715_),
    .B1(_05272_),
    .X(_06716_));
 sky130_fd_sc_hd__a31o_4 _13969_ (.A1(_05270_),
    .A2(_06636_),
    .A3(_06637_),
    .B1(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__buf_4 _13970_ (.A(_04836_),
    .X(_06718_));
 sky130_fd_sc_hd__mux2_1 _13971_ (.A0(\rbzero.wall_tracer.stepDistY[-2] ),
    .A1(_06717_),
    .S(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__clkbuf_1 _13972_ (.A(_06719_),
    .X(_00415_));
 sky130_fd_sc_hd__a21o_1 _13973_ (.A1(_05270_),
    .A2(_06652_),
    .B1(_06629_),
    .X(_06720_));
 sky130_fd_sc_hd__inv_2 _13974_ (.A(_06676_),
    .Y(_06721_));
 sky130_fd_sc_hd__and2_1 _13975_ (.A(_06588_),
    .B(_06587_),
    .X(_06722_));
 sky130_fd_sc_hd__a21oi_2 _13976_ (.A1(_06601_),
    .A2(_06600_),
    .B1(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__mux4_1 _13977_ (.A0(_06721_),
    .A1(_06690_),
    .A2(_06708_),
    .A3(_06723_),
    .S0(_06664_),
    .S1(_05310_),
    .X(_06724_));
 sky130_fd_sc_hd__nor2_1 _13978_ (.A(_05390_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__a21o_2 _13979_ (.A1(_05414_),
    .A2(_06720_),
    .B1(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__mux2_1 _13980_ (.A0(\rbzero.wall_tracer.stepDistY[-1] ),
    .A1(_06726_),
    .S(_06718_),
    .X(_06727_));
 sky130_fd_sc_hd__clkbuf_1 _13981_ (.A(_06727_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _13982_ (.A0(_06598_),
    .A1(_06600_),
    .S(_06588_),
    .X(_06728_));
 sky130_fd_sc_hd__or2_1 _13983_ (.A(_05380_),
    .B(_06714_),
    .X(_06729_));
 sky130_fd_sc_hd__o21ai_1 _13984_ (.A1(_05315_),
    .A2(_06728_),
    .B1(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__mux2_1 _13985_ (.A0(_06701_),
    .A1(_06730_),
    .S(_05310_),
    .X(_06731_));
 sky130_fd_sc_hd__a221oi_2 _13986_ (.A1(_05318_),
    .A2(_06663_),
    .B1(_06667_),
    .B2(_05373_),
    .C1(_06629_),
    .Y(_06732_));
 sky130_fd_sc_hd__o21ai_4 _13987_ (.A1(_05390_),
    .A2(_06731_),
    .B1(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__mux2_1 _13988_ (.A0(\rbzero.wall_tracer.stepDistY[0] ),
    .A1(_06733_),
    .S(_06718_),
    .X(_06734_));
 sky130_fd_sc_hd__clkbuf_1 _13989_ (.A(_06734_),
    .X(_00417_));
 sky130_fd_sc_hd__a21oi_1 _13990_ (.A1(_06588_),
    .A2(_06598_),
    .B1(_06605_),
    .Y(_06735_));
 sky130_fd_sc_hd__mux4_2 _13991_ (.A0(_06690_),
    .A1(_06708_),
    .A2(_06723_),
    .A3(_06735_),
    .S0(_06664_),
    .S1(_06675_),
    .X(_06736_));
 sky130_fd_sc_hd__a21oi_1 _13992_ (.A1(_05373_),
    .A2(_06678_),
    .B1(_06629_),
    .Y(_06737_));
 sky130_fd_sc_hd__o221ai_4 _13993_ (.A1(_05320_),
    .A2(_06673_),
    .B1(_06736_),
    .B2(_05390_),
    .C1(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__mux2_1 _13994_ (.A0(\rbzero.wall_tracer.stepDistY[1] ),
    .A1(_06738_),
    .S(_06718_),
    .X(_06739_));
 sky130_fd_sc_hd__clkbuf_1 _13995_ (.A(_06739_),
    .X(_00418_));
 sky130_fd_sc_hd__and2_1 _13996_ (.A(_06675_),
    .B(_06684_),
    .X(_06740_));
 sky130_fd_sc_hd__or2_1 _13997_ (.A(_05380_),
    .B(_06699_),
    .X(_06741_));
 sky130_fd_sc_hd__o21ai_1 _13998_ (.A1(_05315_),
    .A2(_06714_),
    .B1(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__clkinv_2 _13999_ (.A(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__a22o_1 _14000_ (.A1(_06603_),
    .A2(_06634_),
    .B1(_06728_),
    .B2(_05315_),
    .X(_06744_));
 sky130_fd_sc_hd__mux2_1 _14001_ (.A0(_06743_),
    .A1(_06744_),
    .S(_06675_),
    .X(_06745_));
 sky130_fd_sc_hd__a221o_4 _14002_ (.A1(_05373_),
    .A2(_06740_),
    .B1(_06745_),
    .B2(_05476_),
    .C1(_06629_),
    .X(_06746_));
 sky130_fd_sc_hd__mux2_1 _14003_ (.A0(\rbzero.wall_tracer.stepDistY[2] ),
    .A1(_06746_),
    .S(_06718_),
    .X(_06747_));
 sky130_fd_sc_hd__clkbuf_1 _14004_ (.A(_06747_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _14005_ (.A0(_06708_),
    .A1(_06723_),
    .S(_06664_),
    .X(_06748_));
 sky130_fd_sc_hd__nand2_1 _14006_ (.A(_05376_),
    .B(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__a21o_1 _14007_ (.A1(_06588_),
    .A2(_06598_),
    .B1(_06605_),
    .X(_06750_));
 sky130_fd_sc_hd__a21o_1 _14008_ (.A1(_05315_),
    .A2(_06750_),
    .B1(_05376_),
    .X(_06751_));
 sky130_fd_sc_hd__a32o_1 _14009_ (.A1(_05476_),
    .A2(_06749_),
    .A3(_06751_),
    .B1(_05373_),
    .B2(_06693_),
    .X(_06752_));
 sky130_fd_sc_hd__or2_1 _14010_ (.A(_06630_),
    .B(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__mux2_1 _14011_ (.A0(\rbzero.wall_tracer.stepDistY[3] ),
    .A1(_06753_),
    .S(_06718_),
    .X(_06754_));
 sky130_fd_sc_hd__clkbuf_1 _14012_ (.A(_06754_),
    .X(_00420_));
 sky130_fd_sc_hd__nor2_1 _14013_ (.A(_06675_),
    .B(_06730_),
    .Y(_06755_));
 sky130_fd_sc_hd__a21o_1 _14014_ (.A1(_05447_),
    .A2(_06634_),
    .B1(_05322_),
    .X(_06756_));
 sky130_fd_sc_hd__o221a_1 _14015_ (.A1(_05334_),
    .A2(_06703_),
    .B1(_06755_),
    .B2(_06756_),
    .C1(_05369_),
    .X(_06757_));
 sky130_fd_sc_hd__or2_1 _14016_ (.A(_06630_),
    .B(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__buf_2 _14017_ (.A(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__mux2_1 _14018_ (.A0(\rbzero.wall_tracer.stepDistY[4] ),
    .A1(_06759_),
    .S(_06718_),
    .X(_06760_));
 sky130_fd_sc_hd__clkbuf_1 _14019_ (.A(_06760_),
    .X(_00421_));
 sky130_fd_sc_hd__nand2_1 _14020_ (.A(_05315_),
    .B(_06723_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_1 _14021_ (.A(_06664_),
    .B(_06735_),
    .Y(_06762_));
 sky130_fd_sc_hd__nor2_1 _14022_ (.A(_06675_),
    .B(_05390_),
    .Y(_06763_));
 sky130_fd_sc_hd__a32o_2 _14023_ (.A1(_06761_),
    .A2(_06762_),
    .A3(_06763_),
    .B1(_06711_),
    .B2(_05373_),
    .X(_06764_));
 sky130_fd_sc_hd__or2_1 _14024_ (.A(_06630_),
    .B(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__mux2_1 _14025_ (.A0(\rbzero.wall_tracer.stepDistY[5] ),
    .A1(_06765_),
    .S(_06718_),
    .X(_06766_));
 sky130_fd_sc_hd__clkbuf_1 _14026_ (.A(_06766_),
    .X(_00422_));
 sky130_fd_sc_hd__a221o_2 _14027_ (.A1(_05373_),
    .A2(_06715_),
    .B1(_06744_),
    .B2(_06763_),
    .C1(_06630_),
    .X(_06767_));
 sky130_fd_sc_hd__mux2_1 _14028_ (.A0(\rbzero.wall_tracer.stepDistY[6] ),
    .A1(_06767_),
    .S(_06718_),
    .X(_06768_));
 sky130_fd_sc_hd__clkbuf_1 _14029_ (.A(_06768_),
    .X(_00423_));
 sky130_fd_sc_hd__nand2_1 _14030_ (.A(_05322_),
    .B(_06724_),
    .Y(_06769_));
 sky130_fd_sc_hd__a31o_1 _14031_ (.A1(_05315_),
    .A2(_06750_),
    .A3(_06763_),
    .B1(_05373_),
    .X(_06770_));
 sky130_fd_sc_hd__a21oi_4 _14032_ (.A1(_06769_),
    .A2(_06770_),
    .B1(_06630_),
    .Y(_06771_));
 sky130_fd_sc_hd__inv_2 _14033_ (.A(_06771_),
    .Y(_06772_));
 sky130_fd_sc_hd__mux2_1 _14034_ (.A0(\rbzero.wall_tracer.stepDistY[7] ),
    .A1(_06772_),
    .S(_06718_),
    .X(_06773_));
 sky130_fd_sc_hd__clkbuf_1 _14035_ (.A(_06773_),
    .X(_00424_));
 sky130_fd_sc_hd__nor2_2 _14036_ (.A(_06097_),
    .B(_05305_),
    .Y(_06774_));
 sky130_fd_sc_hd__a21oi_1 _14037_ (.A1(_05395_),
    .A2(_06634_),
    .B1(_05373_),
    .Y(_06775_));
 sky130_fd_sc_hd__a221o_1 _14038_ (.A1(_05210_),
    .A2(_05278_),
    .B1(_05322_),
    .B2(_06731_),
    .C1(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__nand2_1 _14039_ (.A(_06774_),
    .B(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__mux2_1 _14040_ (.A0(\rbzero.wall_tracer.stepDistY[8] ),
    .A1(_06777_),
    .S(_04836_),
    .X(_06778_));
 sky130_fd_sc_hd__clkbuf_1 _14041_ (.A(_06778_),
    .X(_00425_));
 sky130_fd_sc_hd__o31ai_4 _14042_ (.A1(_05210_),
    .A2(_05334_),
    .A3(_06736_),
    .B1(_06774_),
    .Y(_06779_));
 sky130_fd_sc_hd__mux2_1 _14043_ (.A0(\rbzero.wall_tracer.stepDistY[9] ),
    .A1(_06779_),
    .S(_04836_),
    .X(_06780_));
 sky130_fd_sc_hd__clkbuf_1 _14044_ (.A(_06780_),
    .X(_00426_));
 sky130_fd_sc_hd__and3_1 _14045_ (.A(_06774_),
    .B(_05373_),
    .C(_06745_),
    .X(_06781_));
 sky130_fd_sc_hd__mux2_1 _14046_ (.A0(\rbzero.wall_tracer.stepDistY[10] ),
    .A1(_06781_),
    .S(_04836_),
    .X(_06782_));
 sky130_fd_sc_hd__clkbuf_1 _14047_ (.A(_06782_),
    .X(_00427_));
 sky130_fd_sc_hd__inv_2 _14048_ (.A(_03495_),
    .Y(_06783_));
 sky130_fd_sc_hd__or2_1 _14049_ (.A(_06783_),
    .B(_05004_),
    .X(_06784_));
 sky130_fd_sc_hd__clkbuf_4 _14050_ (.A(_06784_),
    .X(_06785_));
 sky130_fd_sc_hd__clkbuf_4 _14051_ (.A(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__buf_4 _14052_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_06787_));
 sky130_fd_sc_hd__clkbuf_4 _14053_ (.A(_05005_),
    .X(_06788_));
 sky130_fd_sc_hd__o221a_1 _14054_ (.A1(_06787_),
    .A2(_03496_),
    .B1(_06788_),
    .B2(\rbzero.wall_tracer.trackDistX[-11] ),
    .C1(_03485_),
    .X(_06789_));
 sky130_fd_sc_hd__o21a_1 _14055_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(_06786_),
    .B1(_06789_),
    .X(_00428_));
 sky130_fd_sc_hd__o221a_1 _14056_ (.A1(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A2(_03496_),
    .B1(_06785_),
    .B2(\rbzero.wall_tracer.trackDistY[-10] ),
    .C1(_03485_),
    .X(_06790_));
 sky130_fd_sc_hd__o21a_1 _14057_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(_06788_),
    .B1(_06790_),
    .X(_00429_));
 sky130_fd_sc_hd__clkbuf_4 _14058_ (.A(_05005_),
    .X(_06791_));
 sky130_fd_sc_hd__o221a_1 _14059_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_03496_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-9] ),
    .C1(_03485_),
    .X(_06792_));
 sky130_fd_sc_hd__o21a_1 _14060_ (.A1(\rbzero.wall_tracer.trackDistY[-9] ),
    .A2(_06786_),
    .B1(_06792_),
    .X(_00430_));
 sky130_fd_sc_hd__o221a_1 _14061_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(_03496_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-8] ),
    .C1(_03485_),
    .X(_06793_));
 sky130_fd_sc_hd__o21a_1 _14062_ (.A1(\rbzero.wall_tracer.trackDistY[-8] ),
    .A2(_06786_),
    .B1(_06793_),
    .X(_00431_));
 sky130_fd_sc_hd__o221a_1 _14063_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_03496_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-7] ),
    .C1(_03485_),
    .X(_06794_));
 sky130_fd_sc_hd__o21a_1 _14064_ (.A1(\rbzero.wall_tracer.trackDistY[-7] ),
    .A2(_06786_),
    .B1(_06794_),
    .X(_00432_));
 sky130_fd_sc_hd__o221a_1 _14065_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_03496_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-6] ),
    .C1(_03485_),
    .X(_06795_));
 sky130_fd_sc_hd__o21a_1 _14066_ (.A1(\rbzero.wall_tracer.trackDistY[-6] ),
    .A2(_06786_),
    .B1(_06795_),
    .X(_00433_));
 sky130_fd_sc_hd__clkbuf_4 _14067_ (.A(_03495_),
    .X(_06796_));
 sky130_fd_sc_hd__clkbuf_4 _14068_ (.A(_03484_),
    .X(_06797_));
 sky130_fd_sc_hd__o221a_1 _14069_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_06796_),
    .B1(_06785_),
    .B2(\rbzero.wall_tracer.trackDistY[-5] ),
    .C1(_06797_),
    .X(_06798_));
 sky130_fd_sc_hd__o21a_1 _14070_ (.A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .A2(_06788_),
    .B1(_06798_),
    .X(_00434_));
 sky130_fd_sc_hd__o221a_1 _14071_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_06796_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-4] ),
    .C1(_06797_),
    .X(_06799_));
 sky130_fd_sc_hd__o21a_1 _14072_ (.A1(\rbzero.wall_tracer.trackDistY[-4] ),
    .A2(_06786_),
    .B1(_06799_),
    .X(_00435_));
 sky130_fd_sc_hd__o221a_1 _14073_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_06796_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-3] ),
    .C1(_06797_),
    .X(_06800_));
 sky130_fd_sc_hd__o21a_1 _14074_ (.A1(\rbzero.wall_tracer.trackDistY[-3] ),
    .A2(_06786_),
    .B1(_06800_),
    .X(_00436_));
 sky130_fd_sc_hd__o221a_1 _14075_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_06796_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-2] ),
    .C1(_06797_),
    .X(_06801_));
 sky130_fd_sc_hd__o21a_1 _14076_ (.A1(\rbzero.wall_tracer.trackDistY[-2] ),
    .A2(_06786_),
    .B1(_06801_),
    .X(_00437_));
 sky130_fd_sc_hd__o221a_1 _14077_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_06796_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[-1] ),
    .C1(_06797_),
    .X(_06802_));
 sky130_fd_sc_hd__o21a_1 _14078_ (.A1(\rbzero.wall_tracer.trackDistY[-1] ),
    .A2(_06786_),
    .B1(_06802_),
    .X(_00438_));
 sky130_fd_sc_hd__o221a_1 _14079_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_06796_),
    .B1(_06785_),
    .B2(\rbzero.wall_tracer.trackDistY[0] ),
    .C1(_06797_),
    .X(_06803_));
 sky130_fd_sc_hd__o21a_1 _14080_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(_06788_),
    .B1(_06803_),
    .X(_00439_));
 sky130_fd_sc_hd__o221a_1 _14081_ (.A1(\rbzero.wall_tracer.visualWallDist[1] ),
    .A2(_06796_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[1] ),
    .C1(_06797_),
    .X(_06804_));
 sky130_fd_sc_hd__o21a_1 _14082_ (.A1(\rbzero.wall_tracer.trackDistY[1] ),
    .A2(_06786_),
    .B1(_06804_),
    .X(_00440_));
 sky130_fd_sc_hd__o221a_1 _14083_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_06796_),
    .B1(_06785_),
    .B2(\rbzero.wall_tracer.trackDistY[2] ),
    .C1(_06797_),
    .X(_06805_));
 sky130_fd_sc_hd__o21a_1 _14084_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_06788_),
    .B1(_06805_),
    .X(_00441_));
 sky130_fd_sc_hd__o221a_1 _14085_ (.A1(\rbzero.wall_tracer.visualWallDist[3] ),
    .A2(_06796_),
    .B1(_06785_),
    .B2(\rbzero.wall_tracer.trackDistY[3] ),
    .C1(_06797_),
    .X(_06806_));
 sky130_fd_sc_hd__o21a_1 _14086_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_06788_),
    .B1(_06806_),
    .X(_00442_));
 sky130_fd_sc_hd__o221a_1 _14087_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_06796_),
    .B1(_06785_),
    .B2(\rbzero.wall_tracer.trackDistY[4] ),
    .C1(_06797_),
    .X(_06807_));
 sky130_fd_sc_hd__o21a_1 _14088_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(_06788_),
    .B1(_06807_),
    .X(_00443_));
 sky130_fd_sc_hd__o221a_1 _14089_ (.A1(\rbzero.wall_tracer.visualWallDist[5] ),
    .A2(_03495_),
    .B1(_06785_),
    .B2(\rbzero.wall_tracer.trackDistY[5] ),
    .C1(_03497_),
    .X(_06808_));
 sky130_fd_sc_hd__o21a_1 _14090_ (.A1(\rbzero.wall_tracer.trackDistX[5] ),
    .A2(_06788_),
    .B1(_06808_),
    .X(_00444_));
 sky130_fd_sc_hd__o221a_1 _14091_ (.A1(\rbzero.wall_tracer.visualWallDist[6] ),
    .A2(_03495_),
    .B1(_06784_),
    .B2(\rbzero.wall_tracer.trackDistY[6] ),
    .C1(_03497_),
    .X(_06809_));
 sky130_fd_sc_hd__o21a_1 _14092_ (.A1(\rbzero.wall_tracer.trackDistX[6] ),
    .A2(_06788_),
    .B1(_06809_),
    .X(_00445_));
 sky130_fd_sc_hd__o221a_1 _14093_ (.A1(\rbzero.wall_tracer.visualWallDist[7] ),
    .A2(_03495_),
    .B1(_06791_),
    .B2(\rbzero.wall_tracer.trackDistX[7] ),
    .C1(_03497_),
    .X(_06810_));
 sky130_fd_sc_hd__o21a_1 _14094_ (.A1(\rbzero.wall_tracer.trackDistY[7] ),
    .A2(_06785_),
    .B1(_06810_),
    .X(_00446_));
 sky130_fd_sc_hd__o221a_1 _14095_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_03495_),
    .B1(_05005_),
    .B2(\rbzero.wall_tracer.trackDistX[8] ),
    .C1(_03497_),
    .X(_06811_));
 sky130_fd_sc_hd__o21a_1 _14096_ (.A1(\rbzero.wall_tracer.trackDistY[8] ),
    .A2(_06785_),
    .B1(_06811_),
    .X(_00447_));
 sky130_fd_sc_hd__o21a_1 _14097_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(_04953_),
    .B1(\rbzero.wall_tracer.trackDistY[9] ),
    .X(_06812_));
 sky130_fd_sc_hd__inv_2 _14098_ (.A(_05003_),
    .Y(_06813_));
 sky130_fd_sc_hd__a221o_1 _14099_ (.A1(\rbzero.wall_tracer.trackDistX[9] ),
    .A2(_05004_),
    .B1(_06812_),
    .B2(_06813_),
    .C1(_06783_),
    .X(_06814_));
 sky130_fd_sc_hd__o211a_1 _14100_ (.A1(\rbzero.wall_tracer.visualWallDist[9] ),
    .A2(_03496_),
    .B1(_06814_),
    .C1(_03498_),
    .X(_00448_));
 sky130_fd_sc_hd__a21o_1 _14101_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(\rbzero.wall_tracer.trackDistY[10] ),
    .B1(_06783_),
    .X(_06815_));
 sky130_fd_sc_hd__o211a_1 _14102_ (.A1(\rbzero.wall_tracer.visualWallDist[10] ),
    .A2(_03496_),
    .B1(_06815_),
    .C1(_03498_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14103_ (.A0(\rbzero.wall_tracer.stepDistX[-11] ),
    .A1(_06631_),
    .S(_00008_),
    .X(_06816_));
 sky130_fd_sc_hd__clkbuf_1 _14104_ (.A(_06816_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _14105_ (.A0(\rbzero.wall_tracer.stepDistX[-10] ),
    .A1(_06649_),
    .S(_00008_),
    .X(_06817_));
 sky130_fd_sc_hd__clkbuf_1 _14106_ (.A(_06817_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _14107_ (.A0(\rbzero.wall_tracer.stepDistX[-9] ),
    .A1(_06658_),
    .S(_00008_),
    .X(_06818_));
 sky130_fd_sc_hd__clkbuf_1 _14108_ (.A(_06818_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _14109_ (.A0(\rbzero.wall_tracer.stepDistX[-8] ),
    .A1(_06669_),
    .S(_00008_),
    .X(_06819_));
 sky130_fd_sc_hd__clkbuf_1 _14110_ (.A(_06819_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _14111_ (.A0(\rbzero.wall_tracer.stepDistX[-7] ),
    .A1(_06679_),
    .S(_00008_),
    .X(_06820_));
 sky130_fd_sc_hd__clkbuf_1 _14112_ (.A(_06820_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _14113_ (.A0(\rbzero.wall_tracer.stepDistX[-6] ),
    .A1(_06686_),
    .S(_00008_),
    .X(_06821_));
 sky130_fd_sc_hd__clkbuf_1 _14114_ (.A(_06821_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _14115_ (.A0(\rbzero.wall_tracer.stepDistX[-5] ),
    .A1(_06695_),
    .S(_00008_),
    .X(_06822_));
 sky130_fd_sc_hd__clkbuf_1 _14116_ (.A(_06822_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _14117_ (.A0(\rbzero.wall_tracer.stepDistX[-4] ),
    .A1(_06705_),
    .S(_00008_),
    .X(_06823_));
 sky130_fd_sc_hd__clkbuf_1 _14118_ (.A(_06823_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _14119_ (.A0(\rbzero.wall_tracer.stepDistX[-3] ),
    .A1(_06712_),
    .S(_00008_),
    .X(_06824_));
 sky130_fd_sc_hd__clkbuf_1 _14120_ (.A(_06824_),
    .X(_00458_));
 sky130_fd_sc_hd__buf_4 _14121_ (.A(_04833_),
    .X(_06825_));
 sky130_fd_sc_hd__mux2_1 _14122_ (.A0(\rbzero.wall_tracer.stepDistX[-2] ),
    .A1(_06717_),
    .S(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__clkbuf_1 _14123_ (.A(_06826_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _14124_ (.A0(\rbzero.wall_tracer.stepDistX[-1] ),
    .A1(_06726_),
    .S(_06825_),
    .X(_06827_));
 sky130_fd_sc_hd__clkbuf_1 _14125_ (.A(_06827_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _14126_ (.A0(\rbzero.wall_tracer.stepDistX[0] ),
    .A1(_06733_),
    .S(_06825_),
    .X(_06828_));
 sky130_fd_sc_hd__clkbuf_1 _14127_ (.A(_06828_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _14128_ (.A0(\rbzero.wall_tracer.stepDistX[1] ),
    .A1(_06738_),
    .S(_06825_),
    .X(_06829_));
 sky130_fd_sc_hd__clkbuf_1 _14129_ (.A(_06829_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _14130_ (.A0(\rbzero.wall_tracer.stepDistX[2] ),
    .A1(_06746_),
    .S(_06825_),
    .X(_06830_));
 sky130_fd_sc_hd__clkbuf_1 _14131_ (.A(_06830_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _14132_ (.A0(\rbzero.wall_tracer.stepDistX[3] ),
    .A1(_06753_),
    .S(_06825_),
    .X(_06831_));
 sky130_fd_sc_hd__clkbuf_1 _14133_ (.A(_06831_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _14134_ (.A0(\rbzero.wall_tracer.stepDistX[4] ),
    .A1(_06759_),
    .S(_06825_),
    .X(_06832_));
 sky130_fd_sc_hd__clkbuf_1 _14135_ (.A(_06832_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _14136_ (.A0(\rbzero.wall_tracer.stepDistX[5] ),
    .A1(_06765_),
    .S(_06825_),
    .X(_06833_));
 sky130_fd_sc_hd__clkbuf_1 _14137_ (.A(_06833_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _14138_ (.A0(\rbzero.wall_tracer.stepDistX[6] ),
    .A1(_06767_),
    .S(_06825_),
    .X(_06834_));
 sky130_fd_sc_hd__clkbuf_1 _14139_ (.A(_06834_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _14140_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_06772_),
    .S(_06825_),
    .X(_06835_));
 sky130_fd_sc_hd__clkbuf_1 _14141_ (.A(_06835_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _14142_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_06777_),
    .S(_04833_),
    .X(_06836_));
 sky130_fd_sc_hd__clkbuf_1 _14143_ (.A(_06836_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _14144_ (.A0(\rbzero.wall_tracer.stepDistX[9] ),
    .A1(_06779_),
    .S(_04833_),
    .X(_06837_));
 sky130_fd_sc_hd__clkbuf_1 _14145_ (.A(_06837_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _14146_ (.A0(\rbzero.wall_tracer.stepDistX[10] ),
    .A1(_06781_),
    .S(_04833_),
    .X(_06838_));
 sky130_fd_sc_hd__clkbuf_1 _14147_ (.A(_06838_),
    .X(_00471_));
 sky130_fd_sc_hd__and2_1 _14148_ (.A(_03389_),
    .B(_03454_),
    .X(_06839_));
 sky130_fd_sc_hd__or2b_1 _14149_ (.A(_03455_),
    .B_N(_03389_),
    .X(_06840_));
 sky130_fd_sc_hd__a22o_1 _14150_ (.A1(\rbzero.mapdyw[0] ),
    .A2(_06839_),
    .B1(_06840_),
    .B2(_03409_),
    .X(_06841_));
 sky130_fd_sc_hd__and2_1 _14151_ (.A(_03389_),
    .B(_03429_),
    .X(_06842_));
 sky130_fd_sc_hd__mux2_1 _14152_ (.A0(_06841_),
    .A1(\rbzero.mapdxw[0] ),
    .S(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__mux2_1 _14153_ (.A0(_06843_),
    .A1(\rbzero.wall_tracer.wall[0] ),
    .S(_03458_),
    .X(_06844_));
 sky130_fd_sc_hd__and2_1 _14154_ (.A(_03485_),
    .B(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__clkbuf_1 _14155_ (.A(_06845_),
    .X(_00472_));
 sky130_fd_sc_hd__a22o_1 _14156_ (.A1(\rbzero.mapdyw[1] ),
    .A2(_06839_),
    .B1(_06840_),
    .B2(_03419_),
    .X(_06846_));
 sky130_fd_sc_hd__mux2_1 _14157_ (.A0(_06846_),
    .A1(\rbzero.mapdxw[1] ),
    .S(_06842_),
    .X(_06847_));
 sky130_fd_sc_hd__and3_1 _14158_ (.A(net72),
    .B(\rbzero.wall_tracer.wall[1] ),
    .C(_04827_),
    .X(_06848_));
 sky130_fd_sc_hd__o22a_1 _14159_ (.A1(_03458_),
    .A2(_06847_),
    .B1(_06848_),
    .B2(_00016_),
    .X(_00473_));
 sky130_fd_sc_hd__buf_2 _14160_ (.A(\rbzero.wall_tracer.side ),
    .X(_06849_));
 sky130_fd_sc_hd__clkbuf_4 _14161_ (.A(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__buf_4 _14162_ (.A(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__o211a_1 _14163_ (.A1(_06851_),
    .A2(_03496_),
    .B1(_06788_),
    .C1(_03498_),
    .X(_00474_));
 sky130_fd_sc_hd__clkbuf_4 _14164_ (.A(\rbzero.wall_tracer.state[3] ),
    .X(_06852_));
 sky130_fd_sc_hd__buf_4 _14165_ (.A(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__nor2_2 _14166_ (.A(\rbzero.wall_tracer.state[6] ),
    .B(\rbzero.wall_tracer.state[13] ),
    .Y(_06854_));
 sky130_fd_sc_hd__buf_6 _14167_ (.A(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__nand2_1 _14168_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__buf_2 _14169_ (.A(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__buf_2 _14170_ (.A(_06857_),
    .X(_06858_));
 sky130_fd_sc_hd__inv_2 _14171_ (.A(\rbzero.wall_tracer.state[13] ),
    .Y(_06859_));
 sky130_fd_sc_hd__buf_2 _14172_ (.A(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__mux2_1 _14173_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(_06849_),
    .X(_06861_));
 sky130_fd_sc_hd__a21o_1 _14174_ (.A1(_06852_),
    .A2(_06861_),
    .B1(_03491_),
    .X(_06862_));
 sky130_fd_sc_hd__a21o_1 _14175_ (.A1(_04831_),
    .A2(_06631_),
    .B1(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__o211a_1 _14176_ (.A1(_06860_),
    .A2(\rbzero.wall_tracer.stepDistY[-11] ),
    .B1(_06863_),
    .C1(_04840_),
    .X(_06864_));
 sky130_fd_sc_hd__a21oi_4 _14177_ (.A1(_04949_),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__buf_4 _14178_ (.A(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__a21oi_1 _14179_ (.A1(_03491_),
    .A2(\rbzero.wall_tracer.stepDistY[-10] ),
    .B1(_04948_),
    .Y(_06867_));
 sky130_fd_sc_hd__mux2_1 _14180_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(_06849_),
    .X(_06868_));
 sky130_fd_sc_hd__o21a_1 _14181_ (.A1(_04831_),
    .A2(_06868_),
    .B1(_06859_),
    .X(_06869_));
 sky130_fd_sc_hd__o21ai_1 _14182_ (.A1(_06853_),
    .A2(_06649_),
    .B1(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__a2bb2o_2 _14183_ (.A1_N(_04840_),
    .A2_N(\rbzero.wall_tracer.stepDistX[-10] ),
    .B1(_06867_),
    .B2(_06870_),
    .X(_06871_));
 sky130_fd_sc_hd__clkbuf_4 _14184_ (.A(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__clkbuf_4 _14185_ (.A(_06872_),
    .X(_06873_));
 sky130_fd_sc_hd__nand2_2 _14186_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_06855_),
    .Y(_06874_));
 sky130_fd_sc_hd__buf_2 _14187_ (.A(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__or4_4 _14188_ (.A(_06858_),
    .B(_06866_),
    .C(_06873_),
    .D(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__or3_1 _14189_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(\rbzero.debug_overlay.playerY[-8] ),
    .C(\rbzero.debug_overlay.playerY[-9] ),
    .X(_06877_));
 sky130_fd_sc_hd__o21ai_1 _14190_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(\rbzero.debug_overlay.playerY[-9] ),
    .B1(\rbzero.debug_overlay.playerY[-7] ),
    .Y(_06878_));
 sky130_fd_sc_hd__and2_1 _14191_ (.A(_06877_),
    .B(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__mux2_1 _14192_ (.A0(\rbzero.debug_overlay.playerY[-7] ),
    .A1(_06879_),
    .S(_04927_),
    .X(_06880_));
 sky130_fd_sc_hd__mux2_1 _14193_ (.A0(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A1(_06880_),
    .S(\rbzero.wall_tracer.state[13] ),
    .X(_06881_));
 sky130_fd_sc_hd__or4_1 _14194_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .C(_05113_),
    .D(_05107_),
    .X(_06882_));
 sky130_fd_sc_hd__nor3_1 _14195_ (.A(_05124_),
    .B(_05102_),
    .C(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__and4_1 _14196_ (.A(_05096_),
    .B(_05128_),
    .C(_05091_),
    .D(_06883_),
    .X(_06884_));
 sky130_fd_sc_hd__and4b_1 _14197_ (.A_N(_05137_),
    .B(_05086_),
    .C(_05143_),
    .D(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__a21oi_1 _14198_ (.A1(_05062_),
    .A2(_05060_),
    .B1(_05061_),
    .Y(_06886_));
 sky130_fd_sc_hd__a31o_2 _14199_ (.A1(_05075_),
    .A2(_05064_),
    .A3(_06885_),
    .B1(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__or3_1 _14200_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(\rbzero.debug_overlay.playerX[-8] ),
    .C(\rbzero.debug_overlay.playerX[-9] ),
    .X(_06888_));
 sky130_fd_sc_hd__o21ai_1 _14201_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(\rbzero.debug_overlay.playerX[-9] ),
    .B1(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_06889_));
 sky130_fd_sc_hd__nand2_1 _14202_ (.A(_06888_),
    .B(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__or2_1 _14203_ (.A(_06887_),
    .B(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__a21oi_1 _14204_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_06887_),
    .B1(_04838_),
    .Y(_06892_));
 sky130_fd_sc_hd__a2bb2o_4 _14205_ (.A1_N(_04947_),
    .A2_N(_06881_),
    .B1(_06891_),
    .B2(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__a21oi_1 _14206_ (.A1(_03490_),
    .A2(\rbzero.wall_tracer.stepDistY[-4] ),
    .B1(_04947_),
    .Y(_06894_));
 sky130_fd_sc_hd__clkinv_2 _14207_ (.A(_04904_),
    .Y(_06895_));
 sky130_fd_sc_hd__mux2_1 _14208_ (.A0(_06895_),
    .A1(_05096_),
    .S(\rbzero.wall_tracer.side ),
    .X(_06896_));
 sky130_fd_sc_hd__a21oi_1 _14209_ (.A1(_06852_),
    .A2(_06896_),
    .B1(_03490_),
    .Y(_06897_));
 sky130_fd_sc_hd__o21ai_1 _14210_ (.A1(_06852_),
    .A2(_06705_),
    .B1(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__a2bb2o_2 _14211_ (.A1_N(_04838_),
    .A2_N(\rbzero.wall_tracer.stepDistX[-4] ),
    .B1(_06894_),
    .B2(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__clkbuf_4 _14212_ (.A(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__nor2_1 _14213_ (.A(_06893_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__a21o_1 _14214_ (.A1(_03490_),
    .A2(\rbzero.wall_tracer.stepDistY[-3] ),
    .B1(_04947_),
    .X(_06902_));
 sky130_fd_sc_hd__mux2_1 _14215_ (.A0(_04907_),
    .A1(_05091_),
    .S(\rbzero.wall_tracer.side ),
    .X(_06903_));
 sky130_fd_sc_hd__nand2_1 _14216_ (.A(\rbzero.wall_tracer.state[3] ),
    .B(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__o211a_2 _14217_ (.A1(_06852_),
    .A2(_06712_),
    .B1(_06904_),
    .C1(_06859_),
    .X(_06905_));
 sky130_fd_sc_hd__buf_4 _14218_ (.A(_04947_),
    .X(_06906_));
 sky130_fd_sc_hd__inv_2 _14219_ (.A(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_06907_));
 sky130_fd_sc_hd__a2bb2o_4 _14220_ (.A1_N(_06902_),
    .A2_N(_06905_),
    .B1(_06906_),
    .B2(_06907_),
    .X(_06908_));
 sky130_fd_sc_hd__xor2_1 _14221_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(\rbzero.debug_overlay.playerY[-9] ),
    .X(_06909_));
 sky130_fd_sc_hd__mux2_1 _14222_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(_06909_),
    .S(_04928_),
    .X(_06910_));
 sky130_fd_sc_hd__mux2_1 _14223_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_06910_),
    .S(_03490_),
    .X(_06911_));
 sky130_fd_sc_hd__xnor2_1 _14224_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_06912_));
 sky130_fd_sc_hd__or2_1 _14225_ (.A(_06887_),
    .B(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__buf_4 _14226_ (.A(_06887_),
    .X(_06914_));
 sky130_fd_sc_hd__a21oi_1 _14227_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(_06914_),
    .B1(_04838_),
    .Y(_06915_));
 sky130_fd_sc_hd__a2bb2o_2 _14228_ (.A1_N(_06906_),
    .A2_N(_06911_),
    .B1(_06913_),
    .B2(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__clkbuf_4 _14229_ (.A(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__nor2_1 _14230_ (.A(_06908_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__or2_1 _14231_ (.A(_06893_),
    .B(_06908_),
    .X(_06919_));
 sky130_fd_sc_hd__or3_2 _14232_ (.A(_06919_),
    .B(_06899_),
    .C(_06917_),
    .X(_06920_));
 sky130_fd_sc_hd__o21ai_2 _14233_ (.A1(_06901_),
    .A2(_06918_),
    .B1(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__or2_1 _14234_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_06877_),
    .X(_06922_));
 sky130_fd_sc_hd__nand2_1 _14235_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_06877_),
    .Y(_06923_));
 sky130_fd_sc_hd__and2_1 _14236_ (.A(_06922_),
    .B(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__mux2_1 _14237_ (.A0(\rbzero.debug_overlay.playerY[-6] ),
    .A1(_06924_),
    .S(_04928_),
    .X(_06925_));
 sky130_fd_sc_hd__mux2_1 _14238_ (.A0(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A1(_06925_),
    .S(_03491_),
    .X(_06926_));
 sky130_fd_sc_hd__or2_1 _14239_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_06888_),
    .X(_06927_));
 sky130_fd_sc_hd__nand2_1 _14240_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_06888_),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _14241_ (.A(_06927_),
    .B(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__or2_1 _14242_ (.A(_06914_),
    .B(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__a21oi_1 _14243_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_06914_),
    .B1(_04839_),
    .Y(_06931_));
 sky130_fd_sc_hd__a2bb2o_2 _14244_ (.A1_N(_04948_),
    .A2_N(_06926_),
    .B1(_06930_),
    .B2(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__clkbuf_4 _14245_ (.A(_06932_),
    .X(_06933_));
 sky130_fd_sc_hd__a21o_1 _14246_ (.A1(_03490_),
    .A2(\rbzero.wall_tracer.stepDistY[-5] ),
    .B1(\rbzero.wall_tracer.state[6] ),
    .X(_06934_));
 sky130_fd_sc_hd__mux2_1 _14247_ (.A0(_04901_),
    .A1(_05128_),
    .S(\rbzero.wall_tracer.side ),
    .X(_06935_));
 sky130_fd_sc_hd__nand2_1 _14248_ (.A(\rbzero.wall_tracer.state[3] ),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__o211a_1 _14249_ (.A1(_06852_),
    .A2(_06695_),
    .B1(_06936_),
    .C1(_06859_),
    .X(_06937_));
 sky130_fd_sc_hd__o22ai_4 _14250_ (.A1(_04838_),
    .A2(\rbzero.wall_tracer.stepDistX[-5] ),
    .B1(_06934_),
    .B2(_06937_),
    .Y(_06938_));
 sky130_fd_sc_hd__buf_2 _14251_ (.A(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__clkbuf_4 _14252_ (.A(_06939_),
    .X(_06940_));
 sky130_fd_sc_hd__o31ai_4 _14253_ (.A1(_06921_),
    .A2(_06933_),
    .A3(_06940_),
    .B1(_06920_),
    .Y(_06941_));
 sky130_fd_sc_hd__inv_2 _14254_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .Y(_06942_));
 sky130_fd_sc_hd__xnor2_1 _14255_ (.A(_06942_),
    .B(_06922_),
    .Y(_06943_));
 sky130_fd_sc_hd__mux2_1 _14256_ (.A0(\rbzero.debug_overlay.playerY[-5] ),
    .A1(_06943_),
    .S(_04927_),
    .X(_06944_));
 sky130_fd_sc_hd__mux2_1 _14257_ (.A0(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A1(_06944_),
    .S(\rbzero.wall_tracer.state[13] ),
    .X(_06945_));
 sky130_fd_sc_hd__xnor2_1 _14258_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_06927_),
    .Y(_06946_));
 sky130_fd_sc_hd__or2_1 _14259_ (.A(_06887_),
    .B(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__a21oi_1 _14260_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_06887_),
    .B1(_04838_),
    .Y(_06948_));
 sky130_fd_sc_hd__a2bb2o_4 _14261_ (.A1_N(_04947_),
    .A2_N(_06945_),
    .B1(_06947_),
    .B2(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__a21o_1 _14262_ (.A1(\rbzero.wall_tracer.state[13] ),
    .A2(\rbzero.wall_tracer.stepDistY[-6] ),
    .B1(\rbzero.wall_tracer.state[6] ),
    .X(_06950_));
 sky130_fd_sc_hd__nor2_1 _14263_ (.A(\rbzero.wall_tracer.side ),
    .B(_04894_),
    .Y(_06951_));
 sky130_fd_sc_hd__a211o_1 _14264_ (.A1(_06849_),
    .A2(_05102_),
    .B1(_06951_),
    .C1(_04830_),
    .X(_06952_));
 sky130_fd_sc_hd__o311a_1 _14265_ (.A1(\rbzero.wall_tracer.state[3] ),
    .A2(_06682_),
    .A3(_06685_),
    .B1(_06952_),
    .C1(_06859_),
    .X(_06953_));
 sky130_fd_sc_hd__o22ai_4 _14266_ (.A1(_04838_),
    .A2(\rbzero.wall_tracer.stepDistX[-6] ),
    .B1(_06950_),
    .B2(_06953_),
    .Y(_06954_));
 sky130_fd_sc_hd__or2_1 _14267_ (.A(_06949_),
    .B(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__or3_1 _14268_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .C(_06922_),
    .X(_06956_));
 sky130_fd_sc_hd__o21ai_1 _14269_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_06922_),
    .B1(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_06957_));
 sky130_fd_sc_hd__and2_1 _14270_ (.A(_06956_),
    .B(_06957_),
    .X(_06958_));
 sky130_fd_sc_hd__mux2_1 _14271_ (.A0(\rbzero.debug_overlay.playerY[-4] ),
    .A1(_06958_),
    .S(_04927_),
    .X(_06959_));
 sky130_fd_sc_hd__mux2_1 _14272_ (.A0(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A1(_06959_),
    .S(\rbzero.wall_tracer.state[13] ),
    .X(_06960_));
 sky130_fd_sc_hd__or3_1 _14273_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(\rbzero.debug_overlay.playerX[-5] ),
    .C(_06927_),
    .X(_06961_));
 sky130_fd_sc_hd__o21ai_1 _14274_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_06927_),
    .B1(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_06962_));
 sky130_fd_sc_hd__nand2_1 _14275_ (.A(_06961_),
    .B(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__or2_1 _14276_ (.A(_06887_),
    .B(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__a21oi_1 _14277_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_06887_),
    .B1(_04838_),
    .Y(_06965_));
 sky130_fd_sc_hd__a2bb2o_4 _14278_ (.A1_N(_04947_),
    .A2_N(_06960_),
    .B1(_06964_),
    .B2(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__or3_1 _14279_ (.A(_06940_),
    .B(_06955_),
    .C(_06966_),
    .X(_06967_));
 sky130_fd_sc_hd__clkbuf_4 _14280_ (.A(_06949_),
    .X(_06968_));
 sky130_fd_sc_hd__buf_4 _14281_ (.A(_06954_),
    .X(_06969_));
 sky130_fd_sc_hd__clkbuf_4 _14282_ (.A(_06966_),
    .X(_06970_));
 sky130_fd_sc_hd__o22ai_1 _14283_ (.A1(_06940_),
    .A2(_06968_),
    .B1(_06969_),
    .B2(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__nand2_1 _14284_ (.A(_06967_),
    .B(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__a21oi_1 _14285_ (.A1(_03490_),
    .A2(\rbzero.wall_tracer.stepDistY[-7] ),
    .B1(_04947_),
    .Y(_06973_));
 sky130_fd_sc_hd__mux2_1 _14286_ (.A0(_04890_),
    .A1(_05124_),
    .S(\rbzero.wall_tracer.side ),
    .X(_06974_));
 sky130_fd_sc_hd__o21a_1 _14287_ (.A1(_04830_),
    .A2(_06974_),
    .B1(_06859_),
    .X(_06975_));
 sky130_fd_sc_hd__o21ai_1 _14288_ (.A1(_06852_),
    .A2(_06679_),
    .B1(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__a2bb2o_4 _14289_ (.A1_N(_04838_),
    .A2_N(\rbzero.wall_tracer.stepDistX[-7] ),
    .B1(_06973_),
    .B2(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__clkbuf_4 _14290_ (.A(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__clkbuf_4 _14291_ (.A(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__or2_1 _14292_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_06956_),
    .X(_06980_));
 sky130_fd_sc_hd__nand2_1 _14293_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_06956_),
    .Y(_06981_));
 sky130_fd_sc_hd__and2_1 _14294_ (.A(_06980_),
    .B(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__mux2_1 _14295_ (.A0(\rbzero.debug_overlay.playerY[-3] ),
    .A1(_06982_),
    .S(_04928_),
    .X(_06983_));
 sky130_fd_sc_hd__nand2_1 _14296_ (.A(_03491_),
    .B(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__clkbuf_4 _14297_ (.A(_06859_),
    .X(_06985_));
 sky130_fd_sc_hd__a21oi_1 _14298_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_06985_),
    .B1(_06906_),
    .Y(_06986_));
 sky130_fd_sc_hd__or2_1 _14299_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_06961_),
    .X(_06987_));
 sky130_fd_sc_hd__nand2_1 _14300_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_06961_),
    .Y(_06988_));
 sky130_fd_sc_hd__nand2_1 _14301_ (.A(_06987_),
    .B(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__inv_2 _14302_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .Y(_06990_));
 sky130_fd_sc_hd__mux2_1 _14303_ (.A0(_06989_),
    .A1(_06990_),
    .S(_06914_),
    .X(_06991_));
 sky130_fd_sc_hd__a22o_1 _14304_ (.A1(_06984_),
    .A2(_06986_),
    .B1(_06991_),
    .B2(_04948_),
    .X(_06992_));
 sky130_fd_sc_hd__buf_4 _14305_ (.A(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__nor2_1 _14306_ (.A(_06979_),
    .B(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__xnor2_1 _14307_ (.A(_06972_),
    .B(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__xnor2_1 _14308_ (.A(_06941_),
    .B(_06995_),
    .Y(_06996_));
 sky130_fd_sc_hd__buf_4 _14309_ (.A(_06993_),
    .X(_06997_));
 sky130_fd_sc_hd__or2_1 _14310_ (.A(_06966_),
    .B(_06977_),
    .X(_06998_));
 sky130_fd_sc_hd__or4_1 _14311_ (.A(_06949_),
    .B(_06954_),
    .C(_06966_),
    .D(_06977_),
    .X(_06999_));
 sky130_fd_sc_hd__a21bo_1 _14312_ (.A1(_06955_),
    .A2(_06998_),
    .B1_N(_06999_),
    .X(_07000_));
 sky130_fd_sc_hd__a21oi_1 _14313_ (.A1(_03491_),
    .A2(\rbzero.wall_tracer.stepDistY[-8] ),
    .B1(_06906_),
    .Y(_07001_));
 sky130_fd_sc_hd__nor2_1 _14314_ (.A(_06849_),
    .B(_04898_),
    .Y(_07002_));
 sky130_fd_sc_hd__a211o_1 _14315_ (.A1(_06850_),
    .A2(_05107_),
    .B1(_07002_),
    .C1(_04830_),
    .X(_07003_));
 sky130_fd_sc_hd__o211ai_1 _14316_ (.A1(_06852_),
    .A2(_06669_),
    .B1(_07003_),
    .C1(_06985_),
    .Y(_07004_));
 sky130_fd_sc_hd__a2bb2o_4 _14317_ (.A1_N(_04839_),
    .A2_N(\rbzero.wall_tracer.stepDistX[-8] ),
    .B1(_07001_),
    .B2(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__buf_2 _14318_ (.A(_07005_),
    .X(_07006_));
 sky130_fd_sc_hd__clkbuf_4 _14319_ (.A(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__o31ai_2 _14320_ (.A1(_06997_),
    .A2(_07000_),
    .A3(_07007_),
    .B1(_06999_),
    .Y(_07008_));
 sky130_fd_sc_hd__or2b_1 _14321_ (.A(_06996_),
    .B_N(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__a21bo_1 _14322_ (.A1(_06941_),
    .A2(_06995_),
    .B1_N(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__clkbuf_4 _14323_ (.A(_06866_),
    .X(_07011_));
 sky130_fd_sc_hd__clkbuf_4 _14324_ (.A(_06875_),
    .X(_07012_));
 sky130_fd_sc_hd__or2_1 _14325_ (.A(_06856_),
    .B(_06872_),
    .X(_07013_));
 sky130_fd_sc_hd__o21ai_2 _14326_ (.A1(_07011_),
    .A2(_07012_),
    .B1(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__nand2_1 _14327_ (.A(_06876_),
    .B(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__inv_2 _14328_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .Y(_07016_));
 sky130_fd_sc_hd__xnor2_1 _14329_ (.A(_07016_),
    .B(_06980_),
    .Y(_07017_));
 sky130_fd_sc_hd__mux2_1 _14330_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(_07017_),
    .S(_04928_),
    .X(_07018_));
 sky130_fd_sc_hd__nand2_1 _14331_ (.A(_03492_),
    .B(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__a21oi_1 _14332_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_06985_),
    .B1(_06906_),
    .Y(_07020_));
 sky130_fd_sc_hd__xnor2_1 _14333_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_06987_),
    .Y(_07021_));
 sky130_fd_sc_hd__inv_2 _14334_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .Y(_07022_));
 sky130_fd_sc_hd__mux2_1 _14335_ (.A0(_07021_),
    .A1(_07022_),
    .S(_06914_),
    .X(_07023_));
 sky130_fd_sc_hd__a22o_4 _14336_ (.A1(_07019_),
    .A2(_07020_),
    .B1(_07023_),
    .B2(_04948_),
    .X(_07024_));
 sky130_fd_sc_hd__or2_1 _14337_ (.A(_06978_),
    .B(_07024_),
    .X(_07025_));
 sky130_fd_sc_hd__or3_4 _14338_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .C(_06980_),
    .X(_07026_));
 sky130_fd_sc_hd__o21ai_1 _14339_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_06980_),
    .B1(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_07027_));
 sky130_fd_sc_hd__nand2_1 _14340_ (.A(_07026_),
    .B(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__nor2_1 _14341_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(_04928_),
    .Y(_07029_));
 sky130_fd_sc_hd__a21oi_1 _14342_ (.A1(_04928_),
    .A2(_07028_),
    .B1(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__mux2_1 _14343_ (.A0(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A1(_07030_),
    .S(_03490_),
    .X(_07031_));
 sky130_fd_sc_hd__or3_4 _14344_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .B(\rbzero.debug_overlay.playerX[-2] ),
    .C(_06987_),
    .X(_07032_));
 sky130_fd_sc_hd__o21ai_1 _14345_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_06987_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_07033_));
 sky130_fd_sc_hd__and2_1 _14346_ (.A(_07032_),
    .B(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__mux2_1 _14347_ (.A0(_07034_),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_06887_),
    .X(_07035_));
 sky130_fd_sc_hd__or2_1 _14348_ (.A(_04839_),
    .B(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__o21ai_4 _14349_ (.A1(_04948_),
    .A2(_07031_),
    .B1(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__or2_1 _14350_ (.A(_07005_),
    .B(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__buf_2 _14351_ (.A(_07024_),
    .X(_07039_));
 sky130_fd_sc_hd__or2_1 _14352_ (.A(_06978_),
    .B(_07037_),
    .X(_07040_));
 sky130_fd_sc_hd__or3_1 _14353_ (.A(_07006_),
    .B(_07039_),
    .C(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__a21bo_1 _14354_ (.A1(_07025_),
    .A2(_07038_),
    .B1_N(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__a21oi_1 _14355_ (.A1(_03491_),
    .A2(\rbzero.wall_tracer.stepDistY[-9] ),
    .B1(_06906_),
    .Y(_07043_));
 sky130_fd_sc_hd__nor2_1 _14356_ (.A(_06849_),
    .B(_04896_),
    .Y(_07044_));
 sky130_fd_sc_hd__a211o_1 _14357_ (.A1(_06850_),
    .A2(_05113_),
    .B1(_07044_),
    .C1(_04830_),
    .X(_07045_));
 sky130_fd_sc_hd__o211ai_1 _14358_ (.A1(_06852_),
    .A2(_06658_),
    .B1(_07045_),
    .C1(_06985_),
    .Y(_07046_));
 sky130_fd_sc_hd__a2bb2o_2 _14359_ (.A1_N(_04839_),
    .A2_N(\rbzero.wall_tracer.stepDistX[-9] ),
    .B1(_07043_),
    .B2(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__buf_2 _14360_ (.A(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__clkbuf_4 _14361_ (.A(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__or3_1 _14362_ (.A(_06985_),
    .B(_04922_),
    .C(_07026_),
    .X(_07050_));
 sky130_fd_sc_hd__o2bb2a_1 _14363_ (.A1_N(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2_N(_06855_),
    .B1(_07050_),
    .B2(_04948_),
    .X(_07051_));
 sky130_fd_sc_hd__o31a_4 _14364_ (.A1(_04840_),
    .A2(_06914_),
    .A3(_07032_),
    .B1(_07051_),
    .X(_07052_));
 sky130_fd_sc_hd__nor2_1 _14365_ (.A(_07049_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__xor2_1 _14366_ (.A(_07042_),
    .B(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__nor2_1 _14367_ (.A(_06871_),
    .B(_07052_),
    .Y(_07055_));
 sky130_fd_sc_hd__nor3_1 _14368_ (.A(_07024_),
    .B(_07038_),
    .C(_07047_),
    .Y(_07056_));
 sky130_fd_sc_hd__o22a_1 _14369_ (.A1(_07005_),
    .A2(_07024_),
    .B1(_07037_),
    .B2(_07047_),
    .X(_07057_));
 sky130_fd_sc_hd__nor2_1 _14370_ (.A(_07056_),
    .B(_07057_),
    .Y(_07058_));
 sky130_fd_sc_hd__a21oi_1 _14371_ (.A1(_07055_),
    .A2(_07058_),
    .B1(_07056_),
    .Y(_07059_));
 sky130_fd_sc_hd__nor2_1 _14372_ (.A(_07054_),
    .B(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_1 _14373_ (.A(_07054_),
    .B(_07059_),
    .Y(_07061_));
 sky130_fd_sc_hd__and2b_1 _14374_ (.A_N(_07060_),
    .B(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__xnor2_1 _14375_ (.A(_07015_),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__xnor2_1 _14376_ (.A(_07010_),
    .B(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__xnor2_1 _14377_ (.A(_07055_),
    .B(_07058_),
    .Y(_07065_));
 sky130_fd_sc_hd__or2_1 _14378_ (.A(_06865_),
    .B(_07052_),
    .X(_07066_));
 sky130_fd_sc_hd__o22a_1 _14379_ (.A1(_06871_),
    .A2(_07037_),
    .B1(_07048_),
    .B2(_07024_),
    .X(_07067_));
 sky130_fd_sc_hd__or4_1 _14380_ (.A(_06871_),
    .B(_07024_),
    .C(_07037_),
    .D(_07047_),
    .X(_07068_));
 sky130_fd_sc_hd__o21a_1 _14381_ (.A1(_07066_),
    .A2(_07067_),
    .B1(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__nor2_2 _14382_ (.A(_06857_),
    .B(_06866_),
    .Y(_07070_));
 sky130_fd_sc_hd__xor2_1 _14383_ (.A(_07065_),
    .B(_07069_),
    .X(_07071_));
 sky130_fd_sc_hd__nand2_1 _14384_ (.A(_07070_),
    .B(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__o21ai_1 _14385_ (.A1(_07065_),
    .A2(_07069_),
    .B1(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__and2b_1 _14386_ (.A_N(_07064_),
    .B(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__a21oi_1 _14387_ (.A1(_07010_),
    .A2(_07063_),
    .B1(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__nor2_2 _14388_ (.A(_06876_),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__nor2_1 _14389_ (.A(_06900_),
    .B(_06970_),
    .Y(_07077_));
 sky130_fd_sc_hd__clkbuf_4 _14390_ (.A(_06908_),
    .X(_07078_));
 sky130_fd_sc_hd__nor2_1 _14391_ (.A(_07078_),
    .B(_06968_),
    .Y(_07079_));
 sky130_fd_sc_hd__nor2_1 _14392_ (.A(_07078_),
    .B(_06970_),
    .Y(_07080_));
 sky130_fd_sc_hd__nor2_1 _14393_ (.A(_06900_),
    .B(_06968_),
    .Y(_07081_));
 sky130_fd_sc_hd__nand2_1 _14394_ (.A(_07080_),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__o21a_1 _14395_ (.A1(_07077_),
    .A2(_07079_),
    .B1(_07082_),
    .X(_07083_));
 sky130_fd_sc_hd__buf_2 _14396_ (.A(_06940_),
    .X(_07084_));
 sky130_fd_sc_hd__nor2_1 _14397_ (.A(_07084_),
    .B(_06993_),
    .Y(_07085_));
 sky130_fd_sc_hd__a21bo_1 _14398_ (.A1(_07083_),
    .A2(_07085_),
    .B1_N(_07082_),
    .X(_07086_));
 sky130_fd_sc_hd__o21ai_1 _14399_ (.A1(_06859_),
    .A2(\rbzero.wall_tracer.stepDistY[-2] ),
    .B1(_04838_),
    .Y(_07087_));
 sky130_fd_sc_hd__mux2_1 _14400_ (.A0(_04911_),
    .A1(_05086_),
    .S(\rbzero.wall_tracer.side ),
    .X(_07088_));
 sky130_fd_sc_hd__or2_1 _14401_ (.A(_04830_),
    .B(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__o211a_1 _14402_ (.A1(\rbzero.wall_tracer.state[3] ),
    .A2(_06717_),
    .B1(_07089_),
    .C1(_06859_),
    .X(_07090_));
 sky130_fd_sc_hd__o2bb2a_2 _14403_ (.A1_N(_04947_),
    .A2_N(\rbzero.wall_tracer.stepDistX[-2] ),
    .B1(_07087_),
    .B2(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__clkbuf_4 _14404_ (.A(_07091_),
    .X(_07092_));
 sky130_fd_sc_hd__nor2_1 _14405_ (.A(_06968_),
    .B(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__or2_1 _14406_ (.A(_06966_),
    .B(_07092_),
    .X(_07094_));
 sky130_fd_sc_hd__or3_1 _14407_ (.A(_07078_),
    .B(_06968_),
    .C(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__o21a_1 _14408_ (.A1(_07080_),
    .A2(_07093_),
    .B1(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__clkbuf_4 _14409_ (.A(_06900_),
    .X(_07097_));
 sky130_fd_sc_hd__nor2_1 _14410_ (.A(_07097_),
    .B(_06993_),
    .Y(_07098_));
 sky130_fd_sc_hd__xnor2_1 _14411_ (.A(_07096_),
    .B(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__clkbuf_4 _14412_ (.A(_06933_),
    .X(_07100_));
 sky130_fd_sc_hd__buf_2 _14413_ (.A(_06917_),
    .X(_07101_));
 sky130_fd_sc_hd__inv_2 _14414_ (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_07102_));
 sky130_fd_sc_hd__a211o_2 _14415_ (.A1(_05414_),
    .A2(_06720_),
    .B1(_06725_),
    .C1(_06717_),
    .X(_07103_));
 sky130_fd_sc_hd__xnor2_1 _14416_ (.A(_06733_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__nand2_1 _14417_ (.A(_06849_),
    .B(_05137_),
    .Y(_07105_));
 sky130_fd_sc_hd__o211a_1 _14418_ (.A1(_06849_),
    .A2(_04915_),
    .B1(_07105_),
    .C1(\rbzero.wall_tracer.state[3] ),
    .X(_07106_));
 sky130_fd_sc_hd__a211o_2 _14419_ (.A1(_04830_),
    .A2(_07104_),
    .B1(_07106_),
    .C1(_03490_),
    .X(_07107_));
 sky130_fd_sc_hd__a21oi_1 _14420_ (.A1(_03492_),
    .A2(\rbzero.wall_tracer.stepDistY[0] ),
    .B1(_04949_),
    .Y(_07108_));
 sky130_fd_sc_hd__a22o_1 _14421_ (.A1(_04949_),
    .A2(_07102_),
    .B1(_07107_),
    .B2(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__or2_1 _14422_ (.A(_07101_),
    .B(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__xnor2_1 _14423_ (.A(_06717_),
    .B(_06726_),
    .Y(_07111_));
 sky130_fd_sc_hd__or2_1 _14424_ (.A(_06849_),
    .B(_04888_),
    .X(_07112_));
 sky130_fd_sc_hd__a21oi_1 _14425_ (.A1(_06850_),
    .A2(_05143_),
    .B1(_04830_),
    .Y(_07113_));
 sky130_fd_sc_hd__a221o_2 _14426_ (.A1(_04831_),
    .A2(_07111_),
    .B1(_07112_),
    .B2(_07113_),
    .C1(_03490_),
    .X(_07114_));
 sky130_fd_sc_hd__inv_2 _14427_ (.A(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_07115_));
 sky130_fd_sc_hd__a21oi_1 _14428_ (.A1(_03491_),
    .A2(_07115_),
    .B1(_06906_),
    .Y(_07116_));
 sky130_fd_sc_hd__a22oi_4 _14429_ (.A1(_06906_),
    .A2(\rbzero.wall_tracer.stepDistX[-1] ),
    .B1(_07114_),
    .B2(_07116_),
    .Y(_07117_));
 sky130_fd_sc_hd__or2_1 _14430_ (.A(_06893_),
    .B(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__buf_2 _14431_ (.A(_06893_),
    .X(_07119_));
 sky130_fd_sc_hd__or2_1 _14432_ (.A(_07101_),
    .B(_07117_),
    .X(_07120_));
 sky130_fd_sc_hd__or3_1 _14433_ (.A(_07119_),
    .B(_07109_),
    .C(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__a21bo_1 _14434_ (.A1(_07110_),
    .A2(_07118_),
    .B1_N(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__clkbuf_4 _14435_ (.A(_07092_),
    .X(_07123_));
 sky130_fd_sc_hd__o31ai_1 _14436_ (.A1(_07100_),
    .A2(_07122_),
    .A3(_07123_),
    .B1(_07121_),
    .Y(_07124_));
 sky130_fd_sc_hd__or2b_1 _14437_ (.A(_07099_),
    .B_N(_07124_),
    .X(_07125_));
 sky130_fd_sc_hd__or2b_1 _14438_ (.A(_07124_),
    .B_N(_07099_),
    .X(_07126_));
 sky130_fd_sc_hd__nand2_1 _14439_ (.A(_07125_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__xnor2_1 _14440_ (.A(_07086_),
    .B(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand3_1 _14441_ (.A(_06733_),
    .B(_06738_),
    .C(_07103_),
    .Y(_07129_));
 sky130_fd_sc_hd__a21o_1 _14442_ (.A1(_06733_),
    .A2(_07103_),
    .B1(_06738_),
    .X(_07130_));
 sky130_fd_sc_hd__nand2_1 _14443_ (.A(_07129_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__mux2_1 _14444_ (.A0(_04920_),
    .A1(_05075_),
    .S(_06850_),
    .X(_07132_));
 sky130_fd_sc_hd__o21ai_1 _14445_ (.A1(_04831_),
    .A2(_07132_),
    .B1(_06985_),
    .Y(_07133_));
 sky130_fd_sc_hd__a21oi_2 _14446_ (.A1(_04831_),
    .A2(_07131_),
    .B1(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__o21ai_1 _14447_ (.A1(_06860_),
    .A2(\rbzero.wall_tracer.stepDistY[1] ),
    .B1(_04840_),
    .Y(_07135_));
 sky130_fd_sc_hd__o2bb2a_2 _14448_ (.A1_N(_04949_),
    .A2_N(\rbzero.wall_tracer.stepDistX[1] ),
    .B1(_07134_),
    .B2(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__clkbuf_4 _14449_ (.A(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__buf_2 _14450_ (.A(_07109_),
    .X(_07138_));
 sky130_fd_sc_hd__o22ai_1 _14451_ (.A1(_07119_),
    .A2(_07138_),
    .B1(_07137_),
    .B2(_07101_),
    .Y(_07139_));
 sky130_fd_sc_hd__o31a_1 _14452_ (.A1(_07119_),
    .A2(_07110_),
    .A3(_07137_),
    .B1(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__buf_4 _14453_ (.A(_07117_),
    .X(_07141_));
 sky130_fd_sc_hd__nor2_1 _14454_ (.A(_07100_),
    .B(_07141_),
    .Y(_07142_));
 sky130_fd_sc_hd__xor2_1 _14455_ (.A(_07140_),
    .B(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__nor2_1 _14456_ (.A(_04947_),
    .B(_06859_),
    .Y(_07144_));
 sky130_fd_sc_hd__clkinv_2 _14457_ (.A(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_07145_));
 sky130_fd_sc_hd__nor2_1 _14458_ (.A(_07145_),
    .B(_04839_),
    .Y(_07146_));
 sky130_fd_sc_hd__a221oi_4 _14459_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_06855_),
    .B1(_07144_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .C1(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__clkbuf_4 _14460_ (.A(_07147_),
    .X(_07148_));
 sky130_fd_sc_hd__xnor2_1 _14461_ (.A(_06746_),
    .B(_07130_),
    .Y(_07149_));
 sky130_fd_sc_hd__nand2_1 _14462_ (.A(_06850_),
    .B(_05064_),
    .Y(_07150_));
 sky130_fd_sc_hd__o211a_1 _14463_ (.A1(_06850_),
    .A2(_04886_),
    .B1(_07150_),
    .C1(_06853_),
    .X(_07151_));
 sky130_fd_sc_hd__a211o_2 _14464_ (.A1(_04831_),
    .A2(_07149_),
    .B1(_07151_),
    .C1(_03492_),
    .X(_07152_));
 sky130_fd_sc_hd__o21a_1 _14465_ (.A1(_06860_),
    .A2(\rbzero.wall_tracer.stepDistY[2] ),
    .B1(_04840_),
    .X(_07153_));
 sky130_fd_sc_hd__a22oi_4 _14466_ (.A1(_04949_),
    .A2(\rbzero.wall_tracer.stepDistX[2] ),
    .B1(_07152_),
    .B2(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__or2_1 _14467_ (.A(_07148_),
    .B(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__nand2_2 _14468_ (.A(_06787_),
    .B(_06855_),
    .Y(_07156_));
 sky130_fd_sc_hd__clkbuf_4 _14469_ (.A(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__nor2_1 _14470_ (.A(_04840_),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_07158_));
 sky130_fd_sc_hd__inv_2 _14471_ (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_07159_));
 sky130_fd_sc_hd__mux2_1 _14472_ (.A0(_04881_),
    .A1(_05171_),
    .S(_06849_),
    .X(_07160_));
 sky130_fd_sc_hd__a21oi_4 _14473_ (.A1(_06852_),
    .A2(_07160_),
    .B1(_03491_),
    .Y(_07161_));
 sky130_fd_sc_hd__inv_2 _14474_ (.A(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__nor2_1 _14475_ (.A(_06630_),
    .B(_06752_),
    .Y(_07163_));
 sky130_fd_sc_hd__a211oi_1 _14476_ (.A1(_06733_),
    .A2(_07103_),
    .B1(_06746_),
    .C1(_06738_),
    .Y(_07164_));
 sky130_fd_sc_hd__a2111o_2 _14477_ (.A1(_06733_),
    .A2(_07103_),
    .B1(_06752_),
    .C1(_06746_),
    .D1(_06738_),
    .X(_07165_));
 sky130_fd_sc_hd__o211a_1 _14478_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07165_),
    .C1(_04831_),
    .X(_07166_));
 sky130_fd_sc_hd__o221a_1 _14479_ (.A1(_06860_),
    .A2(_07159_),
    .B1(_07162_),
    .B2(_07166_),
    .C1(_04840_),
    .X(_07167_));
 sky130_fd_sc_hd__nor3_2 _14480_ (.A(_07157_),
    .B(_07158_),
    .C(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__or2_1 _14481_ (.A(_06759_),
    .B(_07165_),
    .X(_07169_));
 sky130_fd_sc_hd__nand2_1 _14482_ (.A(_06759_),
    .B(_07165_),
    .Y(_07170_));
 sky130_fd_sc_hd__a31o_1 _14483_ (.A1(_04831_),
    .A2(_07169_),
    .A3(_07170_),
    .B1(_07162_),
    .X(_07171_));
 sky130_fd_sc_hd__a21oi_1 _14484_ (.A1(_03492_),
    .A2(\rbzero.wall_tracer.stepDistY[4] ),
    .B1(_04949_),
    .Y(_07172_));
 sky130_fd_sc_hd__o2bb2a_4 _14485_ (.A1_N(_07171_),
    .A2_N(_07172_),
    .B1(_04841_),
    .B2(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_07173_));
 sky130_fd_sc_hd__and2_2 _14486_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_06855_),
    .X(_07174_));
 sky130_fd_sc_hd__inv_2 _14487_ (.A(_06787_),
    .Y(_07175_));
 sky130_fd_sc_hd__or4_2 _14488_ (.A(_07175_),
    .B(_04949_),
    .C(_03492_),
    .D(_07171_),
    .X(_07176_));
 sky130_fd_sc_hd__nand2_2 _14489_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_06854_),
    .Y(_07177_));
 sky130_fd_sc_hd__buf_2 _14490_ (.A(_07177_),
    .X(_07178_));
 sky130_fd_sc_hd__or3_2 _14491_ (.A(_07158_),
    .B(_07167_),
    .C(_07178_),
    .X(_07179_));
 sky130_fd_sc_hd__a32oi_4 _14492_ (.A1(_07168_),
    .A2(_07173_),
    .A3(_07174_),
    .B1(_07176_),
    .B2(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__xnor2_1 _14493_ (.A(_07155_),
    .B(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__nor2_1 _14494_ (.A(_07136_),
    .B(_07148_),
    .Y(_07182_));
 sky130_fd_sc_hd__and4_1 _14495_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_04841_),
    .C(_06860_),
    .D(_07152_),
    .X(_07183_));
 sky130_fd_sc_hd__o32a_1 _14496_ (.A1(_07154_),
    .A2(_07157_),
    .A3(_07179_),
    .B1(_07183_),
    .B2(_07168_),
    .X(_07184_));
 sky130_fd_sc_hd__clkbuf_4 _14497_ (.A(_07157_),
    .X(_07185_));
 sky130_fd_sc_hd__or3_1 _14498_ (.A(_07154_),
    .B(_07185_),
    .C(_07179_),
    .X(_07186_));
 sky130_fd_sc_hd__a21boi_1 _14499_ (.A1(_07182_),
    .A2(_07184_),
    .B1_N(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__xnor2_1 _14500_ (.A(_07181_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__xnor2_1 _14501_ (.A(_07143_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__nor2_1 _14502_ (.A(_07100_),
    .B(_07123_),
    .Y(_07190_));
 sky130_fd_sc_hd__xnor2_1 _14503_ (.A(_07122_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__xnor2_1 _14504_ (.A(_07182_),
    .B(_07184_),
    .Y(_07192_));
 sky130_fd_sc_hd__or2_1 _14505_ (.A(_07109_),
    .B(_07148_),
    .X(_07193_));
 sky130_fd_sc_hd__and4_1 _14506_ (.A(_06787_),
    .B(_04840_),
    .C(_06860_),
    .D(_07152_),
    .X(_07194_));
 sky130_fd_sc_hd__inv_2 _14507_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .Y(_07195_));
 sky130_fd_sc_hd__nor4_2 _14508_ (.A(_07195_),
    .B(_04948_),
    .C(_03492_),
    .D(_07134_),
    .Y(_07196_));
 sky130_fd_sc_hd__nor2_1 _14509_ (.A(_07194_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__clkbuf_4 _14510_ (.A(_07154_),
    .X(_07198_));
 sky130_fd_sc_hd__clkbuf_4 _14511_ (.A(_07178_),
    .X(_07199_));
 sky130_fd_sc_hd__or4_1 _14512_ (.A(_07175_),
    .B(_04948_),
    .C(_03492_),
    .D(_07134_),
    .X(_07200_));
 sky130_fd_sc_hd__or3_1 _14513_ (.A(_07198_),
    .B(_07199_),
    .C(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__o21a_1 _14514_ (.A1(_07193_),
    .A2(_07197_),
    .B1(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__xor2_1 _14515_ (.A(_07192_),
    .B(_07202_),
    .X(_07203_));
 sky130_fd_sc_hd__nor2_1 _14516_ (.A(_07192_),
    .B(_07202_),
    .Y(_07204_));
 sky130_fd_sc_hd__a21oi_1 _14517_ (.A1(_07191_),
    .A2(_07203_),
    .B1(_07204_),
    .Y(_07205_));
 sky130_fd_sc_hd__nor2_1 _14518_ (.A(_07189_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand2_1 _14519_ (.A(_07189_),
    .B(_07205_),
    .Y(_07207_));
 sky130_fd_sc_hd__and2b_1 _14520_ (.A_N(_07206_),
    .B(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__xnor2_1 _14521_ (.A(_07128_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__xnor2_1 _14522_ (.A(_07191_),
    .B(_07203_),
    .Y(_07210_));
 sky130_fd_sc_hd__o32a_1 _14523_ (.A1(_07154_),
    .A2(_07178_),
    .A3(_07200_),
    .B1(_07196_),
    .B2(_07194_),
    .X(_07211_));
 sky130_fd_sc_hd__xnor2_1 _14524_ (.A(_07193_),
    .B(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__clkbuf_4 _14525_ (.A(_07148_),
    .X(_07213_));
 sky130_fd_sc_hd__and4bb_1 _14526_ (.A_N(_06906_),
    .B_N(_07107_),
    .C(_06985_),
    .D(_06787_),
    .X(_07214_));
 sky130_fd_sc_hd__or4_1 _14527_ (.A(_07195_),
    .B(_06906_),
    .C(_03491_),
    .D(_07107_),
    .X(_07215_));
 sky130_fd_sc_hd__a22o_1 _14528_ (.A1(_07196_),
    .A2(_07214_),
    .B1(_07215_),
    .B2(_07200_),
    .X(_07216_));
 sky130_fd_sc_hd__nand2_1 _14529_ (.A(_07196_),
    .B(_07214_),
    .Y(_07217_));
 sky130_fd_sc_hd__o31a_1 _14530_ (.A1(_07141_),
    .A2(_07213_),
    .A3(_07216_),
    .B1(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__xnor2_1 _14531_ (.A(_07212_),
    .B(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__or2_1 _14532_ (.A(_06893_),
    .B(_07092_),
    .X(_07220_));
 sky130_fd_sc_hd__nand2_1 _14533_ (.A(_07120_),
    .B(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__or2_1 _14534_ (.A(_06917_),
    .B(_07092_),
    .X(_07222_));
 sky130_fd_sc_hd__or2_1 _14535_ (.A(_07118_),
    .B(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__or4bb_1 _14536_ (.A(_07078_),
    .B(_06933_),
    .C_N(_07221_),
    .D_N(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__a2bb2o_1 _14537_ (.A1_N(_07078_),
    .A2_N(_06933_),
    .B1(_07221_),
    .B2(_07223_),
    .X(_07225_));
 sky130_fd_sc_hd__and2_1 _14538_ (.A(_07224_),
    .B(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__or2b_1 _14539_ (.A(_07218_),
    .B_N(_07212_),
    .X(_07227_));
 sky130_fd_sc_hd__a21boi_1 _14540_ (.A1(_07219_),
    .A2(_07226_),
    .B1_N(_07227_),
    .Y(_07228_));
 sky130_fd_sc_hd__nor2_1 _14541_ (.A(_07210_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__and2_1 _14542_ (.A(_07210_),
    .B(_07228_),
    .X(_07230_));
 sky130_fd_sc_hd__nor2_1 _14543_ (.A(_07229_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__nor2_1 _14544_ (.A(_06940_),
    .B(_06970_),
    .Y(_07232_));
 sky130_fd_sc_hd__or4_1 _14545_ (.A(_06900_),
    .B(_06940_),
    .C(_06968_),
    .D(_06970_),
    .X(_07233_));
 sky130_fd_sc_hd__o21a_1 _14546_ (.A1(_07232_),
    .A2(_07081_),
    .B1(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__clkbuf_4 _14547_ (.A(_06969_),
    .X(_07235_));
 sky130_fd_sc_hd__nor2_1 _14548_ (.A(_07235_),
    .B(_06993_),
    .Y(_07236_));
 sky130_fd_sc_hd__a21boi_1 _14549_ (.A1(_07234_),
    .A2(_07236_),
    .B1_N(_07233_),
    .Y(_07237_));
 sky130_fd_sc_hd__xnor2_1 _14550_ (.A(_07083_),
    .B(_07085_),
    .Y(_07238_));
 sky130_fd_sc_hd__a21o_1 _14551_ (.A1(_07223_),
    .A2(_07224_),
    .B1(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__nand3_1 _14552_ (.A(_07223_),
    .B(_07224_),
    .C(_07238_),
    .Y(_07240_));
 sky130_fd_sc_hd__and2_1 _14553_ (.A(_07239_),
    .B(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__xnor2_1 _14554_ (.A(_07237_),
    .B(_07241_),
    .Y(_07242_));
 sky130_fd_sc_hd__a21oi_1 _14555_ (.A1(_07231_),
    .A2(_07242_),
    .B1(_07229_),
    .Y(_07243_));
 sky130_fd_sc_hd__nor2_1 _14556_ (.A(_07209_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__and2_1 _14557_ (.A(_07209_),
    .B(_07243_),
    .X(_07245_));
 sky130_fd_sc_hd__nor2_1 _14558_ (.A(_07244_),
    .B(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__or2_1 _14559_ (.A(_06969_),
    .B(_07024_),
    .X(_07247_));
 sky130_fd_sc_hd__or3_1 _14560_ (.A(_07235_),
    .B(_07037_),
    .C(_07025_),
    .X(_07248_));
 sky130_fd_sc_hd__a21bo_1 _14561_ (.A1(_07040_),
    .A2(_07247_),
    .B1_N(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__or2_1 _14562_ (.A(_07007_),
    .B(_07052_),
    .X(_07250_));
 sky130_fd_sc_hd__xnor2_1 _14563_ (.A(_07249_),
    .B(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__o31a_1 _14564_ (.A1(_07042_),
    .A2(_07049_),
    .A3(_07052_),
    .B1(_07041_),
    .X(_07252_));
 sky130_fd_sc_hd__or3_1 _14565_ (.A(_06874_),
    .B(_07013_),
    .C(_07049_),
    .X(_07253_));
 sky130_fd_sc_hd__o22ai_1 _14566_ (.A1(_06873_),
    .A2(_06875_),
    .B1(_07049_),
    .B2(_06857_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand2_1 _14567_ (.A(_07253_),
    .B(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__clkbuf_8 _14568_ (.A(_06855_),
    .X(_07256_));
 sky130_fd_sc_hd__nand2_1 _14569_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__nor2_1 _14570_ (.A(_06866_),
    .B(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__xnor2_1 _14571_ (.A(_07255_),
    .B(_07258_),
    .Y(_07259_));
 sky130_fd_sc_hd__xor2_1 _14572_ (.A(_07251_),
    .B(_07252_),
    .X(_07260_));
 sky130_fd_sc_hd__nand2_1 _14573_ (.A(_07259_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__o21ai_2 _14574_ (.A1(_07251_),
    .A2(_07252_),
    .B1(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__or2b_1 _14575_ (.A(_07237_),
    .B_N(_07241_),
    .X(_07263_));
 sky130_fd_sc_hd__or4_1 _14576_ (.A(_06857_),
    .B(_06875_),
    .C(_07007_),
    .D(_07049_),
    .X(_07264_));
 sky130_fd_sc_hd__clkbuf_4 _14577_ (.A(_07049_),
    .X(_07265_));
 sky130_fd_sc_hd__nor2_1 _14578_ (.A(_06857_),
    .B(_07007_),
    .Y(_07266_));
 sky130_fd_sc_hd__o21bai_1 _14579_ (.A1(_07012_),
    .A2(_07265_),
    .B1_N(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__nand2_1 _14580_ (.A(_07264_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__buf_2 _14581_ (.A(_06873_),
    .X(_07269_));
 sky130_fd_sc_hd__buf_2 _14582_ (.A(_07257_),
    .X(_07270_));
 sky130_fd_sc_hd__nor2_1 _14583_ (.A(_07269_),
    .B(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__xnor2_1 _14584_ (.A(_07268_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__buf_4 _14585_ (.A(_07037_),
    .X(_07273_));
 sky130_fd_sc_hd__or3_1 _14586_ (.A(_06940_),
    .B(_07273_),
    .C(_07247_),
    .X(_07274_));
 sky130_fd_sc_hd__o22a_1 _14587_ (.A1(_06940_),
    .A2(_07024_),
    .B1(_07037_),
    .B2(_06969_),
    .X(_07275_));
 sky130_fd_sc_hd__inv_2 _14588_ (.A(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__nor2_1 _14589_ (.A(_06979_),
    .B(_07052_),
    .Y(_07277_));
 sky130_fd_sc_hd__and3_1 _14590_ (.A(_07274_),
    .B(_07276_),
    .C(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__a21oi_1 _14591_ (.A1(_07274_),
    .A2(_07276_),
    .B1(_07277_),
    .Y(_07279_));
 sky130_fd_sc_hd__or2_1 _14592_ (.A(_07278_),
    .B(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__clkbuf_4 _14593_ (.A(_07052_),
    .X(_07281_));
 sky130_fd_sc_hd__o31a_1 _14594_ (.A1(_07007_),
    .A2(_07281_),
    .A3(_07249_),
    .B1(_07248_),
    .X(_07282_));
 sky130_fd_sc_hd__nor2_1 _14595_ (.A(_07280_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__and2_1 _14596_ (.A(_07280_),
    .B(_07282_),
    .X(_07284_));
 sky130_fd_sc_hd__nor2_1 _14597_ (.A(_07283_),
    .B(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__xnor2_1 _14598_ (.A(_07272_),
    .B(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__a21o_1 _14599_ (.A1(_07239_),
    .A2(_07263_),
    .B1(_07286_),
    .X(_07287_));
 sky130_fd_sc_hd__nand3_1 _14600_ (.A(_07239_),
    .B(_07263_),
    .C(_07286_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand2_1 _14601_ (.A(_07287_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__xnor2_1 _14602_ (.A(_07262_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__xnor2_2 _14603_ (.A(_07246_),
    .B(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__xnor2_1 _14604_ (.A(_07231_),
    .B(_07242_),
    .Y(_07292_));
 sky130_fd_sc_hd__xnor2_1 _14605_ (.A(_07219_),
    .B(_07226_),
    .Y(_07293_));
 sky130_fd_sc_hd__nor2_1 _14606_ (.A(_07141_),
    .B(_07148_),
    .Y(_07294_));
 sky130_fd_sc_hd__xnor2_1 _14607_ (.A(_07216_),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__and4_1 _14608_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_04839_),
    .C(_06985_),
    .D(_07114_),
    .X(_07296_));
 sky130_fd_sc_hd__o32a_1 _14609_ (.A1(_07117_),
    .A2(_07156_),
    .A3(_07215_),
    .B1(_07296_),
    .B2(_07214_),
    .X(_07297_));
 sky130_fd_sc_hd__nor2_1 _14610_ (.A(_07092_),
    .B(_07147_),
    .Y(_07298_));
 sky130_fd_sc_hd__nand2_1 _14611_ (.A(_07297_),
    .B(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__o31a_1 _14612_ (.A1(_07141_),
    .A2(_07157_),
    .A3(_07215_),
    .B1(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__xnor2_1 _14613_ (.A(_07295_),
    .B(_07300_),
    .Y(_07301_));
 sky130_fd_sc_hd__or3_1 _14614_ (.A(_06908_),
    .B(_06917_),
    .C(_07220_),
    .X(_07302_));
 sky130_fd_sc_hd__a21bo_1 _14615_ (.A1(_06919_),
    .A2(_07222_),
    .B1_N(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__nor2_1 _14616_ (.A(_06900_),
    .B(_06933_),
    .Y(_07304_));
 sky130_fd_sc_hd__xnor2_1 _14617_ (.A(_07303_),
    .B(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__or2b_1 _14618_ (.A(_07300_),
    .B_N(_07295_),
    .X(_07306_));
 sky130_fd_sc_hd__a21bo_1 _14619_ (.A1(_07301_),
    .A2(_07305_),
    .B1_N(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__xnor2_1 _14620_ (.A(_07293_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__a21bo_1 _14621_ (.A1(_06971_),
    .A2(_06994_),
    .B1_N(_06967_),
    .X(_07309_));
 sky130_fd_sc_hd__or3_1 _14622_ (.A(_07097_),
    .B(_07100_),
    .C(_07303_),
    .X(_07310_));
 sky130_fd_sc_hd__xnor2_1 _14623_ (.A(_07234_),
    .B(_07236_),
    .Y(_07311_));
 sky130_fd_sc_hd__a21o_1 _14624_ (.A1(_07302_),
    .A2(_07310_),
    .B1(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__nand3_1 _14625_ (.A(_07302_),
    .B(_07310_),
    .C(_07311_),
    .Y(_07313_));
 sky130_fd_sc_hd__nand2_1 _14626_ (.A(_07312_),
    .B(_07313_),
    .Y(_07314_));
 sky130_fd_sc_hd__xnor2_1 _14627_ (.A(_07309_),
    .B(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__and2b_1 _14628_ (.A_N(_07293_),
    .B(_07307_),
    .X(_07316_));
 sky130_fd_sc_hd__a21oi_1 _14629_ (.A1(_07308_),
    .A2(_07315_),
    .B1(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__xor2_1 _14630_ (.A(_07292_),
    .B(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__a31o_1 _14631_ (.A1(_06876_),
    .A2(_07014_),
    .A3(_07061_),
    .B1(_07060_),
    .X(_07319_));
 sky130_fd_sc_hd__or2b_1 _14632_ (.A(_07314_),
    .B_N(_07309_),
    .X(_07320_));
 sky130_fd_sc_hd__or2_1 _14633_ (.A(_07259_),
    .B(_07260_),
    .X(_07321_));
 sky130_fd_sc_hd__nand2_1 _14634_ (.A(_07261_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__a21o_1 _14635_ (.A1(_07312_),
    .A2(_07320_),
    .B1(_07322_),
    .X(_07323_));
 sky130_fd_sc_hd__nand3_1 _14636_ (.A(_07312_),
    .B(_07320_),
    .C(_07322_),
    .Y(_07324_));
 sky130_fd_sc_hd__nand2_1 _14637_ (.A(_07323_),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__xnor2_1 _14638_ (.A(_07319_),
    .B(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__nor2_1 _14639_ (.A(_07292_),
    .B(_07317_),
    .Y(_07327_));
 sky130_fd_sc_hd__a21oi_2 _14640_ (.A1(_07318_),
    .A2(_07326_),
    .B1(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__xor2_2 _14641_ (.A(_07291_),
    .B(_07328_),
    .X(_07329_));
 sky130_fd_sc_hd__or2b_1 _14642_ (.A(_07325_),
    .B_N(_07319_),
    .X(_07330_));
 sky130_fd_sc_hd__a21bo_1 _14643_ (.A1(_07254_),
    .A2(_07258_),
    .B1_N(_07253_),
    .X(_07331_));
 sky130_fd_sc_hd__nand2_2 _14644_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_06855_),
    .Y(_07332_));
 sky130_fd_sc_hd__clkbuf_4 _14645_ (.A(_07332_),
    .X(_07333_));
 sky130_fd_sc_hd__nor2_1 _14646_ (.A(_07011_),
    .B(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__xnor2_2 _14647_ (.A(_07331_),
    .B(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__a21oi_4 _14648_ (.A1(_07323_),
    .A2(_07330_),
    .B1(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__and3_1 _14649_ (.A(_07323_),
    .B(_07330_),
    .C(_07335_),
    .X(_07337_));
 sky130_fd_sc_hd__nor2_2 _14650_ (.A(_07336_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__xnor2_1 _14651_ (.A(_07329_),
    .B(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__xnor2_1 _14652_ (.A(_07318_),
    .B(_07326_),
    .Y(_07340_));
 sky130_fd_sc_hd__xnor2_1 _14653_ (.A(_07308_),
    .B(_07315_),
    .Y(_07341_));
 sky130_fd_sc_hd__xnor2_1 _14654_ (.A(_07301_),
    .B(_07305_),
    .Y(_07342_));
 sky130_fd_sc_hd__xnor2_1 _14655_ (.A(_07297_),
    .B(_07298_),
    .Y(_07343_));
 sky130_fd_sc_hd__nor2_1 _14656_ (.A(_07091_),
    .B(_07156_),
    .Y(_07344_));
 sky130_fd_sc_hd__or2_1 _14657_ (.A(_06908_),
    .B(_07147_),
    .X(_07345_));
 sky130_fd_sc_hd__and4_1 _14658_ (.A(_06787_),
    .B(_04839_),
    .C(_06860_),
    .D(_07114_),
    .X(_07346_));
 sky130_fd_sc_hd__nor2_1 _14659_ (.A(_07091_),
    .B(_07177_),
    .Y(_07347_));
 sky130_fd_sc_hd__nor2_1 _14660_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__o2bb2a_1 _14661_ (.A1_N(_07296_),
    .A2_N(_07344_),
    .B1(_07345_),
    .B2(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__xor2_1 _14662_ (.A(_07343_),
    .B(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__nor2_1 _14663_ (.A(_06933_),
    .B(_06939_),
    .Y(_07351_));
 sky130_fd_sc_hd__xnor2_1 _14664_ (.A(_06921_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__nor2_1 _14665_ (.A(_07343_),
    .B(_07349_),
    .Y(_07353_));
 sky130_fd_sc_hd__a21oi_2 _14666_ (.A1(_07350_),
    .A2(_07352_),
    .B1(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__xor2_1 _14667_ (.A(_07342_),
    .B(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__xnor2_1 _14668_ (.A(_07008_),
    .B(_06996_),
    .Y(_07356_));
 sky130_fd_sc_hd__nor2_1 _14669_ (.A(_07342_),
    .B(_07354_),
    .Y(_07357_));
 sky130_fd_sc_hd__a21oi_1 _14670_ (.A1(_07355_),
    .A2(_07356_),
    .B1(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__nand2_1 _14671_ (.A(_07341_),
    .B(_07358_),
    .Y(_07359_));
 sky130_fd_sc_hd__xnor2_1 _14672_ (.A(_07073_),
    .B(_07064_),
    .Y(_07360_));
 sky130_fd_sc_hd__nor2_1 _14673_ (.A(_07341_),
    .B(_07358_),
    .Y(_07361_));
 sky130_fd_sc_hd__a21oi_1 _14674_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__nor2_1 _14675_ (.A(_07340_),
    .B(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__and2_1 _14676_ (.A(_07340_),
    .B(_07362_),
    .X(_07364_));
 sky130_fd_sc_hd__nor2_1 _14677_ (.A(_07363_),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__and2_1 _14678_ (.A(_06876_),
    .B(_07075_),
    .X(_07366_));
 sky130_fd_sc_hd__nor2_1 _14679_ (.A(_07076_),
    .B(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__a21oi_1 _14680_ (.A1(_07365_),
    .A2(_07367_),
    .B1(_07363_),
    .Y(_07368_));
 sky130_fd_sc_hd__nor2_1 _14681_ (.A(_07339_),
    .B(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__and2_1 _14682_ (.A(_07339_),
    .B(_07368_),
    .X(_07370_));
 sky130_fd_sc_hd__nor2_2 _14683_ (.A(_07369_),
    .B(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__xnor2_4 _14684_ (.A(_07076_),
    .B(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__and2b_1 _14685_ (.A_N(_07361_),
    .B(_07359_),
    .X(_07373_));
 sky130_fd_sc_hd__xnor2_1 _14686_ (.A(_07373_),
    .B(_07360_),
    .Y(_07374_));
 sky130_fd_sc_hd__xnor2_1 _14687_ (.A(_07355_),
    .B(_07356_),
    .Y(_07375_));
 sky130_fd_sc_hd__xnor2_1 _14688_ (.A(_07350_),
    .B(_07352_),
    .Y(_07376_));
 sky130_fd_sc_hd__nor2_1 _14689_ (.A(_06932_),
    .B(_06969_),
    .Y(_07377_));
 sky130_fd_sc_hd__nor2_1 _14690_ (.A(_06917_),
    .B(_06939_),
    .Y(_07378_));
 sky130_fd_sc_hd__o22ai_1 _14691_ (.A1(_06900_),
    .A2(_06917_),
    .B1(_06939_),
    .B2(_06893_),
    .Y(_07379_));
 sky130_fd_sc_hd__a21bo_1 _14692_ (.A1(_06901_),
    .A2(_07378_),
    .B1_N(_07379_),
    .X(_07380_));
 sky130_fd_sc_hd__xnor2_1 _14693_ (.A(_07377_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__o2bb2a_1 _14694_ (.A1_N(_07296_),
    .A2_N(_07344_),
    .B1(_07347_),
    .B2(_07346_),
    .X(_07382_));
 sky130_fd_sc_hd__xnor2_1 _14695_ (.A(_07345_),
    .B(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__and4_1 _14696_ (.A(_06787_),
    .B(_04839_),
    .C(_06985_),
    .D(_06905_),
    .X(_07384_));
 sky130_fd_sc_hd__nor2_1 _14697_ (.A(_06900_),
    .B(_07147_),
    .Y(_07385_));
 sky130_fd_sc_hd__and4_1 _14698_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_04839_),
    .C(_06985_),
    .D(_06905_),
    .X(_07386_));
 sky130_fd_sc_hd__o2bb2a_1 _14699_ (.A1_N(_07347_),
    .A2_N(_07384_),
    .B1(_07386_),
    .B2(_07344_),
    .X(_07387_));
 sky130_fd_sc_hd__nand2_1 _14700_ (.A(_07385_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__a21boi_1 _14701_ (.A1(_07347_),
    .A2(_07384_),
    .B1_N(_07388_),
    .Y(_07389_));
 sky130_fd_sc_hd__xnor2_1 _14702_ (.A(_07383_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__or2b_1 _14703_ (.A(_07389_),
    .B_N(_07383_),
    .X(_07391_));
 sky130_fd_sc_hd__a21bo_1 _14704_ (.A1(_07381_),
    .A2(_07390_),
    .B1_N(_07391_),
    .X(_07392_));
 sky130_fd_sc_hd__xnor2_1 _14705_ (.A(_07376_),
    .B(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__or2_1 _14706_ (.A(_06949_),
    .B(_07005_),
    .X(_07394_));
 sky130_fd_sc_hd__or2_1 _14707_ (.A(_06998_),
    .B(_07394_),
    .X(_07395_));
 sky130_fd_sc_hd__nor2_1 _14708_ (.A(_06993_),
    .B(_07048_),
    .Y(_07396_));
 sky130_fd_sc_hd__o22a_1 _14709_ (.A1(_06949_),
    .A2(_06977_),
    .B1(_07005_),
    .B2(_06966_),
    .X(_07397_));
 sky130_fd_sc_hd__o21ba_1 _14710_ (.A1(_06998_),
    .A2(_07394_),
    .B1_N(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__nand2_1 _14711_ (.A(_07396_),
    .B(_07398_),
    .Y(_07399_));
 sky130_fd_sc_hd__a22o_1 _14712_ (.A1(_07377_),
    .A2(_07379_),
    .B1(_07378_),
    .B2(_06901_),
    .X(_07400_));
 sky130_fd_sc_hd__nor2_1 _14713_ (.A(_06993_),
    .B(_07005_),
    .Y(_07401_));
 sky130_fd_sc_hd__xnor2_1 _14714_ (.A(_07000_),
    .B(_07401_),
    .Y(_07402_));
 sky130_fd_sc_hd__xnor2_1 _14715_ (.A(_07400_),
    .B(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__a21o_1 _14716_ (.A1(_07395_),
    .A2(_07399_),
    .B1(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__nand3_1 _14717_ (.A(_07395_),
    .B(_07399_),
    .C(_07403_),
    .Y(_07405_));
 sky130_fd_sc_hd__and2_1 _14718_ (.A(_07404_),
    .B(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__or2b_1 _14719_ (.A(_07376_),
    .B_N(_07392_),
    .X(_07407_));
 sky130_fd_sc_hd__a21boi_2 _14720_ (.A1(_07393_),
    .A2(_07406_),
    .B1_N(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__xor2_1 _14721_ (.A(_07375_),
    .B(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__or2_1 _14722_ (.A(_06865_),
    .B(_07039_),
    .X(_07410_));
 sky130_fd_sc_hd__nor3_1 _14723_ (.A(_06872_),
    .B(_07273_),
    .C(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__inv_2 _14724_ (.A(_07068_),
    .Y(_07412_));
 sky130_fd_sc_hd__nor2_1 _14725_ (.A(_07412_),
    .B(_07067_),
    .Y(_07413_));
 sky130_fd_sc_hd__xnor2_1 _14726_ (.A(_07066_),
    .B(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__nand2_1 _14727_ (.A(_07411_),
    .B(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__nand2_1 _14728_ (.A(_07400_),
    .B(_07402_),
    .Y(_07416_));
 sky130_fd_sc_hd__or2_1 _14729_ (.A(_07070_),
    .B(_07071_),
    .X(_07417_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(_07072_),
    .B(_07417_),
    .Y(_07418_));
 sky130_fd_sc_hd__a21oi_1 _14731_ (.A1(_07416_),
    .A2(_07404_),
    .B1(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__and3_1 _14732_ (.A(_07416_),
    .B(_07404_),
    .C(_07418_),
    .X(_07420_));
 sky130_fd_sc_hd__nor2_1 _14733_ (.A(_07419_),
    .B(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__xnor2_1 _14734_ (.A(_07415_),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__nor2_1 _14735_ (.A(_07375_),
    .B(_07408_),
    .Y(_07423_));
 sky130_fd_sc_hd__a21oi_2 _14736_ (.A1(_07409_),
    .A2(_07422_),
    .B1(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__xnor2_2 _14737_ (.A(_07374_),
    .B(_07424_),
    .Y(_07425_));
 sky130_fd_sc_hd__o21ba_1 _14738_ (.A1(_07415_),
    .A2(_07420_),
    .B1_N(_07419_),
    .X(_07426_));
 sky130_fd_sc_hd__xnor2_2 _14739_ (.A(_07425_),
    .B(_07426_),
    .Y(_07427_));
 sky130_fd_sc_hd__xnor2_1 _14740_ (.A(_07396_),
    .B(_07398_),
    .Y(_07428_));
 sky130_fd_sc_hd__or2_1 _14741_ (.A(_06932_),
    .B(_06978_),
    .X(_07429_));
 sky130_fd_sc_hd__o22a_1 _14742_ (.A1(_06917_),
    .A2(_06939_),
    .B1(_06969_),
    .B2(_06893_),
    .X(_07430_));
 sky130_fd_sc_hd__or4_1 _14743_ (.A(_06893_),
    .B(_06916_),
    .C(_06939_),
    .D(_06954_),
    .X(_07431_));
 sky130_fd_sc_hd__o21ai_1 _14744_ (.A1(_07429_),
    .A2(_07430_),
    .B1(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__or2b_1 _14745_ (.A(_07428_),
    .B_N(_07432_),
    .X(_07433_));
 sky130_fd_sc_hd__nor2_1 _14746_ (.A(_06871_),
    .B(_06993_),
    .Y(_07434_));
 sky130_fd_sc_hd__or2_1 _14747_ (.A(_06966_),
    .B(_07047_),
    .X(_07435_));
 sky130_fd_sc_hd__nor4_1 _14748_ (.A(_06949_),
    .B(_06966_),
    .C(_07005_),
    .D(_07047_),
    .Y(_07436_));
 sky130_fd_sc_hd__a21oi_1 _14749_ (.A1(_07394_),
    .A2(_07435_),
    .B1(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__a21oi_1 _14750_ (.A1(_07434_),
    .A2(_07437_),
    .B1(_07436_),
    .Y(_07438_));
 sky130_fd_sc_hd__xnor2_1 _14751_ (.A(_07432_),
    .B(_07428_),
    .Y(_07439_));
 sky130_fd_sc_hd__or2b_1 _14752_ (.A(_07438_),
    .B_N(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__or2_1 _14753_ (.A(_07411_),
    .B(_07414_),
    .X(_07441_));
 sky130_fd_sc_hd__nand2_1 _14754_ (.A(_07415_),
    .B(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__a21oi_2 _14755_ (.A1(_07433_),
    .A2(_07440_),
    .B1(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__xnor2_1 _14756_ (.A(_07409_),
    .B(_07422_),
    .Y(_07444_));
 sky130_fd_sc_hd__xnor2_1 _14757_ (.A(_07393_),
    .B(_07406_),
    .Y(_07445_));
 sky130_fd_sc_hd__xnor2_1 _14758_ (.A(_07438_),
    .B(_07439_),
    .Y(_07446_));
 sky130_fd_sc_hd__xnor2_1 _14759_ (.A(_07381_),
    .B(_07390_),
    .Y(_07447_));
 sky130_fd_sc_hd__xnor2_1 _14760_ (.A(_07385_),
    .B(_07387_),
    .Y(_07448_));
 sky130_fd_sc_hd__nor2_1 _14761_ (.A(_06939_),
    .B(_07147_),
    .Y(_07449_));
 sky130_fd_sc_hd__or2_1 _14762_ (.A(_06899_),
    .B(_07156_),
    .X(_07450_));
 sky130_fd_sc_hd__nor2_1 _14763_ (.A(_06899_),
    .B(_07177_),
    .Y(_07451_));
 sky130_fd_sc_hd__o32a_1 _14764_ (.A1(_06908_),
    .A2(_07177_),
    .A3(_07450_),
    .B1(_07451_),
    .B2(_07384_),
    .X(_07452_));
 sky130_fd_sc_hd__nor3_1 _14765_ (.A(_07078_),
    .B(_07178_),
    .C(_07450_),
    .Y(_07453_));
 sky130_fd_sc_hd__a21oi_1 _14766_ (.A1(_07449_),
    .A2(_07452_),
    .B1(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__and2b_1 _14767_ (.A_N(_07430_),
    .B(_07431_),
    .X(_07455_));
 sky130_fd_sc_hd__xnor2_1 _14768_ (.A(_07429_),
    .B(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__xor2_1 _14769_ (.A(_07448_),
    .B(_07454_),
    .X(_07457_));
 sky130_fd_sc_hd__nand2_1 _14770_ (.A(_07456_),
    .B(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__o21ai_1 _14771_ (.A1(_07448_),
    .A2(_07454_),
    .B1(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__xnor2_1 _14772_ (.A(_07447_),
    .B(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__and2b_1 _14773_ (.A_N(_07447_),
    .B(_07459_),
    .X(_07461_));
 sky130_fd_sc_hd__a21oi_1 _14774_ (.A1(_07446_),
    .A2(_07460_),
    .B1(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__xor2_1 _14775_ (.A(_07445_),
    .B(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__and3_1 _14776_ (.A(_07433_),
    .B(_07440_),
    .C(_07442_),
    .X(_07464_));
 sky130_fd_sc_hd__nor2_1 _14777_ (.A(_07443_),
    .B(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__nor2_1 _14778_ (.A(_07445_),
    .B(_07462_),
    .Y(_07466_));
 sky130_fd_sc_hd__a21oi_1 _14779_ (.A1(_07463_),
    .A2(_07465_),
    .B1(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__xor2_1 _14780_ (.A(_07444_),
    .B(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__nor2_1 _14781_ (.A(_07444_),
    .B(_07467_),
    .Y(_07469_));
 sky130_fd_sc_hd__a21oi_2 _14782_ (.A1(_07443_),
    .A2(_07468_),
    .B1(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__nor2_1 _14783_ (.A(_07427_),
    .B(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__xnor2_1 _14784_ (.A(_07365_),
    .B(_07367_),
    .Y(_07472_));
 sky130_fd_sc_hd__or2_1 _14785_ (.A(_07374_),
    .B(_07424_),
    .X(_07473_));
 sky130_fd_sc_hd__o21a_1 _14786_ (.A1(_07425_),
    .A2(_07426_),
    .B1(_07473_),
    .X(_07474_));
 sky130_fd_sc_hd__nor2_1 _14787_ (.A(_07472_),
    .B(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__nand2_1 _14788_ (.A(_07472_),
    .B(_07474_),
    .Y(_07476_));
 sky130_fd_sc_hd__nor2b_2 _14789_ (.A(_07475_),
    .B_N(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__nand2_1 _14790_ (.A(_07471_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__xor2_2 _14791_ (.A(_07427_),
    .B(_07470_),
    .X(_07479_));
 sky130_fd_sc_hd__xnor2_1 _14792_ (.A(_07443_),
    .B(_07468_),
    .Y(_07480_));
 sky130_fd_sc_hd__xnor2_1 _14793_ (.A(_07434_),
    .B(_07437_),
    .Y(_07481_));
 sky130_fd_sc_hd__nor2_1 _14794_ (.A(_07101_),
    .B(_06969_),
    .Y(_07482_));
 sky130_fd_sc_hd__nor2_1 _14795_ (.A(_07119_),
    .B(_06978_),
    .Y(_07483_));
 sky130_fd_sc_hd__or4_1 _14796_ (.A(_06893_),
    .B(_06917_),
    .C(_06954_),
    .D(_06977_),
    .X(_07484_));
 sky130_fd_sc_hd__o21ai_1 _14797_ (.A1(_07482_),
    .A2(_07483_),
    .B1(_07484_),
    .Y(_07485_));
 sky130_fd_sc_hd__o31ai_1 _14798_ (.A1(_06933_),
    .A2(_07006_),
    .A3(_07485_),
    .B1(_07484_),
    .Y(_07486_));
 sky130_fd_sc_hd__or2b_1 _14799_ (.A(_07481_),
    .B_N(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__xor2_1 _14800_ (.A(_07486_),
    .B(_07481_),
    .X(_07488_));
 sky130_fd_sc_hd__nor2_1 _14801_ (.A(_06865_),
    .B(_06993_),
    .Y(_07489_));
 sky130_fd_sc_hd__o22ai_1 _14802_ (.A1(_06871_),
    .A2(_06966_),
    .B1(_07048_),
    .B2(_06949_),
    .Y(_07490_));
 sky130_fd_sc_hd__or3_1 _14803_ (.A(_06871_),
    .B(_06949_),
    .C(_07435_),
    .X(_07491_));
 sky130_fd_sc_hd__a21bo_1 _14804_ (.A1(_07489_),
    .A2(_07490_),
    .B1_N(_07491_),
    .X(_07492_));
 sky130_fd_sc_hd__or2b_1 _14805_ (.A(_07488_),
    .B_N(_07492_),
    .X(_07493_));
 sky130_fd_sc_hd__clkbuf_4 _14806_ (.A(_07039_),
    .X(_07494_));
 sky130_fd_sc_hd__o22a_1 _14807_ (.A1(_06872_),
    .A2(_07494_),
    .B1(_07273_),
    .B2(_06866_),
    .X(_07495_));
 sky130_fd_sc_hd__or2_1 _14808_ (.A(_07411_),
    .B(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__a21oi_2 _14809_ (.A1(_07487_),
    .A2(_07493_),
    .B1(_07496_),
    .Y(_07497_));
 sky130_fd_sc_hd__xnor2_1 _14810_ (.A(_07463_),
    .B(_07465_),
    .Y(_07498_));
 sky130_fd_sc_hd__xnor2_1 _14811_ (.A(_07446_),
    .B(_07460_),
    .Y(_07499_));
 sky130_fd_sc_hd__or2_1 _14812_ (.A(_07456_),
    .B(_07457_),
    .X(_07500_));
 sky130_fd_sc_hd__nor2_1 _14813_ (.A(_06933_),
    .B(_07006_),
    .Y(_07501_));
 sky130_fd_sc_hd__xnor2_1 _14814_ (.A(_07501_),
    .B(_07485_),
    .Y(_07502_));
 sky130_fd_sc_hd__xnor2_1 _14815_ (.A(_07449_),
    .B(_07452_),
    .Y(_07503_));
 sky130_fd_sc_hd__nor2_1 _14816_ (.A(_06969_),
    .B(_07148_),
    .Y(_07504_));
 sky130_fd_sc_hd__nor2_1 _14817_ (.A(_06939_),
    .B(_07157_),
    .Y(_07505_));
 sky130_fd_sc_hd__o22a_1 _14818_ (.A1(_06899_),
    .A2(_07156_),
    .B1(_07177_),
    .B2(_06939_),
    .X(_07506_));
 sky130_fd_sc_hd__a21oi_2 _14819_ (.A1(_07451_),
    .A2(_07505_),
    .B1(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand2_1 _14820_ (.A(_07451_),
    .B(_07505_),
    .Y(_07508_));
 sky130_fd_sc_hd__a21bo_1 _14821_ (.A1(_07504_),
    .A2(_07507_),
    .B1_N(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__xnor2_1 _14822_ (.A(_07503_),
    .B(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__and2b_1 _14823_ (.A_N(_07503_),
    .B(_07509_),
    .X(_07511_));
 sky130_fd_sc_hd__a21o_1 _14824_ (.A1(_07502_),
    .A2(_07510_),
    .B1(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__xnor2_1 _14825_ (.A(_07492_),
    .B(_07488_),
    .Y(_07513_));
 sky130_fd_sc_hd__xnor2_1 _14826_ (.A(_07456_),
    .B(_07457_),
    .Y(_07514_));
 sky130_fd_sc_hd__xnor2_1 _14827_ (.A(_07514_),
    .B(_07512_),
    .Y(_07515_));
 sky130_fd_sc_hd__a32oi_2 _14828_ (.A1(_07458_),
    .A2(_07500_),
    .A3(_07512_),
    .B1(_07513_),
    .B2(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__xor2_1 _14829_ (.A(_07499_),
    .B(_07516_),
    .X(_07517_));
 sky130_fd_sc_hd__and3_1 _14830_ (.A(_07487_),
    .B(_07493_),
    .C(_07496_),
    .X(_07518_));
 sky130_fd_sc_hd__nor2_1 _14831_ (.A(_07497_),
    .B(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__nor2_1 _14832_ (.A(_07499_),
    .B(_07516_),
    .Y(_07520_));
 sky130_fd_sc_hd__a21oi_1 _14833_ (.A1(_07517_),
    .A2(_07519_),
    .B1(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__xor2_1 _14834_ (.A(_07498_),
    .B(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__nor2_1 _14835_ (.A(_07498_),
    .B(_07521_),
    .Y(_07523_));
 sky130_fd_sc_hd__a21oi_1 _14836_ (.A1(_07497_),
    .A2(_07522_),
    .B1(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__nor2_1 _14837_ (.A(_07480_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__and2_1 _14838_ (.A(_07479_),
    .B(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__nor2_1 _14839_ (.A(_07471_),
    .B(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__xnor2_2 _14840_ (.A(_07477_),
    .B(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__xnor2_1 _14841_ (.A(_07497_),
    .B(_07522_),
    .Y(_07529_));
 sky130_fd_sc_hd__clkbuf_4 _14842_ (.A(_06970_),
    .X(_07530_));
 sky130_fd_sc_hd__nor2_1 _14843_ (.A(_06933_),
    .B(_07048_),
    .Y(_07531_));
 sky130_fd_sc_hd__nor2_1 _14844_ (.A(_07101_),
    .B(_06978_),
    .Y(_07532_));
 sky130_fd_sc_hd__nor2_1 _14845_ (.A(_07119_),
    .B(_07005_),
    .Y(_07533_));
 sky130_fd_sc_hd__nor4_1 _14846_ (.A(_07119_),
    .B(_06917_),
    .C(_06978_),
    .D(_07005_),
    .Y(_07534_));
 sky130_fd_sc_hd__o21ba_1 _14847_ (.A1(_07532_),
    .A2(_07533_),
    .B1_N(_07534_),
    .X(_07535_));
 sky130_fd_sc_hd__a21oi_1 _14848_ (.A1(_07531_),
    .A2(_07535_),
    .B1(_07534_),
    .Y(_07536_));
 sky130_fd_sc_hd__nand2_1 _14849_ (.A(_07491_),
    .B(_07490_),
    .Y(_07537_));
 sky130_fd_sc_hd__xor2_1 _14850_ (.A(_07489_),
    .B(_07537_),
    .X(_07538_));
 sky130_fd_sc_hd__xnor2_1 _14851_ (.A(_07536_),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__or2_1 _14852_ (.A(_06865_),
    .B(_06968_),
    .X(_07540_));
 sky130_fd_sc_hd__clkbuf_2 _14853_ (.A(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__or2_1 _14854_ (.A(_07536_),
    .B(_07538_),
    .X(_07542_));
 sky130_fd_sc_hd__o41a_1 _14855_ (.A1(_06873_),
    .A2(_07530_),
    .A3(_07539_),
    .A4(_07541_),
    .B1(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__nor2_1 _14856_ (.A(_07410_),
    .B(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__xnor2_1 _14857_ (.A(_07517_),
    .B(_07519_),
    .Y(_07545_));
 sky130_fd_sc_hd__and2_1 _14858_ (.A(_07410_),
    .B(_07543_),
    .X(_07546_));
 sky130_fd_sc_hd__nor2_1 _14859_ (.A(_07544_),
    .B(_07546_),
    .Y(_07547_));
 sky130_fd_sc_hd__xnor2_1 _14860_ (.A(_07513_),
    .B(_07515_),
    .Y(_07548_));
 sky130_fd_sc_hd__nor3_1 _14861_ (.A(_06872_),
    .B(_06970_),
    .C(_07541_),
    .Y(_07549_));
 sky130_fd_sc_hd__xnor2_1 _14862_ (.A(_07539_),
    .B(_07549_),
    .Y(_07550_));
 sky130_fd_sc_hd__xor2_1 _14863_ (.A(_07502_),
    .B(_07510_),
    .X(_07551_));
 sky130_fd_sc_hd__xor2_1 _14864_ (.A(_07531_),
    .B(_07535_),
    .X(_07552_));
 sky130_fd_sc_hd__xnor2_2 _14865_ (.A(_07504_),
    .B(_07507_),
    .Y(_07553_));
 sky130_fd_sc_hd__nor4_1 _14866_ (.A(_06939_),
    .B(_06954_),
    .C(_07156_),
    .D(_07177_),
    .Y(_07554_));
 sky130_fd_sc_hd__o22a_1 _14867_ (.A1(_06938_),
    .A2(_07156_),
    .B1(_07177_),
    .B2(_06954_),
    .X(_07555_));
 sky130_fd_sc_hd__or4_1 _14868_ (.A(_06977_),
    .B(_07147_),
    .C(_07554_),
    .D(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__or2b_1 _14869_ (.A(_07554_),
    .B_N(_07556_),
    .X(_07557_));
 sky130_fd_sc_hd__xnor2_1 _14870_ (.A(_07553_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__and2b_1 _14871_ (.A_N(_07553_),
    .B(_07557_),
    .X(_07559_));
 sky130_fd_sc_hd__a21oi_1 _14872_ (.A1(_07552_),
    .A2(_07558_),
    .B1(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__xnor2_1 _14873_ (.A(_07551_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__and2b_1 _14874_ (.A_N(_07560_),
    .B(_07551_),
    .X(_07562_));
 sky130_fd_sc_hd__a21oi_1 _14875_ (.A1(_07550_),
    .A2(_07561_),
    .B1(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__nor2_1 _14876_ (.A(_07548_),
    .B(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__and2_1 _14877_ (.A(_07548_),
    .B(_07563_),
    .X(_07565_));
 sky130_fd_sc_hd__nor2_1 _14878_ (.A(_07564_),
    .B(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__a21o_1 _14879_ (.A1(_07547_),
    .A2(_07566_),
    .B1(_07564_),
    .X(_07567_));
 sky130_fd_sc_hd__xnor2_1 _14880_ (.A(_07545_),
    .B(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__or2b_1 _14881_ (.A(_07545_),
    .B_N(_07567_),
    .X(_07569_));
 sky130_fd_sc_hd__a21boi_2 _14882_ (.A1(_07544_),
    .A2(_07568_),
    .B1_N(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__or2_1 _14883_ (.A(_07529_),
    .B(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__xor2_1 _14884_ (.A(_07480_),
    .B(_07524_),
    .X(_07572_));
 sky130_fd_sc_hd__and2b_1 _14885_ (.A_N(_07571_),
    .B(_07572_),
    .X(_07573_));
 sky130_fd_sc_hd__xor2_1 _14886_ (.A(_07529_),
    .B(_07570_),
    .X(_07574_));
 sky130_fd_sc_hd__xor2_1 _14887_ (.A(_07544_),
    .B(_07568_),
    .X(_07575_));
 sky130_fd_sc_hd__xor2_1 _14888_ (.A(_07547_),
    .B(_07566_),
    .X(_07576_));
 sky130_fd_sc_hd__nor2_1 _14889_ (.A(_07101_),
    .B(_07048_),
    .Y(_07577_));
 sky130_fd_sc_hd__o22a_1 _14890_ (.A1(_07101_),
    .A2(_07006_),
    .B1(_07048_),
    .B2(_07119_),
    .X(_07578_));
 sky130_fd_sc_hd__or2_1 _14891_ (.A(_06872_),
    .B(_06933_),
    .X(_07579_));
 sky130_fd_sc_hd__o2bb2a_1 _14892_ (.A1_N(_07533_),
    .A2_N(_07577_),
    .B1(_07578_),
    .B2(_07579_),
    .X(_07580_));
 sky130_fd_sc_hd__buf_2 _14893_ (.A(_06968_),
    .X(_07581_));
 sky130_fd_sc_hd__o22a_1 _14894_ (.A1(_06873_),
    .A2(_07581_),
    .B1(_07530_),
    .B2(_06866_),
    .X(_07582_));
 sky130_fd_sc_hd__nor3_1 _14895_ (.A(_07549_),
    .B(_07580_),
    .C(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__xnor2_1 _14896_ (.A(_07550_),
    .B(_07561_),
    .Y(_07584_));
 sky130_fd_sc_hd__xnor2_1 _14897_ (.A(_07552_),
    .B(_07558_),
    .Y(_07585_));
 sky130_fd_sc_hd__o22a_1 _14898_ (.A1(_06978_),
    .A2(_07148_),
    .B1(_07554_),
    .B2(_07555_),
    .X(_07586_));
 sky130_fd_sc_hd__inv_2 _14899_ (.A(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__nand2_2 _14900_ (.A(_07556_),
    .B(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__or2_1 _14901_ (.A(_07006_),
    .B(_07148_),
    .X(_07589_));
 sky130_fd_sc_hd__or4_1 _14902_ (.A(_06969_),
    .B(_06977_),
    .C(_07157_),
    .D(_07178_),
    .X(_07590_));
 sky130_fd_sc_hd__o22ai_1 _14903_ (.A1(_06969_),
    .A2(_07157_),
    .B1(_07178_),
    .B2(_06978_),
    .Y(_07591_));
 sky130_fd_sc_hd__nand2_1 _14904_ (.A(_07590_),
    .B(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__o21a_1 _14905_ (.A1(_07589_),
    .A2(_07592_),
    .B1(_07590_),
    .X(_07593_));
 sky130_fd_sc_hd__xor2_1 _14906_ (.A(_07588_),
    .B(_07593_),
    .X(_07594_));
 sky130_fd_sc_hd__a21o_1 _14907_ (.A1(_07533_),
    .A2(_07577_),
    .B1(_07578_),
    .X(_07595_));
 sky130_fd_sc_hd__xor2_1 _14908_ (.A(_07579_),
    .B(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__nor2_1 _14909_ (.A(_07588_),
    .B(_07593_),
    .Y(_07597_));
 sky130_fd_sc_hd__a21oi_1 _14910_ (.A1(_07594_),
    .A2(_07596_),
    .B1(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__nor2_1 _14911_ (.A(_07585_),
    .B(_07598_),
    .Y(_07599_));
 sky130_fd_sc_hd__and2_1 _14912_ (.A(_07585_),
    .B(_07598_),
    .X(_07600_));
 sky130_fd_sc_hd__nor2_1 _14913_ (.A(_07599_),
    .B(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__o21a_1 _14914_ (.A1(_07549_),
    .A2(_07582_),
    .B1(_07580_),
    .X(_07602_));
 sky130_fd_sc_hd__nor2_1 _14915_ (.A(_07583_),
    .B(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__a21oi_1 _14916_ (.A1(_07601_),
    .A2(_07603_),
    .B1(_07599_),
    .Y(_07604_));
 sky130_fd_sc_hd__or2_1 _14917_ (.A(_07584_),
    .B(_07604_),
    .X(_07605_));
 sky130_fd_sc_hd__nand2_1 _14918_ (.A(_07584_),
    .B(_07604_),
    .Y(_07606_));
 sky130_fd_sc_hd__and2_1 _14919_ (.A(_07605_),
    .B(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__a21bo_1 _14920_ (.A1(_07583_),
    .A2(_07607_),
    .B1_N(_07605_),
    .X(_07608_));
 sky130_fd_sc_hd__and3_1 _14921_ (.A(_07575_),
    .B(_07576_),
    .C(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__and2_1 _14922_ (.A(_07574_),
    .B(_07609_),
    .X(_07610_));
 sky130_fd_sc_hd__xor2_1 _14923_ (.A(_07574_),
    .B(_07609_),
    .X(_07611_));
 sky130_fd_sc_hd__nand2_1 _14924_ (.A(_07576_),
    .B(_07608_),
    .Y(_07612_));
 sky130_fd_sc_hd__or2b_1 _14925_ (.A(_07576_),
    .B_N(_07605_),
    .X(_07613_));
 sky130_fd_sc_hd__xnor2_1 _14926_ (.A(_07601_),
    .B(_07603_),
    .Y(_07614_));
 sky130_fd_sc_hd__xnor2_1 _14927_ (.A(_07594_),
    .B(_07596_),
    .Y(_07615_));
 sky130_fd_sc_hd__or2_1 _14928_ (.A(_06866_),
    .B(_07100_),
    .X(_07616_));
 sky130_fd_sc_hd__buf_2 _14929_ (.A(_07119_),
    .X(_07617_));
 sky130_fd_sc_hd__nor2_1 _14930_ (.A(_06872_),
    .B(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__or4_1 _14931_ (.A(_06872_),
    .B(_07119_),
    .C(_07101_),
    .D(_07048_),
    .X(_07619_));
 sky130_fd_sc_hd__o21a_1 _14932_ (.A1(_07577_),
    .A2(_07618_),
    .B1(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__xnor2_1 _14933_ (.A(_07616_),
    .B(_07620_),
    .Y(_07621_));
 sky130_fd_sc_hd__xnor2_1 _14934_ (.A(_07589_),
    .B(_07592_),
    .Y(_07622_));
 sky130_fd_sc_hd__or2_1 _14935_ (.A(_07049_),
    .B(_07213_),
    .X(_07623_));
 sky130_fd_sc_hd__o22a_1 _14936_ (.A1(_06979_),
    .A2(_07185_),
    .B1(_07199_),
    .B2(_07006_),
    .X(_07624_));
 sky130_fd_sc_hd__or4_1 _14937_ (.A(_06978_),
    .B(_07006_),
    .C(_07157_),
    .D(_07178_),
    .X(_07625_));
 sky130_fd_sc_hd__o21a_1 _14938_ (.A1(_07623_),
    .A2(_07624_),
    .B1(_07625_),
    .X(_07626_));
 sky130_fd_sc_hd__nand2_1 _14939_ (.A(_07622_),
    .B(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__nor2_1 _14940_ (.A(_07622_),
    .B(_07626_),
    .Y(_07628_));
 sky130_fd_sc_hd__a21oi_1 _14941_ (.A1(_07621_),
    .A2(_07627_),
    .B1(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__xor2_1 _14942_ (.A(_07615_),
    .B(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__inv_2 _14943_ (.A(_07620_),
    .Y(_07631_));
 sky130_fd_sc_hd__o21a_1 _14944_ (.A1(_07616_),
    .A2(_07631_),
    .B1(_07619_),
    .X(_07632_));
 sky130_fd_sc_hd__xor2_1 _14945_ (.A(_07541_),
    .B(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__nand2_1 _14946_ (.A(_07630_),
    .B(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__o21a_1 _14947_ (.A1(_07615_),
    .A2(_07629_),
    .B1(_07634_),
    .X(_07635_));
 sky130_fd_sc_hd__or2_1 _14948_ (.A(_07614_),
    .B(_07635_),
    .X(_07636_));
 sky130_fd_sc_hd__xnor2_1 _14949_ (.A(_07614_),
    .B(_07635_),
    .Y(_07637_));
 sky130_fd_sc_hd__or3_1 _14950_ (.A(_07541_),
    .B(_07632_),
    .C(_07637_),
    .X(_07638_));
 sky130_fd_sc_hd__xnor2_1 _14951_ (.A(_07583_),
    .B(_07607_),
    .Y(_07639_));
 sky130_fd_sc_hd__a21oi_1 _14952_ (.A1(_07636_),
    .A2(_07638_),
    .B1(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__and4_1 _14953_ (.A(_07575_),
    .B(_07612_),
    .C(_07613_),
    .D(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__xor2_1 _14954_ (.A(_07611_),
    .B(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__o21ai_1 _14955_ (.A1(_07541_),
    .A2(_07632_),
    .B1(_07637_),
    .Y(_07643_));
 sky130_fd_sc_hd__or2_1 _14956_ (.A(_07630_),
    .B(_07633_),
    .X(_07644_));
 sky130_fd_sc_hd__nand2_1 _14957_ (.A(_07634_),
    .B(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__buf_2 _14958_ (.A(_07101_),
    .X(_07646_));
 sky130_fd_sc_hd__or2_1 _14959_ (.A(_06866_),
    .B(_07646_),
    .X(_07647_));
 sky130_fd_sc_hd__or3_1 _14960_ (.A(_06873_),
    .B(_07617_),
    .C(_07647_),
    .X(_07648_));
 sky130_fd_sc_hd__and2b_1 _14961_ (.A_N(_07628_),
    .B(_07627_),
    .X(_07649_));
 sky130_fd_sc_hd__xnor2_1 _14962_ (.A(_07621_),
    .B(_07649_),
    .Y(_07650_));
 sky130_fd_sc_hd__inv_2 _14963_ (.A(_07625_),
    .Y(_07651_));
 sky130_fd_sc_hd__nor2_1 _14964_ (.A(_07651_),
    .B(_07624_),
    .Y(_07652_));
 sky130_fd_sc_hd__xor2_1 _14965_ (.A(_07623_),
    .B(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__nor2_1 _14966_ (.A(_06872_),
    .B(_07148_),
    .Y(_07654_));
 sky130_fd_sc_hd__nor2_1 _14967_ (.A(_07048_),
    .B(_07157_),
    .Y(_07655_));
 sky130_fd_sc_hd__and3b_1 _14968_ (.A_N(_07006_),
    .B(_07174_),
    .C(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__o22a_1 _14969_ (.A1(_07006_),
    .A2(_07157_),
    .B1(_07178_),
    .B2(_07048_),
    .X(_07657_));
 sky130_fd_sc_hd__nor2_1 _14970_ (.A(_07656_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__a21oi_1 _14971_ (.A1(_07654_),
    .A2(_07658_),
    .B1(_07656_),
    .Y(_07659_));
 sky130_fd_sc_hd__xor2_1 _14972_ (.A(_07653_),
    .B(_07659_),
    .X(_07660_));
 sky130_fd_sc_hd__buf_2 _14973_ (.A(_07617_),
    .X(_07661_));
 sky130_fd_sc_hd__buf_2 _14974_ (.A(_07646_),
    .X(_07662_));
 sky130_fd_sc_hd__o22ai_1 _14975_ (.A1(_06866_),
    .A2(_07661_),
    .B1(_07662_),
    .B2(_06873_),
    .Y(_07663_));
 sky130_fd_sc_hd__and2_1 _14976_ (.A(_07648_),
    .B(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__and2_1 _14977_ (.A(_07660_),
    .B(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__o21ba_1 _14978_ (.A1(_07653_),
    .A2(_07659_),
    .B1_N(_07665_),
    .X(_07666_));
 sky130_fd_sc_hd__xnor2_1 _14979_ (.A(_07650_),
    .B(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__xor2_1 _14980_ (.A(_07654_),
    .B(_07658_),
    .X(_07668_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(_06872_),
    .B(_07199_),
    .Y(_07669_));
 sky130_fd_sc_hd__nand2_1 _14982_ (.A(_06787_),
    .B(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__nor2_1 _14983_ (.A(_07049_),
    .B(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__inv_2 _14984_ (.A(_06865_),
    .Y(_07672_));
 sky130_fd_sc_hd__a221o_4 _14985_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_06855_),
    .B1(_07144_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .C1(_07146_),
    .X(_07673_));
 sky130_fd_sc_hd__o211a_1 _14986_ (.A1(_07655_),
    .A2(_07669_),
    .B1(_07672_),
    .C1(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__nor3_1 _14987_ (.A(_07668_),
    .B(_07671_),
    .C(_07674_),
    .Y(_07675_));
 sky130_fd_sc_hd__o21ai_1 _14988_ (.A1(_07671_),
    .A2(_07674_),
    .B1(_07668_),
    .Y(_07676_));
 sky130_fd_sc_hd__or3_1 _14989_ (.A(_07668_),
    .B(_07671_),
    .C(_07674_),
    .X(_07677_));
 sky130_fd_sc_hd__nand2_1 _14990_ (.A(_07676_),
    .B(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__nand2_1 _14991_ (.A(_07265_),
    .B(_07213_),
    .Y(_07679_));
 sky130_fd_sc_hd__or2_1 _14992_ (.A(_07011_),
    .B(_07670_),
    .X(_07680_));
 sky130_fd_sc_hd__a221o_1 _14993_ (.A1(_07647_),
    .A2(_07678_),
    .B1(_07679_),
    .B2(_07623_),
    .C1(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__o211a_1 _14994_ (.A1(_07647_),
    .A2(_07675_),
    .B1(_07681_),
    .C1(_07676_),
    .X(_07682_));
 sky130_fd_sc_hd__nor2_1 _14995_ (.A(_07660_),
    .B(_07664_),
    .Y(_07683_));
 sky130_fd_sc_hd__o32a_1 _14996_ (.A1(_07665_),
    .A2(_07682_),
    .A3(_07683_),
    .B1(_07676_),
    .B2(_07681_),
    .X(_07684_));
 sky130_fd_sc_hd__a21o_1 _14997_ (.A1(_07648_),
    .A2(_07667_),
    .B1(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__o21a_1 _14998_ (.A1(_07648_),
    .A2(_07667_),
    .B1(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__a211o_1 _14999_ (.A1(_07645_),
    .A2(_07685_),
    .B1(_07666_),
    .C1(_07650_),
    .X(_07687_));
 sky130_fd_sc_hd__o21ai_1 _15000_ (.A1(_07645_),
    .A2(_07686_),
    .B1(_07687_),
    .Y(_07688_));
 sky130_fd_sc_hd__and4_1 _15001_ (.A(_07612_),
    .B(_07638_),
    .C(_07643_),
    .D(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__o2bb2a_1 _15002_ (.A1_N(_07639_),
    .A2_N(_07636_),
    .B1(_07576_),
    .B2(_07608_),
    .X(_07690_));
 sky130_fd_sc_hd__o2111a_2 _15003_ (.A1(_07639_),
    .A2(_07636_),
    .B1(_07689_),
    .C1(_07690_),
    .D1(_07575_),
    .X(_07691_));
 sky130_fd_sc_hd__and2_1 _15004_ (.A(_07611_),
    .B(_07641_),
    .X(_07692_));
 sky130_fd_sc_hd__a21o_1 _15005_ (.A1(_07642_),
    .A2(_07691_),
    .B1(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__xnor2_1 _15006_ (.A(_07572_),
    .B(_07610_),
    .Y(_07694_));
 sky130_fd_sc_hd__a21oi_1 _15007_ (.A1(_07571_),
    .A2(_07694_),
    .B1(_07573_),
    .Y(_07695_));
 sky130_fd_sc_hd__a22o_2 _15008_ (.A1(_07572_),
    .A2(_07610_),
    .B1(_07693_),
    .B2(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__nor2_1 _15009_ (.A(_07525_),
    .B(_07573_),
    .Y(_07697_));
 sky130_fd_sc_hd__xnor2_2 _15010_ (.A(_07479_),
    .B(_07697_),
    .Y(_07698_));
 sky130_fd_sc_hd__a22o_2 _15011_ (.A1(_07479_),
    .A2(_07573_),
    .B1(_07696_),
    .B2(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__a22o_2 _15012_ (.A1(_07477_),
    .A2(_07526_),
    .B1(_07528_),
    .B2(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__a21o_1 _15013_ (.A1(_07471_),
    .A2(_07476_),
    .B1(_07475_),
    .X(_07701_));
 sky130_fd_sc_hd__xnor2_4 _15014_ (.A(_07372_),
    .B(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__a2bb2o_4 _15015_ (.A1_N(_07372_),
    .A2_N(_07478_),
    .B1(_07700_),
    .B2(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__a21o_1 _15016_ (.A1(_07272_),
    .A2(_07285_),
    .B1(_07283_),
    .X(_07704_));
 sky130_fd_sc_hd__or2b_1 _15017_ (.A(_07127_),
    .B_N(_07086_),
    .X(_07705_));
 sky130_fd_sc_hd__nor2_1 _15018_ (.A(_06875_),
    .B(_07007_),
    .Y(_07706_));
 sky130_fd_sc_hd__nor2_1 _15019_ (.A(_06857_),
    .B(_06979_),
    .Y(_07707_));
 sky130_fd_sc_hd__nor2_1 _15020_ (.A(_06874_),
    .B(_06979_),
    .Y(_07708_));
 sky130_fd_sc_hd__nand2_1 _15021_ (.A(_07266_),
    .B(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__o21ai_1 _15022_ (.A1(_07706_),
    .A2(_07707_),
    .B1(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__nor2_1 _15023_ (.A(_07265_),
    .B(_07270_),
    .Y(_07711_));
 sky130_fd_sc_hd__xnor2_1 _15024_ (.A(_07710_),
    .B(_07711_),
    .Y(_07712_));
 sky130_fd_sc_hd__or2_1 _15025_ (.A(_06900_),
    .B(_07037_),
    .X(_07713_));
 sky130_fd_sc_hd__or3_1 _15026_ (.A(_06940_),
    .B(_07039_),
    .C(_07713_),
    .X(_07714_));
 sky130_fd_sc_hd__o22ai_1 _15027_ (.A1(_07097_),
    .A2(_07039_),
    .B1(_07273_),
    .B2(_06940_),
    .Y(_07715_));
 sky130_fd_sc_hd__nand2_1 _15028_ (.A(_07714_),
    .B(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__or2_1 _15029_ (.A(_07235_),
    .B(_07052_),
    .X(_07717_));
 sky130_fd_sc_hd__xnor2_1 _15030_ (.A(_07716_),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__o31a_1 _15031_ (.A1(_06979_),
    .A2(_07281_),
    .A3(_07275_),
    .B1(_07274_),
    .X(_07719_));
 sky130_fd_sc_hd__nor2_1 _15032_ (.A(_07718_),
    .B(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__and2_1 _15033_ (.A(_07718_),
    .B(_07719_),
    .X(_07721_));
 sky130_fd_sc_hd__nor2_1 _15034_ (.A(_07720_),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__xnor2_1 _15035_ (.A(_07712_),
    .B(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__a21o_1 _15036_ (.A1(_07125_),
    .A2(_07705_),
    .B1(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__nand3_1 _15037_ (.A(_07125_),
    .B(_07705_),
    .C(_07723_),
    .Y(_07725_));
 sky130_fd_sc_hd__nand2_1 _15038_ (.A(_07724_),
    .B(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__xnor2_1 _15039_ (.A(_07704_),
    .B(_07726_),
    .Y(_07727_));
 sky130_fd_sc_hd__a21bo_1 _15040_ (.A1(_07096_),
    .A2(_07098_),
    .B1_N(_07095_),
    .X(_07728_));
 sky130_fd_sc_hd__inv_2 _15041_ (.A(_07110_),
    .Y(_07729_));
 sky130_fd_sc_hd__nor2_1 _15042_ (.A(_07617_),
    .B(_07137_),
    .Y(_07730_));
 sky130_fd_sc_hd__a22o_1 _15043_ (.A1(_07729_),
    .A2(_07730_),
    .B1(_07139_),
    .B2(_07142_),
    .X(_07731_));
 sky130_fd_sc_hd__or2_1 _15044_ (.A(_06968_),
    .B(_07141_),
    .X(_07732_));
 sky130_fd_sc_hd__nor2_1 _15045_ (.A(_06970_),
    .B(_07141_),
    .Y(_07733_));
 sky130_fd_sc_hd__a22o_1 _15046_ (.A1(_07094_),
    .A2(_07732_),
    .B1(_07733_),
    .B2(_07093_),
    .X(_07734_));
 sky130_fd_sc_hd__buf_2 _15047_ (.A(_07078_),
    .X(_07735_));
 sky130_fd_sc_hd__nor2_1 _15048_ (.A(_07735_),
    .B(_06993_),
    .Y(_07736_));
 sky130_fd_sc_hd__xnor2_1 _15049_ (.A(_07734_),
    .B(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__nand2_1 _15050_ (.A(_07731_),
    .B(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__or2_1 _15051_ (.A(_07731_),
    .B(_07737_),
    .X(_07739_));
 sky130_fd_sc_hd__nand2_1 _15052_ (.A(_07738_),
    .B(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__xnor2_1 _15053_ (.A(_07728_),
    .B(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__nor2_1 _15054_ (.A(_07646_),
    .B(_07198_),
    .Y(_07742_));
 sky130_fd_sc_hd__or4_1 _15055_ (.A(_07119_),
    .B(_07101_),
    .C(_07136_),
    .D(_07198_),
    .X(_07743_));
 sky130_fd_sc_hd__o21ai_2 _15056_ (.A1(_07730_),
    .A2(_07742_),
    .B1(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__nor2_1 _15057_ (.A(_07100_),
    .B(_07138_),
    .Y(_07745_));
 sky130_fd_sc_hd__xnor2_2 _15058_ (.A(_07744_),
    .B(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__or2_1 _15059_ (.A(_07158_),
    .B(_07167_),
    .X(_07747_));
 sky130_fd_sc_hd__buf_2 _15060_ (.A(_07747_),
    .X(_07748_));
 sky130_fd_sc_hd__or2_1 _15061_ (.A(_07148_),
    .B(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__or3_1 _15062_ (.A(_06759_),
    .B(_06764_),
    .C(_07165_),
    .X(_07750_));
 sky130_fd_sc_hd__o21ai_1 _15063_ (.A1(_06759_),
    .A2(_07165_),
    .B1(_06765_),
    .Y(_07751_));
 sky130_fd_sc_hd__a31o_1 _15064_ (.A1(_04831_),
    .A2(_07750_),
    .A3(_07751_),
    .B1(_07162_),
    .X(_07752_));
 sky130_fd_sc_hd__a21oi_1 _15065_ (.A1(_03492_),
    .A2(\rbzero.wall_tracer.stepDistY[5] ),
    .B1(_04948_),
    .Y(_07753_));
 sky130_fd_sc_hd__a2bb2o_1 _15066_ (.A1_N(_04840_),
    .A2_N(\rbzero.wall_tracer.stepDistX[5] ),
    .B1(_07752_),
    .B2(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__or3_1 _15067_ (.A(_07178_),
    .B(_07176_),
    .C(_07754_),
    .X(_07755_));
 sky130_fd_sc_hd__a2bb2o_2 _15068_ (.A1_N(_04841_),
    .A2_N(\rbzero.wall_tracer.stepDistX[4] ),
    .B1(_07171_),
    .B2(_07172_),
    .X(_07756_));
 sky130_fd_sc_hd__buf_2 _15069_ (.A(_07754_),
    .X(_07757_));
 sky130_fd_sc_hd__o22ai_1 _15070_ (.A1(_07756_),
    .A2(_07199_),
    .B1(_07757_),
    .B2(_07185_),
    .Y(_07758_));
 sky130_fd_sc_hd__nand2_1 _15071_ (.A(_07755_),
    .B(_07758_),
    .Y(_07759_));
 sky130_fd_sc_hd__xnor2_2 _15072_ (.A(_07749_),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__or2b_1 _15073_ (.A(_07155_),
    .B_N(_07180_),
    .X(_07761_));
 sky130_fd_sc_hd__o41a_1 _15074_ (.A1(_07185_),
    .A2(_07748_),
    .A3(_07756_),
    .A4(_07199_),
    .B1(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__xor2_2 _15075_ (.A(_07760_),
    .B(_07762_),
    .X(_07763_));
 sky130_fd_sc_hd__xnor2_2 _15076_ (.A(_07746_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__inv_2 _15077_ (.A(_07761_),
    .Y(_07765_));
 sky130_fd_sc_hd__clkbuf_4 _15078_ (.A(_07198_),
    .X(_07766_));
 sky130_fd_sc_hd__o21ba_1 _15079_ (.A1(_07213_),
    .A2(_07766_),
    .B1_N(_07180_),
    .X(_07767_));
 sky130_fd_sc_hd__nand2_1 _15080_ (.A(_07143_),
    .B(_07188_),
    .Y(_07768_));
 sky130_fd_sc_hd__o31a_1 _15081_ (.A1(_07765_),
    .A2(_07767_),
    .A3(_07187_),
    .B1(_07768_),
    .X(_07769_));
 sky130_fd_sc_hd__xor2_2 _15082_ (.A(_07764_),
    .B(_07769_),
    .X(_07770_));
 sky130_fd_sc_hd__xnor2_1 _15083_ (.A(_07741_),
    .B(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__a21oi_1 _15084_ (.A1(_07128_),
    .A2(_07207_),
    .B1(_07206_),
    .Y(_07772_));
 sky130_fd_sc_hd__nor2_1 _15085_ (.A(_07771_),
    .B(_07772_),
    .Y(_07773_));
 sky130_fd_sc_hd__nand2_1 _15086_ (.A(_07771_),
    .B(_07772_),
    .Y(_07774_));
 sky130_fd_sc_hd__and2b_1 _15087_ (.A_N(_07773_),
    .B(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__xnor2_1 _15088_ (.A(_07727_),
    .B(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__a21oi_1 _15089_ (.A1(_07246_),
    .A2(_07290_),
    .B1(_07244_),
    .Y(_07777_));
 sky130_fd_sc_hd__nor2_1 _15090_ (.A(_07776_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__and2_1 _15091_ (.A(_07776_),
    .B(_07777_),
    .X(_07779_));
 sky130_fd_sc_hd__nor2_2 _15092_ (.A(_07778_),
    .B(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__or2b_1 _15093_ (.A(_07289_),
    .B_N(_07262_),
    .X(_07781_));
 sky130_fd_sc_hd__and2_1 _15094_ (.A(_07331_),
    .B(_07334_),
    .X(_07782_));
 sky130_fd_sc_hd__a21bo_1 _15095_ (.A1(_07267_),
    .A2(_07271_),
    .B1_N(_07264_),
    .X(_07783_));
 sky130_fd_sc_hd__and2_1 _15096_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_07256_),
    .X(_07784_));
 sky130_fd_sc_hd__and3b_1 _15097_ (.A_N(_07269_),
    .B(_07334_),
    .C(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__nand2_2 _15098_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_06855_),
    .Y(_07786_));
 sky130_fd_sc_hd__buf_2 _15099_ (.A(_07786_),
    .X(_07787_));
 sky130_fd_sc_hd__o22a_1 _15100_ (.A1(_07269_),
    .A2(_07333_),
    .B1(_07787_),
    .B2(_07011_),
    .X(_07788_));
 sky130_fd_sc_hd__nor2_1 _15101_ (.A(_07785_),
    .B(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__nand2_1 _15102_ (.A(_07783_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__or2_1 _15103_ (.A(_07783_),
    .B(_07789_),
    .X(_07791_));
 sky130_fd_sc_hd__and2_1 _15104_ (.A(_07790_),
    .B(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__nand2_1 _15105_ (.A(_07782_),
    .B(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__or2_1 _15106_ (.A(_07782_),
    .B(_07792_),
    .X(_07794_));
 sky130_fd_sc_hd__nand2_1 _15107_ (.A(_07793_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__a21oi_2 _15108_ (.A1(_07287_),
    .A2(_07781_),
    .B1(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__and3_1 _15109_ (.A(_07287_),
    .B(_07781_),
    .C(_07795_),
    .X(_07797_));
 sky130_fd_sc_hd__nor2_2 _15110_ (.A(_07796_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__xnor2_4 _15111_ (.A(_07780_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__nor2_1 _15112_ (.A(_07291_),
    .B(_07328_),
    .Y(_07800_));
 sky130_fd_sc_hd__a21oi_4 _15113_ (.A1(_07329_),
    .A2(_07338_),
    .B1(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__xor2_4 _15114_ (.A(_07799_),
    .B(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__xnor2_4 _15115_ (.A(_07336_),
    .B(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__a21o_2 _15116_ (.A1(_07076_),
    .A2(_07371_),
    .B1(_07369_),
    .X(_07804_));
 sky130_fd_sc_hd__xor2_4 _15117_ (.A(_07803_),
    .B(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__and2b_2 _15118_ (.A_N(_07372_),
    .B(_07475_),
    .X(_07806_));
 sky130_fd_sc_hd__xnor2_4 _15119_ (.A(_07805_),
    .B(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__xor2_4 _15120_ (.A(_07703_),
    .B(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__mux2_1 _15121_ (.A0(\rbzero.debug_overlay.playerY[-6] ),
    .A1(\rbzero.debug_overlay.playerX[-6] ),
    .S(_06851_),
    .X(_07809_));
 sky130_fd_sc_hd__nand2_1 _15122_ (.A(_07808_),
    .B(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__or2_1 _15123_ (.A(_07808_),
    .B(_07809_),
    .X(_07811_));
 sky130_fd_sc_hd__nand2_1 _15124_ (.A(_07810_),
    .B(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__xor2_4 _15125_ (.A(_07700_),
    .B(_07702_),
    .X(_07813_));
 sky130_fd_sc_hd__mux2_1 _15126_ (.A0(\rbzero.debug_overlay.playerY[-7] ),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_06850_),
    .X(_07814_));
 sky130_fd_sc_hd__xor2_4 _15127_ (.A(_07699_),
    .B(_07528_),
    .X(_07815_));
 sky130_fd_sc_hd__mux2_1 _15128_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_06850_),
    .X(_07816_));
 sky130_fd_sc_hd__xor2_4 _15129_ (.A(_07696_),
    .B(_07698_),
    .X(_07817_));
 sky130_fd_sc_hd__mux2_1 _15130_ (.A0(\rbzero.debug_overlay.playerY[-9] ),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_06850_),
    .X(_07818_));
 sky130_fd_sc_hd__a22o_1 _15131_ (.A1(_07817_),
    .A2(_07818_),
    .B1(_07815_),
    .B2(_07816_),
    .X(_07819_));
 sky130_fd_sc_hd__o221a_1 _15132_ (.A1(_07813_),
    .A2(_07814_),
    .B1(_07815_),
    .B2(_07816_),
    .C1(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__a21oi_1 _15133_ (.A1(_07813_),
    .A2(_07814_),
    .B1(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__or2_1 _15134_ (.A(_07812_),
    .B(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__nand2_1 _15135_ (.A(_07812_),
    .B(_07821_),
    .Y(_07823_));
 sky130_fd_sc_hd__nand2_1 _15136_ (.A(_07822_),
    .B(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__clkbuf_4 _15137_ (.A(_06914_),
    .X(_07825_));
 sky130_fd_sc_hd__clkbuf_4 _15138_ (.A(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__mux2_2 _15139_ (.A0(_07826_),
    .A1(_04929_),
    .S(_06851_),
    .X(_07827_));
 sky130_fd_sc_hd__nor2_1 _15140_ (.A(_07824_),
    .B(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__a21o_1 _15141_ (.A1(_07824_),
    .A2(_07827_),
    .B1(_04832_),
    .X(_07829_));
 sky130_fd_sc_hd__o221a_1 _15142_ (.A1(\rbzero.wall_tracer.texu[0] ),
    .A2(_06853_),
    .B1(_07828_),
    .B2(_07829_),
    .C1(_03498_),
    .X(_00475_));
 sky130_fd_sc_hd__or2b_2 _15143_ (.A(_07803_),
    .B_N(_07804_),
    .X(_07830_));
 sky130_fd_sc_hd__and2b_1 _15144_ (.A_N(_07805_),
    .B(_07806_),
    .X(_07831_));
 sky130_fd_sc_hd__a21oi_2 _15145_ (.A1(_07703_),
    .A2(_07807_),
    .B1(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__or2b_1 _15146_ (.A(_07726_),
    .B_N(_07704_),
    .X(_07833_));
 sky130_fd_sc_hd__or3_1 _15147_ (.A(_07265_),
    .B(_07270_),
    .C(_07710_),
    .X(_07834_));
 sky130_fd_sc_hd__nor2_1 _15148_ (.A(_07049_),
    .B(_07786_),
    .Y(_07835_));
 sky130_fd_sc_hd__or3b_1 _15149_ (.A(_06873_),
    .B(_07332_),
    .C_N(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__o22ai_1 _15150_ (.A1(_07265_),
    .A2(_07332_),
    .B1(_07786_),
    .B2(_06873_),
    .Y(_07837_));
 sky130_fd_sc_hd__nand2_1 _15151_ (.A(_07836_),
    .B(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__nand2_1 _15152_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_07256_),
    .Y(_07839_));
 sky130_fd_sc_hd__nor2_1 _15153_ (.A(_06866_),
    .B(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__xor2_1 _15154_ (.A(_07838_),
    .B(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__and3_1 _15155_ (.A(_07709_),
    .B(_07834_),
    .C(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__a21oi_1 _15156_ (.A1(_07709_),
    .A2(_07834_),
    .B1(_07841_),
    .Y(_07843_));
 sky130_fd_sc_hd__or2_1 _15157_ (.A(_07842_),
    .B(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__a21oi_1 _15158_ (.A1(_07783_),
    .A2(_07789_),
    .B1(_07785_),
    .Y(_07845_));
 sky130_fd_sc_hd__xnor2_1 _15159_ (.A(_07844_),
    .B(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__a21oi_1 _15160_ (.A1(_07724_),
    .A2(_07833_),
    .B1(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__and3_1 _15161_ (.A(_07724_),
    .B(_07833_),
    .C(_07846_),
    .X(_07848_));
 sky130_fd_sc_hd__nor2_1 _15162_ (.A(_07847_),
    .B(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__xnor2_1 _15163_ (.A(_07793_),
    .B(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__a21o_1 _15164_ (.A1(_07712_),
    .A2(_07722_),
    .B1(_07720_),
    .X(_07851_));
 sky130_fd_sc_hd__or2b_1 _15165_ (.A(_07740_),
    .B_N(_07728_),
    .X(_07852_));
 sky130_fd_sc_hd__nor2_1 _15166_ (.A(_06857_),
    .B(_07235_),
    .Y(_07853_));
 sky130_fd_sc_hd__or4_1 _15167_ (.A(_06857_),
    .B(_06875_),
    .C(_07235_),
    .D(_06979_),
    .X(_07854_));
 sky130_fd_sc_hd__o21ai_1 _15168_ (.A1(_07708_),
    .A2(_07853_),
    .B1(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__buf_2 _15169_ (.A(_07007_),
    .X(_07856_));
 sky130_fd_sc_hd__clkbuf_4 _15170_ (.A(_07270_),
    .X(_07857_));
 sky130_fd_sc_hd__nor2_1 _15171_ (.A(_07856_),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__xnor2_1 _15172_ (.A(_07855_),
    .B(_07858_),
    .Y(_07859_));
 sky130_fd_sc_hd__or2_1 _15173_ (.A(_07078_),
    .B(_07039_),
    .X(_07860_));
 sky130_fd_sc_hd__or4_1 _15174_ (.A(_07078_),
    .B(_06900_),
    .C(_07039_),
    .D(_07273_),
    .X(_07861_));
 sky130_fd_sc_hd__a21bo_1 _15175_ (.A1(_07713_),
    .A2(_07860_),
    .B1_N(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__nor2_1 _15176_ (.A(_07084_),
    .B(_07281_),
    .Y(_07863_));
 sky130_fd_sc_hd__xor2_1 _15177_ (.A(_07862_),
    .B(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__clkbuf_4 _15178_ (.A(_07235_),
    .X(_07865_));
 sky130_fd_sc_hd__o31a_1 _15179_ (.A1(_07865_),
    .A2(_07281_),
    .A3(_07716_),
    .B1(_07714_),
    .X(_07866_));
 sky130_fd_sc_hd__nor2_1 _15180_ (.A(_07864_),
    .B(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__nand2_1 _15181_ (.A(_07864_),
    .B(_07866_),
    .Y(_07868_));
 sky130_fd_sc_hd__and2b_1 _15182_ (.A_N(_07867_),
    .B(_07868_),
    .X(_07869_));
 sky130_fd_sc_hd__xnor2_1 _15183_ (.A(_07859_),
    .B(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__a21o_1 _15184_ (.A1(_07738_),
    .A2(_07852_),
    .B1(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__nand3_1 _15185_ (.A(_07738_),
    .B(_07852_),
    .C(_07870_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_1 _15186_ (.A(_07871_),
    .B(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__xnor2_1 _15187_ (.A(_07851_),
    .B(_07873_),
    .Y(_07874_));
 sky130_fd_sc_hd__nand2_1 _15188_ (.A(_07094_),
    .B(_07732_),
    .Y(_07875_));
 sky130_fd_sc_hd__a22o_1 _15189_ (.A1(_07093_),
    .A2(_07733_),
    .B1(_07736_),
    .B2(_07875_),
    .X(_07876_));
 sky130_fd_sc_hd__clkbuf_4 _15190_ (.A(_07100_),
    .X(_07877_));
 sky130_fd_sc_hd__clkbuf_4 _15191_ (.A(_07138_),
    .X(_07878_));
 sky130_fd_sc_hd__o31ai_2 _15192_ (.A1(_07877_),
    .A2(_07878_),
    .A3(_07744_),
    .B1(_07743_),
    .Y(_07879_));
 sky130_fd_sc_hd__nor2_1 _15193_ (.A(_07581_),
    .B(_07138_),
    .Y(_07880_));
 sky130_fd_sc_hd__or3_1 _15194_ (.A(_07530_),
    .B(_07138_),
    .C(_07732_),
    .X(_07881_));
 sky130_fd_sc_hd__o21ai_1 _15195_ (.A1(_07733_),
    .A2(_07880_),
    .B1(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__nor2_1 _15196_ (.A(_06997_),
    .B(_07123_),
    .Y(_07883_));
 sky130_fd_sc_hd__xnor2_1 _15197_ (.A(_07882_),
    .B(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__xnor2_1 _15198_ (.A(_07879_),
    .B(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__xnor2_2 _15199_ (.A(_07876_),
    .B(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__or2_1 _15200_ (.A(_07100_),
    .B(_07137_),
    .X(_07887_));
 sky130_fd_sc_hd__or4_1 _15201_ (.A(_07617_),
    .B(_07646_),
    .C(_07198_),
    .D(_07748_),
    .X(_07888_));
 sky130_fd_sc_hd__o22ai_1 _15202_ (.A1(_07661_),
    .A2(_07766_),
    .B1(_07748_),
    .B2(_07662_),
    .Y(_07889_));
 sky130_fd_sc_hd__nand2_1 _15203_ (.A(_07888_),
    .B(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__xor2_2 _15204_ (.A(_07887_),
    .B(_07890_),
    .X(_07891_));
 sky130_fd_sc_hd__nand2_1 _15205_ (.A(_07673_),
    .B(_07173_),
    .Y(_07892_));
 sky130_fd_sc_hd__nor4_4 _15206_ (.A(_06759_),
    .B(_06764_),
    .C(_06767_),
    .D(_07165_),
    .Y(_07893_));
 sky130_fd_sc_hd__o31a_1 _15207_ (.A1(_06759_),
    .A2(_06764_),
    .A3(_07165_),
    .B1(_06767_),
    .X(_07894_));
 sky130_fd_sc_hd__o31a_1 _15208_ (.A1(_06853_),
    .A2(_07893_),
    .A3(_07894_),
    .B1(_07161_),
    .X(_07895_));
 sky130_fd_sc_hd__a21o_1 _15209_ (.A1(_03492_),
    .A2(\rbzero.wall_tracer.stepDistY[6] ),
    .B1(_04949_),
    .X(_07896_));
 sky130_fd_sc_hd__o22ai_4 _15210_ (.A1(_04841_),
    .A2(\rbzero.wall_tracer.stepDistX[6] ),
    .B1(_07895_),
    .B2(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__or2_1 _15211_ (.A(_07178_),
    .B(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__nor3_1 _15212_ (.A(_07185_),
    .B(_07757_),
    .C(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__nor2_1 _15213_ (.A(_07185_),
    .B(_07897_),
    .Y(_07900_));
 sky130_fd_sc_hd__o21bai_1 _15214_ (.A1(_07199_),
    .A2(_07757_),
    .B1_N(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__and2b_1 _15215_ (.A_N(_07899_),
    .B(_07901_),
    .X(_07902_));
 sky130_fd_sc_hd__xnor2_1 _15216_ (.A(_07892_),
    .B(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__o21a_1 _15217_ (.A1(_07749_),
    .A2(_07759_),
    .B1(_07755_),
    .X(_07904_));
 sky130_fd_sc_hd__xnor2_1 _15218_ (.A(_07903_),
    .B(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__xnor2_2 _15219_ (.A(_07891_),
    .B(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__nor2_1 _15220_ (.A(_07760_),
    .B(_07762_),
    .Y(_07907_));
 sky130_fd_sc_hd__a21oi_2 _15221_ (.A1(_07746_),
    .A2(_07763_),
    .B1(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__xor2_2 _15222_ (.A(_07906_),
    .B(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__xnor2_2 _15223_ (.A(_07886_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__nor2_1 _15224_ (.A(_07764_),
    .B(_07769_),
    .Y(_07911_));
 sky130_fd_sc_hd__a21oi_1 _15225_ (.A1(_07741_),
    .A2(_07770_),
    .B1(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__xor2_1 _15226_ (.A(_07910_),
    .B(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__xnor2_1 _15227_ (.A(_07874_),
    .B(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__a21oi_1 _15228_ (.A1(_07727_),
    .A2(_07774_),
    .B1(_07773_),
    .Y(_07915_));
 sky130_fd_sc_hd__nor2_1 _15229_ (.A(_07914_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_07914_),
    .B(_07915_),
    .Y(_07917_));
 sky130_fd_sc_hd__and2b_1 _15231_ (.A_N(_07916_),
    .B(_07917_),
    .X(_07918_));
 sky130_fd_sc_hd__xnor2_1 _15232_ (.A(_07850_),
    .B(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__a21oi_1 _15233_ (.A1(_07780_),
    .A2(_07798_),
    .B1(_07778_),
    .Y(_07920_));
 sky130_fd_sc_hd__nor2_1 _15234_ (.A(_07919_),
    .B(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__and2_1 _15235_ (.A(_07919_),
    .B(_07920_),
    .X(_07922_));
 sky130_fd_sc_hd__nor2_1 _15236_ (.A(_07921_),
    .B(_07922_),
    .Y(_07923_));
 sky130_fd_sc_hd__xnor2_2 _15237_ (.A(_07796_),
    .B(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__nor2_1 _15238_ (.A(_07799_),
    .B(_07801_),
    .Y(_07925_));
 sky130_fd_sc_hd__a21oi_2 _15239_ (.A1(_07336_),
    .A2(_07802_),
    .B1(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__xor2_2 _15240_ (.A(_07924_),
    .B(_07926_),
    .X(_07927_));
 sky130_fd_sc_hd__xnor2_2 _15241_ (.A(_07832_),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__xnor2_4 _15242_ (.A(_07830_),
    .B(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__mux2_1 _15243_ (.A0(\rbzero.debug_overlay.playerY[-5] ),
    .A1(\rbzero.debug_overlay.playerX[-5] ),
    .S(_06851_),
    .X(_07930_));
 sky130_fd_sc_hd__nand2_1 _15244_ (.A(_07929_),
    .B(_07930_),
    .Y(_07931_));
 sky130_fd_sc_hd__or2_1 _15245_ (.A(_07929_),
    .B(_07930_),
    .X(_07932_));
 sky130_fd_sc_hd__nand2_1 _15246_ (.A(_07931_),
    .B(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__a21o_1 _15247_ (.A1(_07810_),
    .A2(_07822_),
    .B1(_07933_),
    .X(_07934_));
 sky130_fd_sc_hd__nand3_1 _15248_ (.A(_07810_),
    .B(_07822_),
    .C(_07933_),
    .Y(_07935_));
 sky130_fd_sc_hd__inv_2 _15249_ (.A(_06914_),
    .Y(_07936_));
 sky130_fd_sc_hd__mux2_2 _15250_ (.A0(_07936_),
    .A1(_04923_),
    .S(_06851_),
    .X(_07937_));
 sky130_fd_sc_hd__a21oi_1 _15251_ (.A1(_07934_),
    .A2(_07935_),
    .B1(_07937_),
    .Y(_07938_));
 sky130_fd_sc_hd__a31o_1 _15252_ (.A1(_07937_),
    .A2(_07934_),
    .A3(_07935_),
    .B1(_04832_),
    .X(_07939_));
 sky130_fd_sc_hd__o221a_1 _15253_ (.A1(\rbzero.wall_tracer.texu[1] ),
    .A2(_06853_),
    .B1(_07938_),
    .B2(_07939_),
    .C1(_03498_),
    .X(_00476_));
 sky130_fd_sc_hd__nor2_2 _15254_ (.A(_07924_),
    .B(_07926_),
    .Y(_07940_));
 sky130_fd_sc_hd__a31o_2 _15255_ (.A1(_07782_),
    .A2(_07792_),
    .A3(_07849_),
    .B1(_07847_),
    .X(_07941_));
 sky130_fd_sc_hd__or2b_1 _15256_ (.A(_07873_),
    .B_N(_07851_),
    .X(_07942_));
 sky130_fd_sc_hd__o31ai_2 _15257_ (.A1(_07856_),
    .A2(_07270_),
    .A3(_07855_),
    .B1(_07854_),
    .Y(_07943_));
 sky130_fd_sc_hd__or4_1 _15258_ (.A(_07007_),
    .B(_07049_),
    .C(_07332_),
    .D(_07786_),
    .X(_07944_));
 sky130_fd_sc_hd__o21bai_1 _15259_ (.A1(_07007_),
    .A2(_07332_),
    .B1_N(_07835_),
    .Y(_07945_));
 sky130_fd_sc_hd__nand2_1 _15260_ (.A(_07944_),
    .B(_07945_),
    .Y(_07946_));
 sky130_fd_sc_hd__nor2_1 _15261_ (.A(_06873_),
    .B(_07839_),
    .Y(_07947_));
 sky130_fd_sc_hd__xor2_1 _15262_ (.A(_07946_),
    .B(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__xor2_1 _15263_ (.A(_07943_),
    .B(_07948_),
    .X(_07949_));
 sky130_fd_sc_hd__a21bo_1 _15264_ (.A1(_07837_),
    .A2(_07840_),
    .B1_N(_07836_),
    .X(_07950_));
 sky130_fd_sc_hd__or2b_1 _15265_ (.A(_07949_),
    .B_N(_07950_),
    .X(_07951_));
 sky130_fd_sc_hd__or2b_1 _15266_ (.A(_07950_),
    .B_N(_07949_),
    .X(_07952_));
 sky130_fd_sc_hd__nand2_1 _15267_ (.A(_07951_),
    .B(_07952_),
    .Y(_07953_));
 sky130_fd_sc_hd__and2b_1 _15268_ (.A_N(_07842_),
    .B(_07785_),
    .X(_07954_));
 sky130_fd_sc_hd__nor2_1 _15269_ (.A(_07843_),
    .B(_07954_),
    .Y(_07955_));
 sky130_fd_sc_hd__nor2_1 _15270_ (.A(_07953_),
    .B(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__and2_1 _15271_ (.A(_07953_),
    .B(_07955_),
    .X(_07957_));
 sky130_fd_sc_hd__nor2_1 _15272_ (.A(_07956_),
    .B(_07957_),
    .Y(_07958_));
 sky130_fd_sc_hd__nand2_2 _15273_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_07256_),
    .Y(_07959_));
 sky130_fd_sc_hd__buf_2 _15274_ (.A(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__clkbuf_4 _15275_ (.A(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__nor2_1 _15276_ (.A(_07011_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__xnor2_1 _15277_ (.A(_07958_),
    .B(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__a21o_1 _15278_ (.A1(_07871_),
    .A2(_07942_),
    .B1(_07963_),
    .X(_07964_));
 sky130_fd_sc_hd__nand3_1 _15279_ (.A(_07871_),
    .B(_07942_),
    .C(_07963_),
    .Y(_07965_));
 sky130_fd_sc_hd__nand2_1 _15280_ (.A(_07964_),
    .B(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__nor2_1 _15281_ (.A(_07790_),
    .B(_07844_),
    .Y(_07967_));
 sky130_fd_sc_hd__xnor2_1 _15282_ (.A(_07966_),
    .B(_07967_),
    .Y(_07968_));
 sky130_fd_sc_hd__a21o_1 _15283_ (.A1(_07859_),
    .A2(_07868_),
    .B1(_07867_),
    .X(_07969_));
 sky130_fd_sc_hd__or2b_1 _15284_ (.A(_07885_),
    .B_N(_07876_),
    .X(_07970_));
 sky130_fd_sc_hd__a21bo_1 _15285_ (.A1(_07879_),
    .A2(_07884_),
    .B1_N(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__buf_2 _15286_ (.A(_06979_),
    .X(_07972_));
 sky130_fd_sc_hd__nor2_1 _15287_ (.A(_06874_),
    .B(_07084_),
    .Y(_07973_));
 sky130_fd_sc_hd__o22a_1 _15288_ (.A1(_06856_),
    .A2(_07084_),
    .B1(_07235_),
    .B2(_06874_),
    .X(_07974_));
 sky130_fd_sc_hd__a21o_1 _15289_ (.A1(_07853_),
    .A2(_07973_),
    .B1(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__or3_1 _15290_ (.A(_07972_),
    .B(_07270_),
    .C(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__o21ai_1 _15291_ (.A1(_07972_),
    .A2(_07270_),
    .B1(_07975_),
    .Y(_07977_));
 sky130_fd_sc_hd__and2_1 _15292_ (.A(_07976_),
    .B(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__or2_1 _15293_ (.A(_07273_),
    .B(_07092_),
    .X(_07979_));
 sky130_fd_sc_hd__o22a_1 _15294_ (.A1(_07078_),
    .A2(_07273_),
    .B1(_07092_),
    .B2(_07039_),
    .X(_07980_));
 sky130_fd_sc_hd__o21bai_1 _15295_ (.A1(_07860_),
    .A2(_07979_),
    .B1_N(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__or2_1 _15296_ (.A(_07097_),
    .B(_07052_),
    .X(_07982_));
 sky130_fd_sc_hd__xnor2_1 _15297_ (.A(_07981_),
    .B(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__clkbuf_4 _15298_ (.A(_07084_),
    .X(_07984_));
 sky130_fd_sc_hd__o31a_1 _15299_ (.A1(_07984_),
    .A2(_07281_),
    .A3(_07862_),
    .B1(_07861_),
    .X(_07985_));
 sky130_fd_sc_hd__xor2_1 _15300_ (.A(_07983_),
    .B(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__nand2_1 _15301_ (.A(_07978_),
    .B(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__or2_1 _15302_ (.A(_07978_),
    .B(_07986_),
    .X(_07988_));
 sky130_fd_sc_hd__and2_1 _15303_ (.A(_07987_),
    .B(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__xnor2_1 _15304_ (.A(_07971_),
    .B(_07989_),
    .Y(_07990_));
 sky130_fd_sc_hd__xnor2_2 _15305_ (.A(_07969_),
    .B(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__clkbuf_4 _15306_ (.A(_06997_),
    .X(_07992_));
 sky130_fd_sc_hd__clkbuf_4 _15307_ (.A(_07123_),
    .X(_07993_));
 sky130_fd_sc_hd__or3_1 _15308_ (.A(_07992_),
    .B(_07993_),
    .C(_07882_),
    .X(_07994_));
 sky130_fd_sc_hd__o21ai_1 _15309_ (.A1(_07887_),
    .A2(_07890_),
    .B1(_07888_),
    .Y(_07995_));
 sky130_fd_sc_hd__o22a_1 _15310_ (.A1(_07530_),
    .A2(_07138_),
    .B1(_07137_),
    .B2(_07581_),
    .X(_07996_));
 sky130_fd_sc_hd__nor2_1 _15311_ (.A(_07530_),
    .B(_07137_),
    .Y(_07997_));
 sky130_fd_sc_hd__and2_1 _15312_ (.A(_07880_),
    .B(_07997_),
    .X(_07998_));
 sky130_fd_sc_hd__nor2_1 _15313_ (.A(_07996_),
    .B(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__clkbuf_4 _15314_ (.A(_07141_),
    .X(_08000_));
 sky130_fd_sc_hd__nor2_1 _15315_ (.A(_06997_),
    .B(_08000_),
    .Y(_08001_));
 sky130_fd_sc_hd__xnor2_1 _15316_ (.A(_07999_),
    .B(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__xor2_1 _15317_ (.A(_07995_),
    .B(_08002_),
    .X(_08003_));
 sky130_fd_sc_hd__a21o_1 _15318_ (.A1(_07881_),
    .A2(_07994_),
    .B1(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__nand3_1 _15319_ (.A(_07881_),
    .B(_07994_),
    .C(_08003_),
    .Y(_08005_));
 sky130_fd_sc_hd__and2_1 _15320_ (.A(_08004_),
    .B(_08005_),
    .X(_08006_));
 sky130_fd_sc_hd__or2_1 _15321_ (.A(_07877_),
    .B(_07766_),
    .X(_08007_));
 sky130_fd_sc_hd__or4_1 _15322_ (.A(_07617_),
    .B(_07646_),
    .C(_07748_),
    .D(_07756_),
    .X(_08008_));
 sky130_fd_sc_hd__o22ai_1 _15323_ (.A1(_07617_),
    .A2(_07748_),
    .B1(_07756_),
    .B2(_07646_),
    .Y(_08009_));
 sky130_fd_sc_hd__and2_1 _15324_ (.A(_08008_),
    .B(_08009_),
    .X(_08010_));
 sky130_fd_sc_hd__xnor2_1 _15325_ (.A(_08007_),
    .B(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__or2_1 _15326_ (.A(_07213_),
    .B(_07757_),
    .X(_08012_));
 sky130_fd_sc_hd__or2_1 _15327_ (.A(_06771_),
    .B(_07893_),
    .X(_08013_));
 sky130_fd_sc_hd__nand2_1 _15328_ (.A(_06771_),
    .B(_07893_),
    .Y(_08014_));
 sky130_fd_sc_hd__a31o_1 _15329_ (.A1(_04832_),
    .A2(_08013_),
    .A3(_08014_),
    .B1(_07162_),
    .X(_08015_));
 sky130_fd_sc_hd__a21oi_1 _15330_ (.A1(_03493_),
    .A2(\rbzero.wall_tracer.stepDistY[7] ),
    .B1(_04950_),
    .Y(_08016_));
 sky130_fd_sc_hd__nor2_1 _15331_ (.A(_04841_),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_08017_));
 sky130_fd_sc_hd__a21o_4 _15332_ (.A1(_08015_),
    .A2(_08016_),
    .B1(_08017_),
    .X(_08018_));
 sky130_fd_sc_hd__nor2_1 _15333_ (.A(_07199_),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__or4_1 _15334_ (.A(_07175_),
    .B(_04950_),
    .C(_03493_),
    .D(_08015_),
    .X(_08020_));
 sky130_fd_sc_hd__and2_1 _15335_ (.A(_07898_),
    .B(_08020_),
    .X(_08021_));
 sky130_fd_sc_hd__a21oi_1 _15336_ (.A1(_07900_),
    .A2(_08019_),
    .B1(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__xnor2_1 _15337_ (.A(_08012_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__a31oi_1 _15338_ (.A1(_07673_),
    .A2(_07173_),
    .A3(_07901_),
    .B1(_07899_),
    .Y(_08024_));
 sky130_fd_sc_hd__xnor2_1 _15339_ (.A(_08023_),
    .B(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__nand2_1 _15340_ (.A(_08011_),
    .B(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__or2_1 _15341_ (.A(_08011_),
    .B(_08025_),
    .X(_08027_));
 sky130_fd_sc_hd__nand2_1 _15342_ (.A(_08026_),
    .B(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__and2b_1 _15343_ (.A_N(_07904_),
    .B(_07903_),
    .X(_08029_));
 sky130_fd_sc_hd__a21o_1 _15344_ (.A1(_07891_),
    .A2(_07905_),
    .B1(_08029_),
    .X(_08030_));
 sky130_fd_sc_hd__xnor2_2 _15345_ (.A(_08028_),
    .B(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__xnor2_2 _15346_ (.A(_08006_),
    .B(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__nor2_1 _15347_ (.A(_07906_),
    .B(_07908_),
    .Y(_08033_));
 sky130_fd_sc_hd__a21oi_1 _15348_ (.A1(_07886_),
    .A2(_07909_),
    .B1(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__xor2_2 _15349_ (.A(_08032_),
    .B(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__xnor2_2 _15350_ (.A(_07991_),
    .B(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__nor2_1 _15351_ (.A(_07910_),
    .B(_07912_),
    .Y(_08037_));
 sky130_fd_sc_hd__a21oi_1 _15352_ (.A1(_07874_),
    .A2(_07913_),
    .B1(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__xor2_1 _15353_ (.A(_08036_),
    .B(_08038_),
    .X(_08039_));
 sky130_fd_sc_hd__xnor2_1 _15354_ (.A(_07968_),
    .B(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__a21oi_1 _15355_ (.A1(_07850_),
    .A2(_07917_),
    .B1(_07916_),
    .Y(_08041_));
 sky130_fd_sc_hd__nor2_1 _15356_ (.A(_08040_),
    .B(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__and2_1 _15357_ (.A(_08040_),
    .B(_08041_),
    .X(_08043_));
 sky130_fd_sc_hd__nor2_2 _15358_ (.A(_08042_),
    .B(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__xnor2_4 _15359_ (.A(_07941_),
    .B(_08044_),
    .Y(_08045_));
 sky130_fd_sc_hd__a21oi_2 _15360_ (.A1(_07796_),
    .A2(_07923_),
    .B1(_07921_),
    .Y(_08046_));
 sky130_fd_sc_hd__xor2_4 _15361_ (.A(_08045_),
    .B(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__xor2_4 _15362_ (.A(_07940_),
    .B(_08047_),
    .X(_08048_));
 sky130_fd_sc_hd__inv_2 _15363_ (.A(_07927_),
    .Y(_08049_));
 sky130_fd_sc_hd__a21oi_1 _15364_ (.A1(_07703_),
    .A2(_07807_),
    .B1(_07927_),
    .Y(_08050_));
 sky130_fd_sc_hd__o22a_2 _15365_ (.A1(_07832_),
    .A2(_08049_),
    .B1(_08050_),
    .B2(_07830_),
    .X(_08051_));
 sky130_fd_sc_hd__xnor2_4 _15366_ (.A(_08048_),
    .B(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__mux2_1 _15367_ (.A0(\rbzero.debug_overlay.playerY[-4] ),
    .A1(\rbzero.debug_overlay.playerX[-4] ),
    .S(_06851_),
    .X(_08053_));
 sky130_fd_sc_hd__nand2_1 _15368_ (.A(_08052_),
    .B(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__or2_1 _15369_ (.A(_08052_),
    .B(_08053_),
    .X(_08055_));
 sky130_fd_sc_hd__nand2_1 _15370_ (.A(_08054_),
    .B(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__a21o_1 _15371_ (.A1(_07931_),
    .A2(_07934_),
    .B1(_08056_),
    .X(_08057_));
 sky130_fd_sc_hd__nand3_1 _15372_ (.A(_07931_),
    .B(_07934_),
    .C(_08056_),
    .Y(_08058_));
 sky130_fd_sc_hd__a21oi_1 _15373_ (.A1(_08057_),
    .A2(_08058_),
    .B1(_07937_),
    .Y(_08059_));
 sky130_fd_sc_hd__a31o_1 _15374_ (.A1(_07937_),
    .A2(_08057_),
    .A3(_08058_),
    .B1(_04832_),
    .X(_08060_));
 sky130_fd_sc_hd__o221a_1 _15375_ (.A1(\rbzero.wall_tracer.texu[2] ),
    .A2(_06853_),
    .B1(_08059_),
    .B2(_08060_),
    .C1(_03498_),
    .X(_00477_));
 sky130_fd_sc_hd__nor2_1 _15376_ (.A(_07940_),
    .B(_08047_),
    .Y(_08061_));
 sky130_fd_sc_hd__nand2_1 _15377_ (.A(_07940_),
    .B(_08047_),
    .Y(_08062_));
 sky130_fd_sc_hd__o21ai_2 _15378_ (.A1(_08061_),
    .A2(_08051_),
    .B1(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__or2_1 _15379_ (.A(_08045_),
    .B(_08046_),
    .X(_08064_));
 sky130_fd_sc_hd__o31ai_2 _15380_ (.A1(_07790_),
    .A2(_07844_),
    .A3(_07966_),
    .B1(_07964_),
    .Y(_08065_));
 sky130_fd_sc_hd__a21o_1 _15381_ (.A1(_07958_),
    .A2(_07962_),
    .B1(_07956_),
    .X(_08066_));
 sky130_fd_sc_hd__or2b_1 _15382_ (.A(_07990_),
    .B_N(_07969_),
    .X(_08067_));
 sky130_fd_sc_hd__a21bo_1 _15383_ (.A1(_07971_),
    .A2(_07989_),
    .B1_N(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__nand2_1 _15384_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_07256_),
    .Y(_08069_));
 sky130_fd_sc_hd__buf_2 _15385_ (.A(_08069_),
    .X(_08070_));
 sky130_fd_sc_hd__clkbuf_4 _15386_ (.A(_08070_),
    .X(_08071_));
 sky130_fd_sc_hd__nor4_1 _15387_ (.A(_07011_),
    .B(_07269_),
    .C(_07961_),
    .D(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__o22a_1 _15388_ (.A1(_07269_),
    .A2(_07961_),
    .B1(_08071_),
    .B2(_07011_),
    .X(_08073_));
 sky130_fd_sc_hd__nor2_1 _15389_ (.A(_08072_),
    .B(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__a21bo_1 _15390_ (.A1(_07945_),
    .A2(_07947_),
    .B1_N(_07944_),
    .X(_08075_));
 sky130_fd_sc_hd__nand2_1 _15391_ (.A(_07853_),
    .B(_07973_),
    .Y(_08076_));
 sky130_fd_sc_hd__nor2_1 _15392_ (.A(_07856_),
    .B(_07787_),
    .Y(_08077_));
 sky130_fd_sc_hd__nor2_1 _15393_ (.A(_06979_),
    .B(_07332_),
    .Y(_08078_));
 sky130_fd_sc_hd__or4_1 _15394_ (.A(_06979_),
    .B(_07007_),
    .C(_07332_),
    .D(_07786_),
    .X(_08079_));
 sky130_fd_sc_hd__o21a_1 _15395_ (.A1(_08077_),
    .A2(_08078_),
    .B1(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__clkbuf_4 _15396_ (.A(_07839_),
    .X(_08081_));
 sky130_fd_sc_hd__nor2_1 _15397_ (.A(_07265_),
    .B(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__xnor2_1 _15398_ (.A(_08080_),
    .B(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__a21oi_1 _15399_ (.A1(_08076_),
    .A2(_07976_),
    .B1(_08083_),
    .Y(_08084_));
 sky130_fd_sc_hd__and3_1 _15400_ (.A(_08076_),
    .B(_07976_),
    .C(_08083_),
    .X(_08085_));
 sky130_fd_sc_hd__nor2_1 _15401_ (.A(_08084_),
    .B(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__xnor2_1 _15402_ (.A(_08075_),
    .B(_08086_),
    .Y(_08087_));
 sky130_fd_sc_hd__inv_2 _15403_ (.A(_07943_),
    .Y(_08088_));
 sky130_fd_sc_hd__o21a_1 _15404_ (.A1(_08088_),
    .A2(_07948_),
    .B1(_07951_),
    .X(_08089_));
 sky130_fd_sc_hd__xor2_1 _15405_ (.A(_08087_),
    .B(_08089_),
    .X(_08090_));
 sky130_fd_sc_hd__xor2_1 _15406_ (.A(_08074_),
    .B(_08090_),
    .X(_08091_));
 sky130_fd_sc_hd__xnor2_1 _15407_ (.A(_08068_),
    .B(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__xnor2_2 _15408_ (.A(_08066_),
    .B(_08092_),
    .Y(_08093_));
 sky130_fd_sc_hd__o21ai_1 _15409_ (.A1(_07983_),
    .A2(_07985_),
    .B1(_07987_),
    .Y(_08094_));
 sky130_fd_sc_hd__or2b_1 _15410_ (.A(_08002_),
    .B_N(_07995_),
    .X(_08095_));
 sky130_fd_sc_hd__nand2_1 _15411_ (.A(_08095_),
    .B(_08004_),
    .Y(_08096_));
 sky130_fd_sc_hd__nor2_1 _15412_ (.A(_06858_),
    .B(_07097_),
    .Y(_08097_));
 sky130_fd_sc_hd__or4_1 _15413_ (.A(_06857_),
    .B(_06875_),
    .C(_07097_),
    .D(_07084_),
    .X(_08098_));
 sky130_fd_sc_hd__o21ai_1 _15414_ (.A1(_07973_),
    .A2(_08097_),
    .B1(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__nor2_1 _15415_ (.A(_07865_),
    .B(_07857_),
    .Y(_08100_));
 sky130_fd_sc_hd__xnor2_1 _15416_ (.A(_08099_),
    .B(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__or2_1 _15417_ (.A(_07039_),
    .B(_07141_),
    .X(_08102_));
 sky130_fd_sc_hd__or4_1 _15418_ (.A(_07039_),
    .B(_07273_),
    .C(_07141_),
    .D(_07092_),
    .X(_08103_));
 sky130_fd_sc_hd__a21bo_1 _15419_ (.A1(_07979_),
    .A2(_08102_),
    .B1_N(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__or2_1 _15420_ (.A(_07735_),
    .B(_07281_),
    .X(_08105_));
 sky130_fd_sc_hd__xnor2_1 _15421_ (.A(_08104_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__clkbuf_4 _15422_ (.A(_07097_),
    .X(_08107_));
 sky130_fd_sc_hd__buf_2 _15423_ (.A(_07281_),
    .X(_08108_));
 sky130_fd_sc_hd__o32a_1 _15424_ (.A1(_08107_),
    .A2(_08108_),
    .A3(_07980_),
    .B1(_07979_),
    .B2(_07860_),
    .X(_08109_));
 sky130_fd_sc_hd__nor2_1 _15425_ (.A(_08106_),
    .B(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__and2_1 _15426_ (.A(_08106_),
    .B(_08109_),
    .X(_08111_));
 sky130_fd_sc_hd__nor2_1 _15427_ (.A(_08110_),
    .B(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__xor2_1 _15428_ (.A(_08101_),
    .B(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__xnor2_1 _15429_ (.A(_08096_),
    .B(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__xnor2_2 _15430_ (.A(_08094_),
    .B(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__a21o_1 _15431_ (.A1(_07999_),
    .A2(_08001_),
    .B1(_07998_),
    .X(_08116_));
 sky130_fd_sc_hd__or2b_1 _15432_ (.A(_08007_),
    .B_N(_08010_),
    .X(_08117_));
 sky130_fd_sc_hd__nor2_1 _15433_ (.A(_07581_),
    .B(_07198_),
    .Y(_08118_));
 sky130_fd_sc_hd__or4_1 _15434_ (.A(_06968_),
    .B(_06970_),
    .C(_07137_),
    .D(_07198_),
    .X(_08119_));
 sky130_fd_sc_hd__o21a_1 _15435_ (.A1(_07997_),
    .A2(_08118_),
    .B1(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__nor2_1 _15436_ (.A(_06997_),
    .B(_07138_),
    .Y(_08121_));
 sky130_fd_sc_hd__nand2_1 _15437_ (.A(_08120_),
    .B(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__or2_1 _15438_ (.A(_08120_),
    .B(_08121_),
    .X(_08123_));
 sky130_fd_sc_hd__nand2_1 _15439_ (.A(_08122_),
    .B(_08123_),
    .Y(_08124_));
 sky130_fd_sc_hd__a21o_1 _15440_ (.A1(_08008_),
    .A2(_08117_),
    .B1(_08124_),
    .X(_08125_));
 sky130_fd_sc_hd__nand3_1 _15441_ (.A(_08008_),
    .B(_08117_),
    .C(_08124_),
    .Y(_08126_));
 sky130_fd_sc_hd__and2_1 _15442_ (.A(_08125_),
    .B(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__xor2_1 _15443_ (.A(_08116_),
    .B(_08127_),
    .X(_08128_));
 sky130_fd_sc_hd__or2b_1 _15444_ (.A(_08024_),
    .B_N(_08023_),
    .X(_08129_));
 sky130_fd_sc_hd__buf_2 _15445_ (.A(_07748_),
    .X(_08130_));
 sky130_fd_sc_hd__nor2_1 _15446_ (.A(_07877_),
    .B(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__or4_1 _15447_ (.A(_07617_),
    .B(_07646_),
    .C(_07756_),
    .D(_07757_),
    .X(_08132_));
 sky130_fd_sc_hd__buf_2 _15448_ (.A(_07756_),
    .X(_08133_));
 sky130_fd_sc_hd__buf_2 _15449_ (.A(_07757_),
    .X(_08134_));
 sky130_fd_sc_hd__o22ai_1 _15450_ (.A1(_07661_),
    .A2(_08133_),
    .B1(_08134_),
    .B2(_07662_),
    .Y(_08135_));
 sky130_fd_sc_hd__nand2_1 _15451_ (.A(_08132_),
    .B(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__xnor2_1 _15452_ (.A(_08131_),
    .B(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__nor2_1 _15453_ (.A(_07213_),
    .B(_07897_),
    .Y(_08138_));
 sky130_fd_sc_hd__a21boi_1 _15454_ (.A1(_06771_),
    .A2(_07893_),
    .B1_N(_06777_),
    .Y(_08139_));
 sky130_fd_sc_hd__a31o_1 _15455_ (.A1(_06771_),
    .A2(_06776_),
    .A3(_07893_),
    .B1(_06853_),
    .X(_08140_));
 sky130_fd_sc_hd__o21ai_2 _15456_ (.A1(_08139_),
    .A2(_08140_),
    .B1(_07161_),
    .Y(_08141_));
 sky130_fd_sc_hd__or4_2 _15457_ (.A(_07195_),
    .B(_04949_),
    .C(_03493_),
    .D(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__or2_1 _15458_ (.A(_08020_),
    .B(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__a21oi_2 _15459_ (.A1(_08015_),
    .A2(_08016_),
    .B1(_08017_),
    .Y(_08144_));
 sky130_fd_sc_hd__and4bb_1 _15460_ (.A_N(_04950_),
    .B_N(_08141_),
    .C(_06860_),
    .D(_06787_),
    .X(_08145_));
 sky130_fd_sc_hd__a21o_1 _15461_ (.A1(_07174_),
    .A2(_08144_),
    .B1(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__and3_1 _15462_ (.A(_08138_),
    .B(_08143_),
    .C(_08146_),
    .X(_08147_));
 sky130_fd_sc_hd__a21oi_1 _15463_ (.A1(_08143_),
    .A2(_08146_),
    .B1(_08138_),
    .Y(_08148_));
 sky130_fd_sc_hd__o2bb2a_1 _15464_ (.A1_N(_07900_),
    .A2_N(_08019_),
    .B1(_08021_),
    .B2(_08012_),
    .X(_08149_));
 sky130_fd_sc_hd__or3_1 _15465_ (.A(_08147_),
    .B(_08148_),
    .C(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__o21ai_1 _15466_ (.A1(_08147_),
    .A2(_08148_),
    .B1(_08149_),
    .Y(_08151_));
 sky130_fd_sc_hd__nand2_1 _15467_ (.A(_08150_),
    .B(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__xor2_1 _15468_ (.A(_08137_),
    .B(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__a21oi_1 _15469_ (.A1(_08129_),
    .A2(_08026_),
    .B1(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__and3_1 _15470_ (.A(_08129_),
    .B(_08026_),
    .C(_08153_),
    .X(_08155_));
 sky130_fd_sc_hd__nor2_1 _15471_ (.A(_08154_),
    .B(_08155_),
    .Y(_08156_));
 sky130_fd_sc_hd__xnor2_1 _15472_ (.A(_08128_),
    .B(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__a32oi_2 _15473_ (.A1(_08026_),
    .A2(_08027_),
    .A3(_08030_),
    .B1(_08031_),
    .B2(_08006_),
    .Y(_08158_));
 sky130_fd_sc_hd__nor2_1 _15474_ (.A(_08157_),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__and2_1 _15475_ (.A(_08157_),
    .B(_08158_),
    .X(_08160_));
 sky130_fd_sc_hd__nor2_1 _15476_ (.A(_08159_),
    .B(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__xnor2_2 _15477_ (.A(_08115_),
    .B(_08161_),
    .Y(_08162_));
 sky130_fd_sc_hd__nor2_1 _15478_ (.A(_08032_),
    .B(_08034_),
    .Y(_08163_));
 sky130_fd_sc_hd__a21oi_2 _15479_ (.A1(_07991_),
    .A2(_08035_),
    .B1(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__xor2_2 _15480_ (.A(_08162_),
    .B(_08164_),
    .X(_08165_));
 sky130_fd_sc_hd__xnor2_2 _15481_ (.A(_08093_),
    .B(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__nor2_1 _15482_ (.A(_08036_),
    .B(_08038_),
    .Y(_08167_));
 sky130_fd_sc_hd__a21oi_2 _15483_ (.A1(_07968_),
    .A2(_08039_),
    .B1(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__xor2_2 _15484_ (.A(_08166_),
    .B(_08168_),
    .X(_08169_));
 sky130_fd_sc_hd__xnor2_2 _15485_ (.A(_08065_),
    .B(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__a21oi_2 _15486_ (.A1(_07941_),
    .A2(_08044_),
    .B1(_08042_),
    .Y(_08171_));
 sky130_fd_sc_hd__xor2_2 _15487_ (.A(_08170_),
    .B(_08171_),
    .X(_08172_));
 sky130_fd_sc_hd__xnor2_2 _15488_ (.A(_08064_),
    .B(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__xor2_4 _15489_ (.A(_08063_),
    .B(_08173_),
    .X(_08174_));
 sky130_fd_sc_hd__mux2_1 _15490_ (.A0(\rbzero.debug_overlay.playerY[-3] ),
    .A1(\rbzero.debug_overlay.playerX[-3] ),
    .S(_06851_),
    .X(_08175_));
 sky130_fd_sc_hd__xnor2_1 _15491_ (.A(_08174_),
    .B(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__a21oi_1 _15492_ (.A1(_08054_),
    .A2(_08057_),
    .B1(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__and3_1 _15493_ (.A(_08054_),
    .B(_08057_),
    .C(_08176_),
    .X(_08178_));
 sky130_fd_sc_hd__or2_1 _15494_ (.A(_08177_),
    .B(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__nor2_1 _15495_ (.A(_07827_),
    .B(_08179_),
    .Y(_08180_));
 sky130_fd_sc_hd__a21o_1 _15496_ (.A1(_07827_),
    .A2(_08179_),
    .B1(_04832_),
    .X(_08181_));
 sky130_fd_sc_hd__o221a_1 _15497_ (.A1(\rbzero.wall_tracer.texu[3] ),
    .A2(_06853_),
    .B1(_08180_),
    .B2(_08181_),
    .C1(_03498_),
    .X(_00478_));
 sky130_fd_sc_hd__a21oi_1 _15498_ (.A1(_08174_),
    .A2(_08175_),
    .B1(_08177_),
    .Y(_08182_));
 sky130_fd_sc_hd__nor2_1 _15499_ (.A(_08170_),
    .B(_08171_),
    .Y(_08183_));
 sky130_fd_sc_hd__nor2_1 _15500_ (.A(_08166_),
    .B(_08168_),
    .Y(_08184_));
 sky130_fd_sc_hd__a21o_1 _15501_ (.A1(_08065_),
    .A2(_08169_),
    .B1(_08184_),
    .X(_08185_));
 sky130_fd_sc_hd__or2b_1 _15502_ (.A(_08092_),
    .B_N(_08066_),
    .X(_08186_));
 sky130_fd_sc_hd__a21bo_1 _15503_ (.A1(_08068_),
    .A2(_08091_),
    .B1_N(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__a2bb2o_1 _15504_ (.A1_N(_08087_),
    .A2_N(_08089_),
    .B1(_08090_),
    .B2(_08074_),
    .X(_08188_));
 sky130_fd_sc_hd__or2b_1 _15505_ (.A(_08114_),
    .B_N(_08094_),
    .X(_08189_));
 sky130_fd_sc_hd__a21bo_1 _15506_ (.A1(_08096_),
    .A2(_08113_),
    .B1_N(_08189_),
    .X(_08190_));
 sky130_fd_sc_hd__nand2_4 _15507_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_07256_),
    .Y(_08191_));
 sky130_fd_sc_hd__or2_1 _15508_ (.A(_07011_),
    .B(_08191_),
    .X(_08192_));
 sky130_fd_sc_hd__nor2_1 _15509_ (.A(_07265_),
    .B(_08069_),
    .Y(_08193_));
 sky130_fd_sc_hd__or3b_1 _15510_ (.A(_07269_),
    .B(_07959_),
    .C_N(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__inv_2 _15511_ (.A(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__o22a_1 _15512_ (.A1(_07265_),
    .A2(_07960_),
    .B1(_08070_),
    .B2(_07269_),
    .X(_08196_));
 sky130_fd_sc_hd__nor2_1 _15513_ (.A(_08195_),
    .B(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__xnor2_1 _15514_ (.A(_08192_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__nand2_1 _15515_ (.A(_08072_),
    .B(_08198_),
    .Y(_08199_));
 sky130_fd_sc_hd__or2_1 _15516_ (.A(_08072_),
    .B(_08198_),
    .X(_08200_));
 sky130_fd_sc_hd__and2_1 _15517_ (.A(_08199_),
    .B(_08200_),
    .X(_08201_));
 sky130_fd_sc_hd__a21bo_1 _15518_ (.A1(_08080_),
    .A2(_08082_),
    .B1_N(_08079_),
    .X(_08202_));
 sky130_fd_sc_hd__o31a_1 _15519_ (.A1(_07865_),
    .A2(_07857_),
    .A3(_08099_),
    .B1(_08098_),
    .X(_08203_));
 sky130_fd_sc_hd__nor2_1 _15520_ (.A(_07972_),
    .B(_07787_),
    .Y(_08204_));
 sky130_fd_sc_hd__nor2_1 _15521_ (.A(_07235_),
    .B(_07333_),
    .Y(_08205_));
 sky130_fd_sc_hd__nor2_1 _15522_ (.A(_07235_),
    .B(_07786_),
    .Y(_08206_));
 sky130_fd_sc_hd__nand2_1 _15523_ (.A(_08078_),
    .B(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__o21ai_1 _15524_ (.A1(_08204_),
    .A2(_08205_),
    .B1(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__nor2_1 _15525_ (.A(_07856_),
    .B(_08081_),
    .Y(_08209_));
 sky130_fd_sc_hd__xnor2_1 _15526_ (.A(_08208_),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__and2b_1 _15527_ (.A_N(_08203_),
    .B(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__and2b_1 _15528_ (.A_N(_08210_),
    .B(_08203_),
    .X(_08212_));
 sky130_fd_sc_hd__nor2_1 _15529_ (.A(_08211_),
    .B(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__xnor2_1 _15530_ (.A(_08202_),
    .B(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__a21oi_1 _15531_ (.A1(_08075_),
    .A2(_08086_),
    .B1(_08084_),
    .Y(_08215_));
 sky130_fd_sc_hd__nor2_1 _15532_ (.A(_08214_),
    .B(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__and2_1 _15533_ (.A(_08214_),
    .B(_08215_),
    .X(_08217_));
 sky130_fd_sc_hd__nor2_1 _15534_ (.A(_08216_),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__xor2_1 _15535_ (.A(_08201_),
    .B(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__xnor2_1 _15536_ (.A(_08190_),
    .B(_08219_),
    .Y(_08220_));
 sky130_fd_sc_hd__xnor2_1 _15537_ (.A(_08188_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__a21o_1 _15538_ (.A1(_08101_),
    .A2(_08112_),
    .B1(_08110_),
    .X(_08222_));
 sky130_fd_sc_hd__nand2_1 _15539_ (.A(_08116_),
    .B(_08127_),
    .Y(_08223_));
 sky130_fd_sc_hd__nor2_1 _15540_ (.A(_06875_),
    .B(_07735_),
    .Y(_08224_));
 sky130_fd_sc_hd__o22a_1 _15541_ (.A1(_06858_),
    .A2(_07735_),
    .B1(_07097_),
    .B2(_06875_),
    .X(_08225_));
 sky130_fd_sc_hd__a21o_1 _15542_ (.A1(_08097_),
    .A2(_08224_),
    .B1(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__nor2_1 _15543_ (.A(_07984_),
    .B(_07857_),
    .Y(_08227_));
 sky130_fd_sc_hd__xnor2_1 _15544_ (.A(_08226_),
    .B(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__buf_2 _15545_ (.A(_07273_),
    .X(_08229_));
 sky130_fd_sc_hd__or3_1 _15546_ (.A(_08229_),
    .B(_07138_),
    .C(_08102_),
    .X(_08230_));
 sky130_fd_sc_hd__o22ai_1 _15547_ (.A1(_07494_),
    .A2(_07138_),
    .B1(_08000_),
    .B2(_08229_),
    .Y(_08231_));
 sky130_fd_sc_hd__nand2_1 _15548_ (.A(_08230_),
    .B(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__or2_1 _15549_ (.A(_07281_),
    .B(_07123_),
    .X(_08233_));
 sky130_fd_sc_hd__xnor2_1 _15550_ (.A(_08232_),
    .B(_08233_),
    .Y(_08234_));
 sky130_fd_sc_hd__o31a_1 _15551_ (.A1(_07735_),
    .A2(_08108_),
    .A3(_08104_),
    .B1(_08103_),
    .X(_08235_));
 sky130_fd_sc_hd__nor2_1 _15552_ (.A(_08234_),
    .B(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__and2_1 _15553_ (.A(_08234_),
    .B(_08235_),
    .X(_08237_));
 sky130_fd_sc_hd__nor2_1 _15554_ (.A(_08236_),
    .B(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__xnor2_1 _15555_ (.A(_08228_),
    .B(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__a21o_1 _15556_ (.A1(_08125_),
    .A2(_08223_),
    .B1(_08239_),
    .X(_08240_));
 sky130_fd_sc_hd__nand3_1 _15557_ (.A(_08125_),
    .B(_08223_),
    .C(_08239_),
    .Y(_08241_));
 sky130_fd_sc_hd__nand2_1 _15558_ (.A(_08240_),
    .B(_08241_),
    .Y(_08242_));
 sky130_fd_sc_hd__xnor2_1 _15559_ (.A(_08222_),
    .B(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__a21bo_1 _15560_ (.A1(_08131_),
    .A2(_08135_),
    .B1_N(_08132_),
    .X(_08244_));
 sky130_fd_sc_hd__buf_2 _15561_ (.A(_07530_),
    .X(_08245_));
 sky130_fd_sc_hd__nor2_1 _15562_ (.A(_08245_),
    .B(_07766_),
    .Y(_08246_));
 sky130_fd_sc_hd__buf_2 _15563_ (.A(_07581_),
    .X(_08247_));
 sky130_fd_sc_hd__nor2_1 _15564_ (.A(_08247_),
    .B(_08130_),
    .Y(_08248_));
 sky130_fd_sc_hd__or2_1 _15565_ (.A(_06970_),
    .B(_07748_),
    .X(_08249_));
 sky130_fd_sc_hd__or3_1 _15566_ (.A(_07581_),
    .B(_07198_),
    .C(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__o21ai_1 _15567_ (.A1(_08246_),
    .A2(_08248_),
    .B1(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__buf_2 _15568_ (.A(_07137_),
    .X(_08252_));
 sky130_fd_sc_hd__nor2_1 _15569_ (.A(_06997_),
    .B(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__xnor2_1 _15570_ (.A(_08251_),
    .B(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__xnor2_1 _15571_ (.A(_08244_),
    .B(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__a21o_1 _15572_ (.A1(_08119_),
    .A2(_08122_),
    .B1(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__nand3_1 _15573_ (.A(_08119_),
    .B(_08122_),
    .C(_08255_),
    .Y(_08257_));
 sky130_fd_sc_hd__and2_1 _15574_ (.A(_08256_),
    .B(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__or4_1 _15575_ (.A(_07617_),
    .B(_07646_),
    .C(_07757_),
    .D(_07897_),
    .X(_08259_));
 sky130_fd_sc_hd__buf_2 _15576_ (.A(_07897_),
    .X(_08260_));
 sky130_fd_sc_hd__o22ai_1 _15577_ (.A1(_07661_),
    .A2(_08134_),
    .B1(_08260_),
    .B2(_07662_),
    .Y(_08261_));
 sky130_fd_sc_hd__nand2_1 _15578_ (.A(_08259_),
    .B(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__nor2_1 _15579_ (.A(_07877_),
    .B(_08133_),
    .Y(_08263_));
 sky130_fd_sc_hd__xnor2_1 _15580_ (.A(_08262_),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__nand2_1 _15581_ (.A(_07673_),
    .B(_08144_),
    .Y(_08265_));
 sky130_fd_sc_hd__inv_2 _15582_ (.A(_06779_),
    .Y(_08266_));
 sky130_fd_sc_hd__nand4_1 _15583_ (.A(_06771_),
    .B(_06776_),
    .C(_08266_),
    .D(_07893_),
    .Y(_08267_));
 sky130_fd_sc_hd__a31o_1 _15584_ (.A1(_06771_),
    .A2(_06776_),
    .A3(_07893_),
    .B1(_08266_),
    .X(_08268_));
 sky130_fd_sc_hd__a31o_1 _15585_ (.A1(_04832_),
    .A2(_08267_),
    .A3(_08268_),
    .B1(_07162_),
    .X(_08269_));
 sky130_fd_sc_hd__and4bb_2 _15586_ (.A_N(_04950_),
    .B_N(_08269_),
    .C(_06860_),
    .D(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_08270_));
 sky130_fd_sc_hd__or4_1 _15587_ (.A(_07175_),
    .B(_04950_),
    .C(_03493_),
    .D(_08269_),
    .X(_08271_));
 sky130_fd_sc_hd__a22oi_2 _15588_ (.A1(_08145_),
    .A2(_08270_),
    .B1(_08271_),
    .B2(_08142_),
    .Y(_08272_));
 sky130_fd_sc_hd__xnor2_1 _15589_ (.A(_08265_),
    .B(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__a21bo_1 _15590_ (.A1(_08138_),
    .A2(_08146_),
    .B1_N(_08143_),
    .X(_08274_));
 sky130_fd_sc_hd__xor2_1 _15591_ (.A(_08273_),
    .B(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__xnor2_1 _15592_ (.A(_08264_),
    .B(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__a21boi_1 _15593_ (.A1(_08137_),
    .A2(_08151_),
    .B1_N(_08150_),
    .Y(_08277_));
 sky130_fd_sc_hd__nor2_1 _15594_ (.A(_08276_),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__and2_1 _15595_ (.A(_08276_),
    .B(_08277_),
    .X(_08279_));
 sky130_fd_sc_hd__nor2_1 _15596_ (.A(_08278_),
    .B(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__xnor2_2 _15597_ (.A(_08258_),
    .B(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__a21oi_2 _15598_ (.A1(_08128_),
    .A2(_08156_),
    .B1(_08154_),
    .Y(_08282_));
 sky130_fd_sc_hd__xor2_1 _15599_ (.A(_08281_),
    .B(_08282_),
    .X(_08283_));
 sky130_fd_sc_hd__nand2_1 _15600_ (.A(_08243_),
    .B(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__or2_1 _15601_ (.A(_08243_),
    .B(_08283_),
    .X(_08285_));
 sky130_fd_sc_hd__nand2_1 _15602_ (.A(_08284_),
    .B(_08285_),
    .Y(_08286_));
 sky130_fd_sc_hd__a21oi_2 _15603_ (.A1(_08115_),
    .A2(_08161_),
    .B1(_08159_),
    .Y(_08287_));
 sky130_fd_sc_hd__xor2_1 _15604_ (.A(_08286_),
    .B(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__xnor2_1 _15605_ (.A(_08221_),
    .B(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__nor2_1 _15606_ (.A(_08162_),
    .B(_08164_),
    .Y(_08290_));
 sky130_fd_sc_hd__a21oi_1 _15607_ (.A1(_08093_),
    .A2(_08165_),
    .B1(_08290_),
    .Y(_08291_));
 sky130_fd_sc_hd__xnor2_1 _15608_ (.A(_08289_),
    .B(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__xnor2_1 _15609_ (.A(_08187_),
    .B(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__nand2_2 _15610_ (.A(_08185_),
    .B(_08293_),
    .Y(_08294_));
 sky130_fd_sc_hd__or2_1 _15611_ (.A(_08185_),
    .B(_08293_),
    .X(_08295_));
 sky130_fd_sc_hd__and2_1 _15612_ (.A(_08294_),
    .B(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__nand2_1 _15613_ (.A(_08183_),
    .B(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__or2_1 _15614_ (.A(_08183_),
    .B(_08296_),
    .X(_08298_));
 sky130_fd_sc_hd__and2_2 _15615_ (.A(_08297_),
    .B(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__nand2_1 _15616_ (.A(_08048_),
    .B(_08173_),
    .Y(_08300_));
 sky130_fd_sc_hd__nand2_1 _15617_ (.A(_08064_),
    .B(_08062_),
    .Y(_08301_));
 sky130_fd_sc_hd__a2bb2o_2 _15618_ (.A1_N(_08051_),
    .A2_N(_08300_),
    .B1(_08301_),
    .B2(_08172_),
    .X(_08302_));
 sky130_fd_sc_hd__xor2_4 _15619_ (.A(_08299_),
    .B(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__mux2_1 _15620_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_06851_),
    .X(_08304_));
 sky130_fd_sc_hd__nor2_1 _15621_ (.A(_08303_),
    .B(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _15622_ (.A(_08303_),
    .B(_08304_),
    .Y(_08306_));
 sky130_fd_sc_hd__and2b_1 _15623_ (.A_N(_08305_),
    .B(_08306_),
    .X(_08307_));
 sky130_fd_sc_hd__xnor2_1 _15624_ (.A(_07937_),
    .B(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__nor2_1 _15625_ (.A(_08182_),
    .B(_08308_),
    .Y(_08309_));
 sky130_fd_sc_hd__a21o_1 _15626_ (.A1(_08182_),
    .A2(_08308_),
    .B1(_04832_),
    .X(_08310_));
 sky130_fd_sc_hd__o221a_1 _15627_ (.A1(\rbzero.wall_tracer.texu[4] ),
    .A2(_06853_),
    .B1(_08309_),
    .B2(_08310_),
    .C1(_03498_),
    .X(_00479_));
 sky130_fd_sc_hd__a21o_1 _15628_ (.A1(_08182_),
    .A2(_08306_),
    .B1(_08305_),
    .X(_08311_));
 sky130_fd_sc_hd__a21bo_1 _15629_ (.A1(_08299_),
    .A2(_08302_),
    .B1_N(_08297_),
    .X(_08312_));
 sky130_fd_sc_hd__or2b_1 _15630_ (.A(_08220_),
    .B_N(_08188_),
    .X(_08313_));
 sky130_fd_sc_hd__a21boi_1 _15631_ (.A1(_08190_),
    .A2(_08219_),
    .B1_N(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__nand2_2 _15632_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_07256_),
    .Y(_08315_));
 sky130_fd_sc_hd__and2_1 _15633_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_07256_),
    .X(_08316_));
 sky130_fd_sc_hd__clkbuf_4 _15634_ (.A(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__xor2_1 _15635_ (.A(_08199_),
    .B(_08314_),
    .X(_08318_));
 sky130_fd_sc_hd__a21o_1 _15636_ (.A1(_07011_),
    .A2(_08317_),
    .B1(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__o31a_1 _15637_ (.A1(_07672_),
    .A2(_08314_),
    .A3(_08315_),
    .B1(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__or2_1 _15638_ (.A(_08286_),
    .B(_08287_),
    .X(_08321_));
 sky130_fd_sc_hd__nand2_1 _15639_ (.A(_08221_),
    .B(_08288_),
    .Y(_08322_));
 sky130_fd_sc_hd__a21o_1 _15640_ (.A1(_08201_),
    .A2(_08218_),
    .B1(_08216_),
    .X(_08323_));
 sky130_fd_sc_hd__or2b_1 _15641_ (.A(_08242_),
    .B_N(_08222_),
    .X(_08324_));
 sky130_fd_sc_hd__nor2_1 _15642_ (.A(_07972_),
    .B(_07959_),
    .Y(_08325_));
 sky130_fd_sc_hd__o22a_1 _15643_ (.A1(_07972_),
    .A2(_08081_),
    .B1(_07959_),
    .B2(_07856_),
    .X(_08326_));
 sky130_fd_sc_hd__a21oi_1 _15644_ (.A1(_08209_),
    .A2(_08325_),
    .B1(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__xnor2_1 _15645_ (.A(_08193_),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__o21a_1 _15646_ (.A1(_08192_),
    .A2(_08196_),
    .B1(_08194_),
    .X(_08329_));
 sky130_fd_sc_hd__or2_1 _15647_ (.A(_08328_),
    .B(_08329_),
    .X(_08330_));
 sky130_fd_sc_hd__nand2_1 _15648_ (.A(_08328_),
    .B(_08329_),
    .Y(_08331_));
 sky130_fd_sc_hd__nand2_1 _15649_ (.A(_08330_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__clkbuf_4 _15650_ (.A(_08191_),
    .X(_08333_));
 sky130_fd_sc_hd__nor2_1 _15651_ (.A(_07269_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__xnor2_1 _15652_ (.A(_08332_),
    .B(_08334_),
    .Y(_08335_));
 sky130_fd_sc_hd__o31ai_1 _15653_ (.A1(_07856_),
    .A2(_08081_),
    .A3(_08208_),
    .B1(_08207_),
    .Y(_08336_));
 sky130_fd_sc_hd__nand2_1 _15654_ (.A(_08097_),
    .B(_08224_),
    .Y(_08337_));
 sky130_fd_sc_hd__or3_1 _15655_ (.A(_07984_),
    .B(_07270_),
    .C(_08226_),
    .X(_08338_));
 sky130_fd_sc_hd__or2_1 _15656_ (.A(_07097_),
    .B(_07332_),
    .X(_08339_));
 sky130_fd_sc_hd__o22ai_1 _15657_ (.A1(_08107_),
    .A2(_07257_),
    .B1(_07333_),
    .B2(_07084_),
    .Y(_08340_));
 sky130_fd_sc_hd__o31a_1 _15658_ (.A1(_07084_),
    .A2(_07270_),
    .A3(_08339_),
    .B1(_08340_),
    .X(_08341_));
 sky130_fd_sc_hd__xnor2_1 _15659_ (.A(_08206_),
    .B(_08341_),
    .Y(_08342_));
 sky130_fd_sc_hd__a21oi_1 _15660_ (.A1(_08337_),
    .A2(_08338_),
    .B1(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__and3_1 _15661_ (.A(_08337_),
    .B(_08338_),
    .C(_08342_),
    .X(_08344_));
 sky130_fd_sc_hd__nor2_1 _15662_ (.A(_08343_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__xnor2_1 _15663_ (.A(_08336_),
    .B(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__a21oi_1 _15664_ (.A1(_08202_),
    .A2(_08213_),
    .B1(_08211_),
    .Y(_08347_));
 sky130_fd_sc_hd__nor2_1 _15665_ (.A(_08346_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__and2_1 _15666_ (.A(_08346_),
    .B(_08347_),
    .X(_08349_));
 sky130_fd_sc_hd__nor2_1 _15667_ (.A(_08348_),
    .B(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__xnor2_1 _15668_ (.A(_08335_),
    .B(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__a21o_1 _15669_ (.A1(_08240_),
    .A2(_08324_),
    .B1(_08351_),
    .X(_08352_));
 sky130_fd_sc_hd__nand3_1 _15670_ (.A(_08240_),
    .B(_08324_),
    .C(_08351_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand2_1 _15671_ (.A(_08352_),
    .B(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__xnor2_1 _15672_ (.A(_08323_),
    .B(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__or2_1 _15673_ (.A(_08281_),
    .B(_08282_),
    .X(_08356_));
 sky130_fd_sc_hd__a21o_1 _15674_ (.A1(_08228_),
    .A2(_08238_),
    .B1(_08236_),
    .X(_08357_));
 sky130_fd_sc_hd__a21bo_1 _15675_ (.A1(_08244_),
    .A2(_08254_),
    .B1_N(_08256_),
    .X(_08358_));
 sky130_fd_sc_hd__or2_1 _15676_ (.A(_06857_),
    .B(_08000_),
    .X(_08359_));
 sky130_fd_sc_hd__o22a_1 _15677_ (.A1(_07281_),
    .A2(_08000_),
    .B1(_07123_),
    .B2(_06858_),
    .X(_08360_));
 sky130_fd_sc_hd__o21ba_1 _15678_ (.A1(_08233_),
    .A2(_08359_),
    .B1_N(_08360_),
    .X(_08361_));
 sky130_fd_sc_hd__nand2_1 _15679_ (.A(_08224_),
    .B(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__or2_1 _15680_ (.A(_08224_),
    .B(_08361_),
    .X(_08363_));
 sky130_fd_sc_hd__and2_1 _15681_ (.A(_08362_),
    .B(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__nor2_1 _15682_ (.A(_08229_),
    .B(_07878_),
    .Y(_08365_));
 sky130_fd_sc_hd__or2_1 _15683_ (.A(_07494_),
    .B(_07198_),
    .X(_08366_));
 sky130_fd_sc_hd__or3_1 _15684_ (.A(_06997_),
    .B(_08252_),
    .C(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__o22ai_1 _15685_ (.A1(_07494_),
    .A2(_08252_),
    .B1(_07766_),
    .B2(_06997_),
    .Y(_08368_));
 sky130_fd_sc_hd__nand2_1 _15686_ (.A(_08367_),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__xor2_1 _15687_ (.A(_08365_),
    .B(_08369_),
    .X(_08370_));
 sky130_fd_sc_hd__o21a_1 _15688_ (.A1(_08232_),
    .A2(_08233_),
    .B1(_08230_),
    .X(_08371_));
 sky130_fd_sc_hd__xor2_1 _15689_ (.A(_08370_),
    .B(_08371_),
    .X(_08372_));
 sky130_fd_sc_hd__nand2_1 _15690_ (.A(_08364_),
    .B(_08372_),
    .Y(_08373_));
 sky130_fd_sc_hd__or2_1 _15691_ (.A(_08364_),
    .B(_08372_),
    .X(_08374_));
 sky130_fd_sc_hd__nand2_1 _15692_ (.A(_08373_),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__xor2_1 _15693_ (.A(_08358_),
    .B(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__xnor2_2 _15694_ (.A(_08357_),
    .B(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__or3_1 _15695_ (.A(_07992_),
    .B(_08252_),
    .C(_08251_),
    .X(_08378_));
 sky130_fd_sc_hd__a21bo_1 _15696_ (.A1(_08261_),
    .A2(_08263_),
    .B1_N(_08259_),
    .X(_08379_));
 sky130_fd_sc_hd__or2_1 _15697_ (.A(_07581_),
    .B(_07757_),
    .X(_08380_));
 sky130_fd_sc_hd__nor3_1 _15698_ (.A(_07100_),
    .B(_08133_),
    .C(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__o22a_1 _15699_ (.A1(_07581_),
    .A2(_07756_),
    .B1(_07757_),
    .B2(_07100_),
    .X(_08382_));
 sky130_fd_sc_hd__nor2_1 _15700_ (.A(_08381_),
    .B(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__xnor2_1 _15701_ (.A(_08249_),
    .B(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__xnor2_1 _15702_ (.A(_08379_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__a21o_1 _15703_ (.A1(_08250_),
    .A2(_08378_),
    .B1(_08385_),
    .X(_08386_));
 sky130_fd_sc_hd__nand3_1 _15704_ (.A(_08250_),
    .B(_08378_),
    .C(_08385_),
    .Y(_08387_));
 sky130_fd_sc_hd__and2_1 _15705_ (.A(_08386_),
    .B(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__nor2_1 _15706_ (.A(_07661_),
    .B(_08260_),
    .Y(_08389_));
 sky130_fd_sc_hd__a21oi_1 _15707_ (.A1(_03493_),
    .A2(\rbzero.wall_tracer.stepDistY[8] ),
    .B1(_04950_),
    .Y(_08390_));
 sky130_fd_sc_hd__a2bb2o_4 _15708_ (.A1_N(_04841_),
    .A2_N(\rbzero.wall_tracer.stepDistX[8] ),
    .B1(_08141_),
    .B2(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__or2_1 _15709_ (.A(_07646_),
    .B(_08391_),
    .X(_08392_));
 sky130_fd_sc_hd__o22ai_1 _15710_ (.A1(_07662_),
    .A2(_08018_),
    .B1(_08391_),
    .B2(_07213_),
    .Y(_08393_));
 sky130_fd_sc_hd__o21ai_1 _15711_ (.A1(_08265_),
    .A2(_08392_),
    .B1(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__xnor2_2 _15712_ (.A(_08389_),
    .B(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__nor2_1 _15713_ (.A(_04841_),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_08396_));
 sky130_fd_sc_hd__inv_2 _15714_ (.A(\rbzero.wall_tracer.stepDistY[10] ),
    .Y(_08397_));
 sky130_fd_sc_hd__o21a_1 _15715_ (.A1(_06781_),
    .A2(_08267_),
    .B1(_04832_),
    .X(_08398_));
 sky130_fd_sc_hd__o221a_1 _15716_ (.A1(_06860_),
    .A2(_08397_),
    .B1(_07162_),
    .B2(_08398_),
    .C1(_04841_),
    .X(_08399_));
 sky130_fd_sc_hd__or4_1 _15717_ (.A(_03388_),
    .B(_07185_),
    .C(_08396_),
    .D(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__o41ai_1 _15718_ (.A1(_07175_),
    .A2(_04950_),
    .A3(_03493_),
    .A4(_08399_),
    .B1(_08315_),
    .Y(_08401_));
 sky130_fd_sc_hd__nand2_1 _15719_ (.A(_08400_),
    .B(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__xnor2_2 _15720_ (.A(_08270_),
    .B(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__and3_1 _15721_ (.A(_07673_),
    .B(_08144_),
    .C(_08272_),
    .X(_08404_));
 sky130_fd_sc_hd__a21o_1 _15722_ (.A1(_08145_),
    .A2(_08270_),
    .B1(_08404_),
    .X(_08405_));
 sky130_fd_sc_hd__xor2_2 _15723_ (.A(_08403_),
    .B(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__xnor2_2 _15724_ (.A(_08395_),
    .B(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__and2_1 _15725_ (.A(_08273_),
    .B(_08274_),
    .X(_08408_));
 sky130_fd_sc_hd__a21oi_2 _15726_ (.A1(_08264_),
    .A2(_08275_),
    .B1(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__xor2_2 _15727_ (.A(_08407_),
    .B(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__xnor2_1 _15728_ (.A(_08388_),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__a21oi_1 _15729_ (.A1(_08258_),
    .A2(_08280_),
    .B1(_08278_),
    .Y(_08412_));
 sky130_fd_sc_hd__nor2_1 _15730_ (.A(_08411_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__nand2_1 _15731_ (.A(_08411_),
    .B(_08412_),
    .Y(_08414_));
 sky130_fd_sc_hd__and2b_1 _15732_ (.A_N(_08413_),
    .B(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__xnor2_2 _15733_ (.A(_08377_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__a21oi_1 _15734_ (.A1(_08356_),
    .A2(_08284_),
    .B1(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__and3_1 _15735_ (.A(_08356_),
    .B(_08284_),
    .C(_08416_),
    .X(_08418_));
 sky130_fd_sc_hd__nor2_1 _15736_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__xnor2_1 _15737_ (.A(_08355_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__a21oi_1 _15738_ (.A1(_08321_),
    .A2(_08322_),
    .B1(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__and3_1 _15739_ (.A(_08321_),
    .B(_08322_),
    .C(_08420_),
    .X(_08422_));
 sky130_fd_sc_hd__nor2_1 _15740_ (.A(_08421_),
    .B(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__xnor2_1 _15741_ (.A(_08320_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__or2b_1 _15742_ (.A(_08292_),
    .B_N(_08187_),
    .X(_08425_));
 sky130_fd_sc_hd__o21a_1 _15743_ (.A1(_08289_),
    .A2(_08291_),
    .B1(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__nor2_1 _15744_ (.A(_08424_),
    .B(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__and2_1 _15745_ (.A(_08424_),
    .B(_08426_),
    .X(_08428_));
 sky130_fd_sc_hd__nor2_2 _15746_ (.A(_08427_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__xnor2_4 _15747_ (.A(_08294_),
    .B(_08429_),
    .Y(_08430_));
 sky130_fd_sc_hd__xor2_4 _15748_ (.A(_08312_),
    .B(_08430_),
    .X(_08431_));
 sky130_fd_sc_hd__mux2_1 _15749_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_06851_),
    .X(_08432_));
 sky130_fd_sc_hd__xnor2_1 _15750_ (.A(_07827_),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__xnor2_1 _15751_ (.A(_08431_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__nor2_1 _15752_ (.A(_08311_),
    .B(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__a21o_1 _15753_ (.A1(_08311_),
    .A2(_08434_),
    .B1(_04832_),
    .X(_08436_));
 sky130_fd_sc_hd__o221a_1 _15754_ (.A1(\rbzero.wall_tracer.texu[5] ),
    .A2(_06853_),
    .B1(_08435_),
    .B2(_08436_),
    .C1(_03485_),
    .X(_00480_));
 sky130_fd_sc_hd__or2_1 _15755_ (.A(_03337_),
    .B(_03506_),
    .X(_08437_));
 sky130_fd_sc_hd__clkbuf_2 _15756_ (.A(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__nor2_1 _15757_ (.A(_02899_),
    .B(_08438_),
    .Y(_00481_));
 sky130_fd_sc_hd__nor2_8 _15758_ (.A(_02981_),
    .B(_03506_),
    .Y(_08439_));
 sky130_fd_sc_hd__and3b_1 _15759_ (.A_N(_03501_),
    .B(_03809_),
    .C(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__clkbuf_1 _15760_ (.A(_08440_),
    .X(_00482_));
 sky130_fd_sc_hd__or2_1 _15761_ (.A(_03526_),
    .B(_03501_),
    .X(_08441_));
 sky130_fd_sc_hd__and3_1 _15762_ (.A(_03502_),
    .B(_08441_),
    .C(_08439_),
    .X(_08442_));
 sky130_fd_sc_hd__clkbuf_1 _15763_ (.A(_08442_),
    .X(_00483_));
 sky130_fd_sc_hd__nor2_1 _15764_ (.A(_04040_),
    .B(_08438_),
    .Y(_00484_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(net61),
    .B(_04054_),
    .Y(_00485_));
 sky130_fd_sc_hd__nor2_1 _15766_ (.A(_04062_),
    .B(_08438_),
    .Y(_00486_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_04035_),
    .B(_08438_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_1 _15768_ (.A(_04076_),
    .B(_08438_),
    .Y(_00488_));
 sky130_fd_sc_hd__and4_1 _15769_ (.A(_02901_),
    .B(_03838_),
    .C(_03459_),
    .D(_04034_),
    .X(_08443_));
 sky130_fd_sc_hd__a31o_1 _15770_ (.A1(_02901_),
    .A2(_03838_),
    .A3(_04034_),
    .B1(_03459_),
    .X(_08444_));
 sky130_fd_sc_hd__and3b_1 _15771_ (.A_N(_08443_),
    .B(_08439_),
    .C(_08444_),
    .X(_08445_));
 sky130_fd_sc_hd__clkbuf_1 _15772_ (.A(_08445_),
    .X(_00489_));
 sky130_fd_sc_hd__a21oi_1 _15773_ (.A1(_03469_),
    .A2(_08443_),
    .B1(_08438_),
    .Y(_08446_));
 sky130_fd_sc_hd__o21a_1 _15774_ (.A1(_03469_),
    .A2(_08443_),
    .B1(_08446_),
    .X(_00490_));
 sky130_fd_sc_hd__buf_4 _15775_ (.A(_03508_),
    .X(_08447_));
 sky130_fd_sc_hd__buf_4 _15776_ (.A(_08447_),
    .X(_08448_));
 sky130_fd_sc_hd__buf_4 _15777_ (.A(_08448_),
    .X(_08449_));
 sky130_fd_sc_hd__and4_2 _15778_ (.A(_03474_),
    .B(_04019_),
    .C(_04053_),
    .D(_03911_),
    .X(_08450_));
 sky130_fd_sc_hd__and3_1 _15779_ (.A(\rbzero.wall_tracer.state[14] ),
    .B(_03484_),
    .C(_08450_),
    .X(_08451_));
 sky130_fd_sc_hd__clkbuf_4 _15780_ (.A(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__buf_4 _15781_ (.A(_08452_),
    .X(_08453_));
 sky130_fd_sc_hd__a22o_1 _15782_ (.A1(\rbzero.row_render.side ),
    .A2(_08449_),
    .B1(_08453_),
    .B2(_06851_),
    .X(_00491_));
 sky130_fd_sc_hd__buf_4 _15783_ (.A(_08452_),
    .X(_08454_));
 sky130_fd_sc_hd__a22o_1 _15784_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_08449_),
    .B1(_06669_),
    .B2(_08454_),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _15785_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_08449_),
    .B1(_06679_),
    .B2(_08454_),
    .X(_00493_));
 sky130_fd_sc_hd__a22o_1 _15786_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_08449_),
    .B1(_06686_),
    .B2(_08454_),
    .X(_00494_));
 sky130_fd_sc_hd__buf_2 _15787_ (.A(_08452_),
    .X(_08455_));
 sky130_fd_sc_hd__a22o_1 _15788_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_08449_),
    .B1(_06695_),
    .B2(_08455_),
    .X(_00495_));
 sky130_fd_sc_hd__clkbuf_4 _15789_ (.A(_08448_),
    .X(_08456_));
 sky130_fd_sc_hd__a22o_1 _15790_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_08456_),
    .B1(_06705_),
    .B2(_08455_),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_1 _15791_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_08456_),
    .B1(_06712_),
    .B2(_08455_),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _15792_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_08456_),
    .B1(_06717_),
    .B2(_08455_),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_1 _15793_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_08456_),
    .B1(_06726_),
    .B2(_08455_),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _15794_ (.A1(\rbzero.row_render.size[8] ),
    .A2(_08456_),
    .B1(_06733_),
    .B2(_08455_),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _15795_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_08456_),
    .B1(_06738_),
    .B2(_08455_),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_1 _15796_ (.A1(\rbzero.row_render.size[10] ),
    .A2(_08456_),
    .B1(_06746_),
    .B2(_08455_),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _15797_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_08456_),
    .B1(_08453_),
    .B2(\rbzero.wall_tracer.texu[0] ),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _15798_ (.A1(\rbzero.row_render.texu[1] ),
    .A2(_08456_),
    .B1(_08453_),
    .B2(\rbzero.wall_tracer.texu[1] ),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _15799_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_08456_),
    .B1(_08453_),
    .B2(\rbzero.wall_tracer.texu[2] ),
    .X(_00505_));
 sky130_fd_sc_hd__clkbuf_4 _15800_ (.A(_08448_),
    .X(_08457_));
 sky130_fd_sc_hd__a22o_1 _15801_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(_08457_),
    .B1(_08453_),
    .B2(\rbzero.wall_tracer.texu[3] ),
    .X(_00506_));
 sky130_fd_sc_hd__a22o_1 _15802_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_08457_),
    .B1(_08453_),
    .B2(\rbzero.wall_tracer.texu[4] ),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _15803_ (.A1(\rbzero.row_render.texu[5] ),
    .A2(_08457_),
    .B1(_08453_),
    .B2(\rbzero.wall_tracer.texu[5] ),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _15804_ (.A1(\rbzero.traced_texa[-11] ),
    .A2(_08457_),
    .B1(_08453_),
    .B2(_06787_),
    .X(_00509_));
 sky130_fd_sc_hd__a22o_1 _15805_ (.A1(\rbzero.traced_texa[-10] ),
    .A2(_08457_),
    .B1(_08453_),
    .B2(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_00510_));
 sky130_fd_sc_hd__buf_4 _15806_ (.A(_08452_),
    .X(_08458_));
 sky130_fd_sc_hd__buf_2 _15807_ (.A(_08458_),
    .X(_08459_));
 sky130_fd_sc_hd__a22o_1 _15808_ (.A1(\rbzero.traced_texa[-9] ),
    .A2(_08457_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00511_));
 sky130_fd_sc_hd__a22o_1 _15809_ (.A1(\rbzero.traced_texa[-8] ),
    .A2(_08457_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _15810_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(_08457_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(_00513_));
 sky130_fd_sc_hd__a22o_1 _15811_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(_08457_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_1 _15812_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(_08457_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(_00515_));
 sky130_fd_sc_hd__clkbuf_4 _15813_ (.A(_08447_),
    .X(_08460_));
 sky130_fd_sc_hd__clkbuf_4 _15814_ (.A(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__a22o_1 _15815_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(_08461_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(_00516_));
 sky130_fd_sc_hd__a22o_1 _15816_ (.A1(\rbzero.traced_texa[-3] ),
    .A2(_08461_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _15817_ (.A1(\rbzero.traced_texa[-2] ),
    .A2(_08461_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_00518_));
 sky130_fd_sc_hd__a22o_1 _15818_ (.A1(\rbzero.traced_texa[-1] ),
    .A2(_08461_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_00519_));
 sky130_fd_sc_hd__a22o_1 _15819_ (.A1(\rbzero.traced_texa[0] ),
    .A2(_08461_),
    .B1(_08459_),
    .B2(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_00520_));
 sky130_fd_sc_hd__clkbuf_4 _15820_ (.A(_08458_),
    .X(_08462_));
 sky130_fd_sc_hd__a22o_1 _15821_ (.A1(\rbzero.traced_texa[1] ),
    .A2(_08461_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_00521_));
 sky130_fd_sc_hd__a22o_1 _15822_ (.A1(\rbzero.traced_texa[2] ),
    .A2(_08461_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_00522_));
 sky130_fd_sc_hd__a22o_1 _15823_ (.A1(\rbzero.traced_texa[3] ),
    .A2(_08461_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(_00523_));
 sky130_fd_sc_hd__a22o_1 _15824_ (.A1(\rbzero.traced_texa[4] ),
    .A2(_08461_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_00524_));
 sky130_fd_sc_hd__a22o_1 _15825_ (.A1(\rbzero.traced_texa[5] ),
    .A2(_08461_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_00525_));
 sky130_fd_sc_hd__buf_4 _15826_ (.A(_08460_),
    .X(_08463_));
 sky130_fd_sc_hd__a22o_1 _15827_ (.A1(\rbzero.traced_texa[6] ),
    .A2(_08463_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_00526_));
 sky130_fd_sc_hd__a22o_1 _15828_ (.A1(\rbzero.traced_texa[7] ),
    .A2(_08463_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_00527_));
 sky130_fd_sc_hd__a22o_1 _15829_ (.A1(\rbzero.traced_texa[8] ),
    .A2(_08463_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_00528_));
 sky130_fd_sc_hd__a22o_1 _15830_ (.A1(\rbzero.traced_texa[9] ),
    .A2(_08463_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_00529_));
 sky130_fd_sc_hd__a22o_1 _15831_ (.A1(\rbzero.traced_texa[10] ),
    .A2(_08463_),
    .B1(_08462_),
    .B2(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_00530_));
 sky130_fd_sc_hd__nand3_4 _15832_ (.A(\rbzero.wall_tracer.state[14] ),
    .B(_03484_),
    .C(_08450_),
    .Y(_08464_));
 sky130_fd_sc_hd__mux2_1 _15833_ (.A0(\rbzero.wall_tracer.wall[0] ),
    .A1(\rbzero.row_render.wall[0] ),
    .S(_08464_),
    .X(_08465_));
 sky130_fd_sc_hd__clkbuf_1 _15834_ (.A(_08465_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _15835_ (.A0(\rbzero.wall_tracer.wall[1] ),
    .A1(\rbzero.row_render.wall[1] ),
    .S(_08464_),
    .X(_08466_));
 sky130_fd_sc_hd__clkbuf_1 _15836_ (.A(_08466_),
    .X(_00532_));
 sky130_fd_sc_hd__o21a_1 _15837_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(\rbzero.wall_tracer.mapX[5] ),
    .B1(_07825_),
    .X(_08467_));
 sky130_fd_sc_hd__xor2_1 _15838_ (.A(\rbzero.wall_tracer.mapX[5] ),
    .B(_07825_),
    .X(_08468_));
 sky130_fd_sc_hd__nor2_1 _15839_ (.A(_03364_),
    .B(_07936_),
    .Y(_08469_));
 sky130_fd_sc_hd__nor2_1 _15840_ (.A(\rbzero.map_rom.i_col[4] ),
    .B(_07825_),
    .Y(_08470_));
 sky130_fd_sc_hd__nor2_1 _15841_ (.A(_08469_),
    .B(_08470_),
    .Y(_08471_));
 sky130_fd_sc_hd__xnor2_1 _15842_ (.A(_03362_),
    .B(_06914_),
    .Y(_08472_));
 sky130_fd_sc_hd__nand2_1 _15843_ (.A(_03395_),
    .B(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__o21ai_1 _15844_ (.A1(_03362_),
    .A2(_07936_),
    .B1(_08473_),
    .Y(_08474_));
 sky130_fd_sc_hd__nand2_1 _15845_ (.A(_03353_),
    .B(_07825_),
    .Y(_08475_));
 sky130_fd_sc_hd__or2_1 _15846_ (.A(_03353_),
    .B(_06914_),
    .X(_08476_));
 sky130_fd_sc_hd__and2_1 _15847_ (.A(_08475_),
    .B(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__a21bo_1 _15848_ (.A1(_08474_),
    .A2(_08477_),
    .B1_N(_08475_),
    .X(_08478_));
 sky130_fd_sc_hd__a21o_1 _15849_ (.A1(_03369_),
    .A2(_07825_),
    .B1(_08478_),
    .X(_08479_));
 sky130_fd_sc_hd__o21a_1 _15850_ (.A1(_03369_),
    .A2(_07825_),
    .B1(_08479_),
    .X(_08480_));
 sky130_fd_sc_hd__and3_1 _15851_ (.A(_08468_),
    .B(_08471_),
    .C(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__xor2_1 _15852_ (.A(\rbzero.wall_tracer.mapX[6] ),
    .B(_07825_),
    .X(_08482_));
 sky130_fd_sc_hd__o21ai_1 _15853_ (.A1(_08467_),
    .A2(_08481_),
    .B1(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__or3_1 _15854_ (.A(_08482_),
    .B(_08467_),
    .C(_08481_),
    .X(_08484_));
 sky130_fd_sc_hd__buf_4 _15855_ (.A(_03341_),
    .X(_08485_));
 sky130_fd_sc_hd__or3b_1 _15856_ (.A(_04951_),
    .B(_04952_),
    .C_N(_06784_),
    .X(_08486_));
 sky130_fd_sc_hd__buf_2 _15857_ (.A(_08486_),
    .X(_08487_));
 sky130_fd_sc_hd__nor2_2 _15858_ (.A(_08485_),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__buf_4 _15859_ (.A(_08487_),
    .X(_08489_));
 sky130_fd_sc_hd__a32o_1 _15860_ (.A1(_08483_),
    .A2(_08484_),
    .A3(_08488_),
    .B1(_08489_),
    .B2(\rbzero.wall_tracer.mapX[6] ),
    .X(_00533_));
 sky130_fd_sc_hd__xor2_1 _15861_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(_07825_),
    .X(_08490_));
 sky130_fd_sc_hd__a21boi_1 _15862_ (.A1(\rbzero.wall_tracer.mapX[6] ),
    .A2(_07826_),
    .B1_N(_08483_),
    .Y(_08491_));
 sky130_fd_sc_hd__xnor2_1 _15863_ (.A(_08490_),
    .B(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__a22o_1 _15864_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(_08489_),
    .B1(_08488_),
    .B2(_08492_),
    .X(_00534_));
 sky130_fd_sc_hd__xor2_1 _15865_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(_07826_),
    .X(_08493_));
 sky130_fd_sc_hd__and3_1 _15866_ (.A(_08482_),
    .B(_08481_),
    .C(_08490_),
    .X(_08494_));
 sky130_fd_sc_hd__o21a_1 _15867_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(\rbzero.wall_tracer.mapX[6] ),
    .B1(_07825_),
    .X(_08495_));
 sky130_fd_sc_hd__or3_1 _15868_ (.A(_08467_),
    .B(_08494_),
    .C(_08495_),
    .X(_08496_));
 sky130_fd_sc_hd__xor2_1 _15869_ (.A(_08493_),
    .B(_08496_),
    .X(_08497_));
 sky130_fd_sc_hd__a22o_1 _15870_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_08489_),
    .B1(_08488_),
    .B2(_08497_),
    .X(_00535_));
 sky130_fd_sc_hd__a22o_1 _15871_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_07826_),
    .B1(_08493_),
    .B2(_08496_),
    .X(_08498_));
 sky130_fd_sc_hd__xnor2_1 _15872_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(_07826_),
    .Y(_08499_));
 sky130_fd_sc_hd__xnor2_1 _15873_ (.A(_08498_),
    .B(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__a22o_1 _15874_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_08489_),
    .B1(_08488_),
    .B2(_08500_),
    .X(_00536_));
 sky130_fd_sc_hd__o21a_1 _15875_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_07826_),
    .B1(_08498_),
    .X(_08501_));
 sky130_fd_sc_hd__a21oi_1 _15876_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_07826_),
    .B1(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__xnor2_1 _15877_ (.A(\rbzero.wall_tracer.mapX[10] ),
    .B(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__nand2_1 _15878_ (.A(_07826_),
    .B(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__or2_1 _15879_ (.A(_07826_),
    .B(_08503_),
    .X(_08505_));
 sky130_fd_sc_hd__a32o_1 _15880_ (.A1(_08488_),
    .A2(_08504_),
    .A3(_08505_),
    .B1(_08489_),
    .B2(\rbzero.wall_tracer.mapX[10] ),
    .X(_00537_));
 sky130_fd_sc_hd__and4b_4 _15881_ (.A_N(_04951_),
    .B(_03484_),
    .C(_03458_),
    .D(_06784_),
    .X(_08506_));
 sky130_fd_sc_hd__buf_4 _15882_ (.A(_08506_),
    .X(_08507_));
 sky130_fd_sc_hd__clkbuf_4 _15883_ (.A(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__buf_8 _15884_ (.A(\rbzero.wall_tracer.state[1] ),
    .X(_08509_));
 sky130_fd_sc_hd__a21oi_1 _15885_ (.A1(_07642_),
    .A2(_07691_),
    .B1(_08509_),
    .Y(_08510_));
 sky130_fd_sc_hd__o21a_1 _15886_ (.A1(_07642_),
    .A2(_07691_),
    .B1(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__buf_4 _15887_ (.A(_08509_),
    .X(_08512_));
 sky130_fd_sc_hd__nand2_1 _15888_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .Y(_08513_));
 sky130_fd_sc_hd__or2_1 _15889_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .X(_08514_));
 sky130_fd_sc_hd__a31o_1 _15890_ (.A1(_08512_),
    .A2(_08513_),
    .A3(_08514_),
    .B1(_08489_),
    .X(_08515_));
 sky130_fd_sc_hd__o22a_1 _15891_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(_08508_),
    .B1(_08511_),
    .B2(_08515_),
    .X(_00538_));
 sky130_fd_sc_hd__a21oi_1 _15892_ (.A1(_07693_),
    .A2(_07695_),
    .B1(_08509_),
    .Y(_08516_));
 sky130_fd_sc_hd__o21a_1 _15893_ (.A1(_07693_),
    .A2(_07695_),
    .B1(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__or2_1 _15894_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_08518_));
 sky130_fd_sc_hd__nand2_1 _15895_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_08519_));
 sky130_fd_sc_hd__nand3b_1 _15896_ (.A_N(_08513_),
    .B(_08518_),
    .C(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__a21bo_1 _15897_ (.A1(_08518_),
    .A2(_08519_),
    .B1_N(_08513_),
    .X(_08521_));
 sky130_fd_sc_hd__clkbuf_4 _15898_ (.A(_08487_),
    .X(_08522_));
 sky130_fd_sc_hd__a31o_1 _15899_ (.A1(_08512_),
    .A2(_08520_),
    .A3(_08521_),
    .B1(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__o22a_1 _15900_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(_08508_),
    .B1(_08517_),
    .B2(_08523_),
    .X(_00539_));
 sky130_fd_sc_hd__clkbuf_4 _15901_ (.A(_03341_),
    .X(_08524_));
 sky130_fd_sc_hd__and2_1 _15902_ (.A(_08524_),
    .B(_07817_),
    .X(_08525_));
 sky130_fd_sc_hd__and2_1 _15903_ (.A(_08519_),
    .B(_08520_),
    .X(_08526_));
 sky130_fd_sc_hd__nor2_1 _15904_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .Y(_08527_));
 sky130_fd_sc_hd__and2_1 _15905_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_08528_));
 sky130_fd_sc_hd__or3_1 _15906_ (.A(_08526_),
    .B(_08527_),
    .C(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__o21ai_1 _15907_ (.A1(_08527_),
    .A2(_08528_),
    .B1(_08526_),
    .Y(_08530_));
 sky130_fd_sc_hd__a31o_1 _15908_ (.A1(_08512_),
    .A2(_08529_),
    .A3(_08530_),
    .B1(_08522_),
    .X(_08531_));
 sky130_fd_sc_hd__o22a_1 _15909_ (.A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .A2(_08508_),
    .B1(_08525_),
    .B2(_08531_),
    .X(_00540_));
 sky130_fd_sc_hd__and2_1 _15910_ (.A(_08524_),
    .B(_07815_),
    .X(_08532_));
 sky130_fd_sc_hd__or2_1 _15911_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_08533_));
 sky130_fd_sc_hd__nand2_1 _15912_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_08534_));
 sky130_fd_sc_hd__o21bai_1 _15913_ (.A1(_08526_),
    .A2(_08527_),
    .B1_N(_08528_),
    .Y(_08535_));
 sky130_fd_sc_hd__nand3_1 _15914_ (.A(_08533_),
    .B(_08534_),
    .C(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__a21o_1 _15915_ (.A1(_08533_),
    .A2(_08534_),
    .B1(_08535_),
    .X(_08537_));
 sky130_fd_sc_hd__a31o_1 _15916_ (.A1(_08512_),
    .A2(_08536_),
    .A3(_08537_),
    .B1(_08522_),
    .X(_08538_));
 sky130_fd_sc_hd__o22a_1 _15917_ (.A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .A2(_08508_),
    .B1(_08532_),
    .B2(_08538_),
    .X(_00541_));
 sky130_fd_sc_hd__and2_1 _15918_ (.A(_08524_),
    .B(_07813_),
    .X(_08539_));
 sky130_fd_sc_hd__nor2_1 _15919_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_08540_));
 sky130_fd_sc_hd__and2_1 _15920_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .X(_08541_));
 sky130_fd_sc_hd__a21boi_1 _15921_ (.A1(_08533_),
    .A2(_08535_),
    .B1_N(_08534_),
    .Y(_08542_));
 sky130_fd_sc_hd__or3_1 _15922_ (.A(_08540_),
    .B(_08541_),
    .C(_08542_),
    .X(_08543_));
 sky130_fd_sc_hd__o21ai_1 _15923_ (.A1(_08540_),
    .A2(_08541_),
    .B1(_08542_),
    .Y(_08544_));
 sky130_fd_sc_hd__a31o_1 _15924_ (.A1(_08512_),
    .A2(_08543_),
    .A3(_08544_),
    .B1(_08522_),
    .X(_08545_));
 sky130_fd_sc_hd__o22a_1 _15925_ (.A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .A2(_08508_),
    .B1(_08539_),
    .B2(_08545_),
    .X(_00542_));
 sky130_fd_sc_hd__and2_1 _15926_ (.A(_08524_),
    .B(_07808_),
    .X(_08546_));
 sky130_fd_sc_hd__or2_1 _15927_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_08547_));
 sky130_fd_sc_hd__nand2_1 _15928_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_08548_));
 sky130_fd_sc_hd__o21bai_1 _15929_ (.A1(_08540_),
    .A2(_08542_),
    .B1_N(_08541_),
    .Y(_08549_));
 sky130_fd_sc_hd__a21oi_1 _15930_ (.A1(_08547_),
    .A2(_08548_),
    .B1(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__a31o_1 _15931_ (.A1(_08547_),
    .A2(_08548_),
    .A3(_08549_),
    .B1(_04946_),
    .X(_08551_));
 sky130_fd_sc_hd__o21ai_1 _15932_ (.A1(_08550_),
    .A2(_08551_),
    .B1(_08507_),
    .Y(_08552_));
 sky130_fd_sc_hd__o22a_1 _15933_ (.A1(\rbzero.wall_tracer.trackDistX[-6] ),
    .A2(_08508_),
    .B1(_08546_),
    .B2(_08552_),
    .X(_00543_));
 sky130_fd_sc_hd__clkbuf_4 _15934_ (.A(_08507_),
    .X(_08553_));
 sky130_fd_sc_hd__and2_1 _15935_ (.A(_08524_),
    .B(_07929_),
    .X(_08554_));
 sky130_fd_sc_hd__nor2_1 _15936_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_08555_));
 sky130_fd_sc_hd__and2_1 _15937_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .X(_08556_));
 sky130_fd_sc_hd__a21boi_1 _15938_ (.A1(_08547_),
    .A2(_08549_),
    .B1_N(_08548_),
    .Y(_08557_));
 sky130_fd_sc_hd__or3_1 _15939_ (.A(_08555_),
    .B(_08556_),
    .C(_08557_),
    .X(_08558_));
 sky130_fd_sc_hd__o21ai_1 _15940_ (.A1(_08555_),
    .A2(_08556_),
    .B1(_08557_),
    .Y(_08559_));
 sky130_fd_sc_hd__a31o_1 _15941_ (.A1(_08512_),
    .A2(_08558_),
    .A3(_08559_),
    .B1(_08522_),
    .X(_08560_));
 sky130_fd_sc_hd__o22a_1 _15942_ (.A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .A2(_08553_),
    .B1(_08554_),
    .B2(_08560_),
    .X(_00544_));
 sky130_fd_sc_hd__and2_1 _15943_ (.A(_08524_),
    .B(_08052_),
    .X(_08561_));
 sky130_fd_sc_hd__clkbuf_4 _15944_ (.A(_08509_),
    .X(_08562_));
 sky130_fd_sc_hd__or2_1 _15945_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(_08563_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_08564_));
 sky130_fd_sc_hd__o21bai_1 _15947_ (.A1(_08555_),
    .A2(_08557_),
    .B1_N(_08556_),
    .Y(_08565_));
 sky130_fd_sc_hd__nand3_1 _15948_ (.A(_08563_),
    .B(_08564_),
    .C(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__a21o_1 _15949_ (.A1(_08563_),
    .A2(_08564_),
    .B1(_08565_),
    .X(_08567_));
 sky130_fd_sc_hd__a31o_1 _15950_ (.A1(_08562_),
    .A2(_08566_),
    .A3(_08567_),
    .B1(_08522_),
    .X(_08568_));
 sky130_fd_sc_hd__o22a_1 _15951_ (.A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .A2(_08553_),
    .B1(_08561_),
    .B2(_08568_),
    .X(_00545_));
 sky130_fd_sc_hd__inv_2 _15952_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .Y(_08569_));
 sky130_fd_sc_hd__nor2_1 _15953_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_08570_));
 sky130_fd_sc_hd__nor2_1 _15954_ (.A(_08569_),
    .B(_06907_),
    .Y(_08571_));
 sky130_fd_sc_hd__a21boi_1 _15955_ (.A1(_08563_),
    .A2(_08565_),
    .B1_N(_08564_),
    .Y(_08572_));
 sky130_fd_sc_hd__nor3_1 _15956_ (.A(_08570_),
    .B(_08571_),
    .C(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__o21a_1 _15957_ (.A1(_08570_),
    .A2(_08571_),
    .B1(_08572_),
    .X(_08574_));
 sky130_fd_sc_hd__nand2_1 _15958_ (.A(_04946_),
    .B(_08174_),
    .Y(_08575_));
 sky130_fd_sc_hd__o311a_1 _15959_ (.A1(_08485_),
    .A2(_08573_),
    .A3(_08574_),
    .B1(_08507_),
    .C1(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__a21oi_1 _15960_ (.A1(_08569_),
    .A2(_08489_),
    .B1(_08576_),
    .Y(_00546_));
 sky130_fd_sc_hd__and2_1 _15961_ (.A(_08524_),
    .B(_08303_),
    .X(_08577_));
 sky130_fd_sc_hd__or2_1 _15962_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_08578_));
 sky130_fd_sc_hd__nand2_1 _15963_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_08579_));
 sky130_fd_sc_hd__o21bai_2 _15964_ (.A1(_08570_),
    .A2(_08572_),
    .B1_N(_08571_),
    .Y(_08580_));
 sky130_fd_sc_hd__nand3_1 _15965_ (.A(_08578_),
    .B(_08579_),
    .C(_08580_),
    .Y(_08581_));
 sky130_fd_sc_hd__a21o_1 _15966_ (.A1(_08578_),
    .A2(_08579_),
    .B1(_08580_),
    .X(_08582_));
 sky130_fd_sc_hd__a31o_1 _15967_ (.A1(_08562_),
    .A2(_08581_),
    .A3(_08582_),
    .B1(_08522_),
    .X(_08583_));
 sky130_fd_sc_hd__o22a_1 _15968_ (.A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .A2(_08553_),
    .B1(_08577_),
    .B2(_08583_),
    .X(_00547_));
 sky130_fd_sc_hd__nand2_1 _15969_ (.A(_04946_),
    .B(_08431_),
    .Y(_08584_));
 sky130_fd_sc_hd__inv_2 _15970_ (.A(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__and2_1 _15971_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(_08586_));
 sky130_fd_sc_hd__nor2_1 _15972_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_08587_));
 sky130_fd_sc_hd__a21boi_1 _15973_ (.A1(_08578_),
    .A2(_08580_),
    .B1_N(_08579_),
    .Y(_08588_));
 sky130_fd_sc_hd__or3_1 _15974_ (.A(_08586_),
    .B(_08587_),
    .C(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__o21ai_1 _15975_ (.A1(_08586_),
    .A2(_08587_),
    .B1(_08588_),
    .Y(_08590_));
 sky130_fd_sc_hd__a31o_1 _15976_ (.A1(_08562_),
    .A2(_08589_),
    .A3(_08590_),
    .B1(_08522_),
    .X(_08591_));
 sky130_fd_sc_hd__o22a_1 _15977_ (.A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .A2(_08553_),
    .B1(_08585_),
    .B2(_08591_),
    .X(_00548_));
 sky130_fd_sc_hd__nor2_1 _15978_ (.A(_04966_),
    .B(_07102_),
    .Y(_08592_));
 sky130_fd_sc_hd__nor2_1 _15979_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_08593_));
 sky130_fd_sc_hd__nand2_1 _15980_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_08594_));
 sky130_fd_sc_hd__o211a_1 _15981_ (.A1(_08592_),
    .A2(_08593_),
    .B1(_08594_),
    .C1(_08589_),
    .X(_08595_));
 sky130_fd_sc_hd__a211oi_2 _15982_ (.A1(_08594_),
    .A2(_08589_),
    .B1(_08592_),
    .C1(_08593_),
    .Y(_08596_));
 sky130_fd_sc_hd__nor2_1 _15983_ (.A(_08199_),
    .B(_08314_),
    .Y(_08597_));
 sky130_fd_sc_hd__a31o_1 _15984_ (.A1(_07011_),
    .A2(_08318_),
    .A3(_08317_),
    .B1(_08597_),
    .X(_08598_));
 sky130_fd_sc_hd__or2b_1 _15985_ (.A(_08354_),
    .B_N(_08323_),
    .X(_08599_));
 sky130_fd_sc_hd__o31a_1 _15986_ (.A1(_07269_),
    .A2(_08333_),
    .A3(_08332_),
    .B1(_08330_),
    .X(_08600_));
 sky130_fd_sc_hd__a21oi_1 _15987_ (.A1(_08352_),
    .A2(_08599_),
    .B1(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__and3_1 _15988_ (.A(_08352_),
    .B(_08599_),
    .C(_08600_),
    .X(_08602_));
 sky130_fd_sc_hd__nor2_1 _15989_ (.A(_08601_),
    .B(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__a21o_1 _15990_ (.A1(_08335_),
    .A2(_08350_),
    .B1(_08348_),
    .X(_08604_));
 sky130_fd_sc_hd__or2b_1 _15991_ (.A(_08375_),
    .B_N(_08358_),
    .X(_08605_));
 sky130_fd_sc_hd__or2b_1 _15992_ (.A(_08376_),
    .B_N(_08357_),
    .X(_08606_));
 sky130_fd_sc_hd__nor2_1 _15993_ (.A(_07265_),
    .B(_08191_),
    .Y(_08607_));
 sky130_fd_sc_hd__nor2_1 _15994_ (.A(_07856_),
    .B(_08070_),
    .Y(_08608_));
 sky130_fd_sc_hd__or4_1 _15995_ (.A(_07972_),
    .B(_07856_),
    .C(_07959_),
    .D(_08069_),
    .X(_08609_));
 sky130_fd_sc_hd__o21a_1 _15996_ (.A1(_08325_),
    .A2(_08608_),
    .B1(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__xnor2_1 _15997_ (.A(_08607_),
    .B(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__a22oi_2 _15998_ (.A1(_08209_),
    .A2(_08325_),
    .B1(_08327_),
    .B2(_08193_),
    .Y(_08612_));
 sky130_fd_sc_hd__xnor2_1 _15999_ (.A(_08611_),
    .B(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__and2_1 _16000_ (.A(_07269_),
    .B(_08316_),
    .X(_08614_));
 sky130_fd_sc_hd__xnor2_1 _16001_ (.A(_08613_),
    .B(_08614_),
    .Y(_08615_));
 sky130_fd_sc_hd__inv_2 _16002_ (.A(_08339_),
    .Y(_08616_));
 sky130_fd_sc_hd__a22o_1 _16003_ (.A1(_08227_),
    .A2(_08616_),
    .B1(_08340_),
    .B2(_08206_),
    .X(_08617_));
 sky130_fd_sc_hd__or2_1 _16004_ (.A(_08233_),
    .B(_08359_),
    .X(_08618_));
 sky130_fd_sc_hd__or4_1 _16005_ (.A(_07097_),
    .B(_07084_),
    .C(_07332_),
    .D(_07786_),
    .X(_08619_));
 sky130_fd_sc_hd__o21ai_1 _16006_ (.A1(_07084_),
    .A2(_07787_),
    .B1(_08339_),
    .Y(_08620_));
 sky130_fd_sc_hd__nand2_1 _16007_ (.A(_08619_),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__nor2_1 _16008_ (.A(_07865_),
    .B(_08081_),
    .Y(_08622_));
 sky130_fd_sc_hd__xor2_1 _16009_ (.A(_08621_),
    .B(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__a21oi_1 _16010_ (.A1(_08618_),
    .A2(_08362_),
    .B1(_08623_),
    .Y(_08624_));
 sky130_fd_sc_hd__and3_1 _16011_ (.A(_08618_),
    .B(_08362_),
    .C(_08623_),
    .X(_08625_));
 sky130_fd_sc_hd__nor2_1 _16012_ (.A(_08624_),
    .B(_08625_),
    .Y(_08626_));
 sky130_fd_sc_hd__xnor2_1 _16013_ (.A(_08617_),
    .B(_08626_),
    .Y(_08627_));
 sky130_fd_sc_hd__a21oi_1 _16014_ (.A1(_08336_),
    .A2(_08345_),
    .B1(_08343_),
    .Y(_08628_));
 sky130_fd_sc_hd__nor2_1 _16015_ (.A(_08627_),
    .B(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__and2_1 _16016_ (.A(_08627_),
    .B(_08628_),
    .X(_08630_));
 sky130_fd_sc_hd__nor2_1 _16017_ (.A(_08629_),
    .B(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__xnor2_1 _16018_ (.A(_08615_),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__a21o_1 _16019_ (.A1(_08605_),
    .A2(_08606_),
    .B1(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__nand3_1 _16020_ (.A(_08605_),
    .B(_08606_),
    .C(_08632_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand2_1 _16021_ (.A(_08633_),
    .B(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__xnor2_1 _16022_ (.A(_08604_),
    .B(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__o21ai_1 _16023_ (.A1(_08370_),
    .A2(_08371_),
    .B1(_08373_),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_1 _16024_ (.A(_08379_),
    .B(_08384_),
    .Y(_08638_));
 sky130_fd_sc_hd__or2_1 _16025_ (.A(_06875_),
    .B(_07123_),
    .X(_08639_));
 sky130_fd_sc_hd__or4_2 _16026_ (.A(_06856_),
    .B(_06874_),
    .C(_07141_),
    .D(_07092_),
    .X(_08640_));
 sky130_fd_sc_hd__a21bo_1 _16027_ (.A1(_08359_),
    .A2(_08639_),
    .B1_N(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__or3_1 _16028_ (.A(_07735_),
    .B(_07270_),
    .C(_08641_),
    .X(_08642_));
 sky130_fd_sc_hd__buf_2 _16029_ (.A(_07735_),
    .X(_08643_));
 sky130_fd_sc_hd__o21ai_1 _16030_ (.A1(_08643_),
    .A2(_07857_),
    .B1(_08641_),
    .Y(_08644_));
 sky130_fd_sc_hd__and2_1 _16031_ (.A(_08642_),
    .B(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__or2_1 _16032_ (.A(_08229_),
    .B(_07137_),
    .X(_08646_));
 sky130_fd_sc_hd__or2_1 _16033_ (.A(_07273_),
    .B(_07198_),
    .X(_08647_));
 sky130_fd_sc_hd__or3_1 _16034_ (.A(_07494_),
    .B(_07137_),
    .C(_08647_),
    .X(_08648_));
 sky130_fd_sc_hd__a21bo_1 _16035_ (.A1(_08366_),
    .A2(_08646_),
    .B1_N(_08648_),
    .X(_08649_));
 sky130_fd_sc_hd__or2_1 _16036_ (.A(_07281_),
    .B(_07138_),
    .X(_08650_));
 sky130_fd_sc_hd__xnor2_1 _16037_ (.A(_08649_),
    .B(_08650_),
    .Y(_08651_));
 sky130_fd_sc_hd__a21boi_1 _16038_ (.A1(_08365_),
    .A2(_08368_),
    .B1_N(_08367_),
    .Y(_08652_));
 sky130_fd_sc_hd__nor2_1 _16039_ (.A(_08651_),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__and2_1 _16040_ (.A(_08651_),
    .B(_08652_),
    .X(_08654_));
 sky130_fd_sc_hd__nor2_1 _16041_ (.A(_08653_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__xnor2_1 _16042_ (.A(_08645_),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__a21o_1 _16043_ (.A1(_08638_),
    .A2(_08386_),
    .B1(_08656_),
    .X(_08657_));
 sky130_fd_sc_hd__nand3_1 _16044_ (.A(_08638_),
    .B(_08386_),
    .C(_08656_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(_08657_),
    .B(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__xnor2_2 _16046_ (.A(_08637_),
    .B(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__o21ba_1 _16047_ (.A1(_08249_),
    .A2(_08382_),
    .B1_N(_08381_),
    .X(_08661_));
 sky130_fd_sc_hd__a2bb2o_1 _16048_ (.A1_N(_08265_),
    .A2_N(_08392_),
    .B1(_08393_),
    .B2(_08389_),
    .X(_08662_));
 sky130_fd_sc_hd__or4_1 _16049_ (.A(_07581_),
    .B(_07530_),
    .C(_07756_),
    .D(_07757_),
    .X(_08663_));
 sky130_fd_sc_hd__o21ai_1 _16050_ (.A1(_07530_),
    .A2(_08133_),
    .B1(_08380_),
    .Y(_08664_));
 sky130_fd_sc_hd__nand2_1 _16051_ (.A(_08663_),
    .B(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__nor2_1 _16052_ (.A(_06997_),
    .B(_08130_),
    .Y(_08666_));
 sky130_fd_sc_hd__xnor2_1 _16053_ (.A(_08665_),
    .B(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__nand2_1 _16054_ (.A(_08662_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__or2_1 _16055_ (.A(_08662_),
    .B(_08667_),
    .X(_08669_));
 sky130_fd_sc_hd__and2_1 _16056_ (.A(_08668_),
    .B(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__xnor2_2 _16057_ (.A(_08661_),
    .B(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__nor2_1 _16058_ (.A(_07877_),
    .B(_08260_),
    .Y(_08672_));
 sky130_fd_sc_hd__or4_1 _16059_ (.A(_07661_),
    .B(_07662_),
    .C(_08018_),
    .D(_08391_),
    .X(_08673_));
 sky130_fd_sc_hd__o21ai_1 _16060_ (.A1(_07661_),
    .A2(_08018_),
    .B1(_08392_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand2_1 _16061_ (.A(_08673_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__xnor2_1 _16062_ (.A(_08672_),
    .B(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__a21oi_1 _16063_ (.A1(_03493_),
    .A2(\rbzero.wall_tracer.stepDistY[9] ),
    .B1(_04950_),
    .Y(_08677_));
 sky130_fd_sc_hd__a2bb2o_4 _16064_ (.A1_N(_04841_),
    .A2_N(\rbzero.wall_tracer.stepDistX[9] ),
    .B1(_08269_),
    .B2(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__o31a_1 _16065_ (.A1(_07199_),
    .A2(_08678_),
    .A3(_08402_),
    .B1(_08400_),
    .X(_08679_));
 sky130_fd_sc_hd__or2_1 _16066_ (.A(_07213_),
    .B(_08678_),
    .X(_08680_));
 sky130_fd_sc_hd__or2_2 _16067_ (.A(_08396_),
    .B(_08399_),
    .X(_08681_));
 sky130_fd_sc_hd__or4_2 _16068_ (.A(_07195_),
    .B(_04950_),
    .C(_07185_),
    .D(_08399_),
    .X(_08682_));
 sky130_fd_sc_hd__nand2_1 _16069_ (.A(_07185_),
    .B(_07199_),
    .Y(_08683_));
 sky130_fd_sc_hd__and3b_1 _16070_ (.A_N(_08681_),
    .B(_08682_),
    .C(_08683_),
    .X(_08684_));
 sky130_fd_sc_hd__mux2_1 _16071_ (.A0(_08680_),
    .A1(_07673_),
    .S(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__xor2_1 _16072_ (.A(_08679_),
    .B(_08685_),
    .X(_08686_));
 sky130_fd_sc_hd__xnor2_1 _16073_ (.A(_08676_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__nand2_1 _16074_ (.A(_08403_),
    .B(_08405_),
    .Y(_08688_));
 sky130_fd_sc_hd__a21boi_1 _16075_ (.A1(_08395_),
    .A2(_08406_),
    .B1_N(_08688_),
    .Y(_08689_));
 sky130_fd_sc_hd__nor2_1 _16076_ (.A(_08687_),
    .B(_08689_),
    .Y(_08690_));
 sky130_fd_sc_hd__nand2_1 _16077_ (.A(_08687_),
    .B(_08689_),
    .Y(_08691_));
 sky130_fd_sc_hd__and2b_1 _16078_ (.A_N(_08690_),
    .B(_08691_),
    .X(_08692_));
 sky130_fd_sc_hd__xnor2_2 _16079_ (.A(_08671_),
    .B(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__nor2_1 _16080_ (.A(_08407_),
    .B(_08409_),
    .Y(_08694_));
 sky130_fd_sc_hd__a21oi_2 _16081_ (.A1(_08388_),
    .A2(_08410_),
    .B1(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__xor2_2 _16082_ (.A(_08693_),
    .B(_08695_),
    .X(_08696_));
 sky130_fd_sc_hd__xnor2_2 _16083_ (.A(_08660_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__a21oi_2 _16084_ (.A1(_08377_),
    .A2(_08414_),
    .B1(_08413_),
    .Y(_08698_));
 sky130_fd_sc_hd__nor2_1 _16085_ (.A(_08697_),
    .B(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(_08697_),
    .B(_08698_),
    .Y(_08700_));
 sky130_fd_sc_hd__and2b_1 _16087_ (.A_N(_08699_),
    .B(_08700_),
    .X(_08701_));
 sky130_fd_sc_hd__xor2_1 _16088_ (.A(_08636_),
    .B(_08701_),
    .X(_08702_));
 sky130_fd_sc_hd__a21o_1 _16089_ (.A1(_08355_),
    .A2(_08419_),
    .B1(_08417_),
    .X(_08703_));
 sky130_fd_sc_hd__xor2_1 _16090_ (.A(_08702_),
    .B(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__and2_1 _16091_ (.A(_08603_),
    .B(_08704_),
    .X(_08705_));
 sky130_fd_sc_hd__nor2_1 _16092_ (.A(_08603_),
    .B(_08704_),
    .Y(_08706_));
 sky130_fd_sc_hd__or2_1 _16093_ (.A(_08705_),
    .B(_08706_),
    .X(_08707_));
 sky130_fd_sc_hd__a21oi_1 _16094_ (.A1(_08320_),
    .A2(_08423_),
    .B1(_08421_),
    .Y(_08708_));
 sky130_fd_sc_hd__xor2_1 _16095_ (.A(_08707_),
    .B(_08708_),
    .X(_08709_));
 sky130_fd_sc_hd__xor2_1 _16096_ (.A(_08598_),
    .B(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(_08427_),
    .B(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__or2_1 _16098_ (.A(_08427_),
    .B(_08710_),
    .X(_08712_));
 sky130_fd_sc_hd__nand2_2 _16099_ (.A(_08711_),
    .B(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__nand2_1 _16100_ (.A(_08294_),
    .B(_08297_),
    .Y(_08714_));
 sky130_fd_sc_hd__a32oi_4 _16101_ (.A1(_08299_),
    .A2(_08302_),
    .A3(_08430_),
    .B1(_08714_),
    .B2(_08429_),
    .Y(_08715_));
 sky130_fd_sc_hd__xor2_2 _16102_ (.A(_08713_),
    .B(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__nand2_1 _16103_ (.A(_04946_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__o311a_1 _16104_ (.A1(_08485_),
    .A2(_08595_),
    .A3(_08596_),
    .B1(_08507_),
    .C1(_08717_),
    .X(_08718_));
 sky130_fd_sc_hd__a21oi_1 _16105_ (.A1(_04966_),
    .A2(_08489_),
    .B1(_08718_),
    .Y(_00549_));
 sky130_fd_sc_hd__or2_1 _16106_ (.A(_08707_),
    .B(_08708_),
    .X(_08719_));
 sky130_fd_sc_hd__nand2_1 _16107_ (.A(_08598_),
    .B(_08709_),
    .Y(_08720_));
 sky130_fd_sc_hd__nand2_2 _16108_ (.A(_08719_),
    .B(_08720_),
    .Y(_08721_));
 sky130_fd_sc_hd__or2b_1 _16109_ (.A(_08635_),
    .B_N(_08604_),
    .X(_08722_));
 sky130_fd_sc_hd__or2b_1 _16110_ (.A(_08613_),
    .B_N(_08614_),
    .X(_08723_));
 sky130_fd_sc_hd__o21a_1 _16111_ (.A1(_08611_),
    .A2(_08612_),
    .B1(_08723_),
    .X(_08724_));
 sky130_fd_sc_hd__a21oi_4 _16112_ (.A1(_08633_),
    .A2(_08722_),
    .B1(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__and3_1 _16113_ (.A(_08633_),
    .B(_08722_),
    .C(_08724_),
    .X(_08726_));
 sky130_fd_sc_hd__nor2_1 _16114_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__a21o_1 _16115_ (.A1(_08615_),
    .A2(_08631_),
    .B1(_08629_),
    .X(_08728_));
 sky130_fd_sc_hd__or2b_1 _16116_ (.A(_08659_),
    .B_N(_08637_),
    .X(_08729_));
 sky130_fd_sc_hd__nor2_1 _16117_ (.A(_07856_),
    .B(_08191_),
    .Y(_08730_));
 sky130_fd_sc_hd__or4_1 _16118_ (.A(_07235_),
    .B(_07972_),
    .C(_07959_),
    .D(_08069_),
    .X(_08731_));
 sky130_fd_sc_hd__inv_2 _16119_ (.A(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__o22a_1 _16120_ (.A1(_07865_),
    .A2(_07959_),
    .B1(_08070_),
    .B2(_07972_),
    .X(_08733_));
 sky130_fd_sc_hd__nor2_1 _16121_ (.A(_08732_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__xnor2_1 _16122_ (.A(_08730_),
    .B(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__a21boi_1 _16123_ (.A1(_08607_),
    .A2(_08610_),
    .B1_N(_08609_),
    .Y(_08736_));
 sky130_fd_sc_hd__xor2_1 _16124_ (.A(_08735_),
    .B(_08736_),
    .X(_08737_));
 sky130_fd_sc_hd__and2_1 _16125_ (.A(_07265_),
    .B(_08316_),
    .X(_08738_));
 sky130_fd_sc_hd__nand2_1 _16126_ (.A(_08737_),
    .B(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__or2_1 _16127_ (.A(_08737_),
    .B(_08738_),
    .X(_08740_));
 sky130_fd_sc_hd__and2_1 _16128_ (.A(_08739_),
    .B(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__a21bo_1 _16129_ (.A1(_08620_),
    .A2(_08622_),
    .B1_N(_08619_),
    .X(_08742_));
 sky130_fd_sc_hd__nor2_1 _16130_ (.A(_08107_),
    .B(_07787_),
    .Y(_08743_));
 sky130_fd_sc_hd__nor2_1 _16131_ (.A(_07735_),
    .B(_07332_),
    .Y(_08744_));
 sky130_fd_sc_hd__or3_1 _16132_ (.A(_07735_),
    .B(_07786_),
    .C(_08339_),
    .X(_08745_));
 sky130_fd_sc_hd__o21a_1 _16133_ (.A1(_08743_),
    .A2(_08744_),
    .B1(_08745_),
    .X(_08746_));
 sky130_fd_sc_hd__nor2_1 _16134_ (.A(_07984_),
    .B(_08081_),
    .Y(_08747_));
 sky130_fd_sc_hd__xnor2_1 _16135_ (.A(_08746_),
    .B(_08747_),
    .Y(_08748_));
 sky130_fd_sc_hd__a21o_1 _16136_ (.A1(_08640_),
    .A2(_08642_),
    .B1(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__nand3_1 _16137_ (.A(_08640_),
    .B(_08642_),
    .C(_08748_),
    .Y(_08750_));
 sky130_fd_sc_hd__and2_1 _16138_ (.A(_08749_),
    .B(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__nand2_1 _16139_ (.A(_08742_),
    .B(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__or2_1 _16140_ (.A(_08742_),
    .B(_08751_),
    .X(_08753_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(_08752_),
    .B(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__a21oi_1 _16142_ (.A1(_08617_),
    .A2(_08626_),
    .B1(_08624_),
    .Y(_08755_));
 sky130_fd_sc_hd__nor2_1 _16143_ (.A(_08754_),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__and2_1 _16144_ (.A(_08754_),
    .B(_08755_),
    .X(_08757_));
 sky130_fd_sc_hd__nor2_1 _16145_ (.A(_08756_),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__xnor2_1 _16146_ (.A(_08741_),
    .B(_08758_),
    .Y(_08759_));
 sky130_fd_sc_hd__a21o_1 _16147_ (.A1(_08657_),
    .A2(_08729_),
    .B1(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__nand3_1 _16148_ (.A(_08657_),
    .B(_08729_),
    .C(_08759_),
    .Y(_08761_));
 sky130_fd_sc_hd__nand2_1 _16149_ (.A(_08760_),
    .B(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__xnor2_1 _16150_ (.A(_08728_),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__a21o_1 _16151_ (.A1(_08645_),
    .A2(_08655_),
    .B1(_08653_),
    .X(_08764_));
 sky130_fd_sc_hd__or2b_1 _16152_ (.A(_08661_),
    .B_N(_08670_),
    .X(_08765_));
 sky130_fd_sc_hd__and2_1 _16153_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_07256_),
    .X(_08766_));
 sky130_fd_sc_hd__inv_2 _16154_ (.A(_08000_),
    .Y(_08767_));
 sky130_fd_sc_hd__nor2_1 _16155_ (.A(_07012_),
    .B(_07878_),
    .Y(_08768_));
 sky130_fd_sc_hd__o22a_1 _16156_ (.A1(_06858_),
    .A2(_07878_),
    .B1(_08000_),
    .B2(_07012_),
    .X(_08769_));
 sky130_fd_sc_hd__a31o_1 _16157_ (.A1(_08766_),
    .A2(_08767_),
    .A3(_08768_),
    .B1(_08769_),
    .X(_08770_));
 sky130_fd_sc_hd__nor2_1 _16158_ (.A(_07993_),
    .B(_07857_),
    .Y(_08771_));
 sky130_fd_sc_hd__xnor2_1 _16159_ (.A(_08770_),
    .B(_08771_),
    .Y(_08772_));
 sky130_fd_sc_hd__or2_1 _16160_ (.A(_07494_),
    .B(_08130_),
    .X(_08773_));
 sky130_fd_sc_hd__or3_1 _16161_ (.A(_08229_),
    .B(_07748_),
    .C(_08366_),
    .X(_08774_));
 sky130_fd_sc_hd__a21bo_1 _16162_ (.A1(_08647_),
    .A2(_08773_),
    .B1_N(_08774_),
    .X(_08775_));
 sky130_fd_sc_hd__or2_1 _16163_ (.A(_08108_),
    .B(_08252_),
    .X(_08776_));
 sky130_fd_sc_hd__xnor2_1 _16164_ (.A(_08775_),
    .B(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__o31a_1 _16165_ (.A1(_08108_),
    .A2(_07878_),
    .A3(_08649_),
    .B1(_08648_),
    .X(_08778_));
 sky130_fd_sc_hd__nor2_1 _16166_ (.A(_08777_),
    .B(_08778_),
    .Y(_08779_));
 sky130_fd_sc_hd__and2_1 _16167_ (.A(_08777_),
    .B(_08778_),
    .X(_08780_));
 sky130_fd_sc_hd__nor2_1 _16168_ (.A(_08779_),
    .B(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__xnor2_1 _16169_ (.A(_08772_),
    .B(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__a21o_1 _16170_ (.A1(_08668_),
    .A2(_08765_),
    .B1(_08782_),
    .X(_08783_));
 sky130_fd_sc_hd__nand3_1 _16171_ (.A(_08668_),
    .B(_08765_),
    .C(_08782_),
    .Y(_08784_));
 sky130_fd_sc_hd__nand2_1 _16172_ (.A(_08783_),
    .B(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__xnor2_1 _16173_ (.A(_08764_),
    .B(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__a21bo_1 _16174_ (.A1(_08664_),
    .A2(_08666_),
    .B1_N(_08663_),
    .X(_08787_));
 sky130_fd_sc_hd__a21bo_1 _16175_ (.A1(_08672_),
    .A2(_08674_),
    .B1_N(_08673_),
    .X(_08788_));
 sky130_fd_sc_hd__nor3_1 _16176_ (.A(_08245_),
    .B(_08260_),
    .C(_08380_),
    .Y(_08789_));
 sky130_fd_sc_hd__o22a_1 _16177_ (.A1(_08245_),
    .A2(_08134_),
    .B1(_08260_),
    .B2(_08247_),
    .X(_08790_));
 sky130_fd_sc_hd__nor2_1 _16178_ (.A(_08789_),
    .B(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__nor2_1 _16179_ (.A(_07992_),
    .B(_08133_),
    .Y(_08792_));
 sky130_fd_sc_hd__xor2_1 _16180_ (.A(_08791_),
    .B(_08792_),
    .X(_08793_));
 sky130_fd_sc_hd__nand2_1 _16181_ (.A(_08788_),
    .B(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__or2_1 _16182_ (.A(_08788_),
    .B(_08793_),
    .X(_08795_));
 sky130_fd_sc_hd__and2_1 _16183_ (.A(_08794_),
    .B(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__xor2_2 _16184_ (.A(_08787_),
    .B(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_07877_),
    .B(_08018_),
    .Y(_08798_));
 sky130_fd_sc_hd__or2_1 _16186_ (.A(_07661_),
    .B(_08678_),
    .X(_08799_));
 sky130_fd_sc_hd__o22ai_1 _16187_ (.A1(_07661_),
    .A2(_08391_),
    .B1(_08678_),
    .B2(_07662_),
    .Y(_08800_));
 sky130_fd_sc_hd__o21ai_1 _16188_ (.A1(_08392_),
    .A2(_08799_),
    .B1(_08800_),
    .Y(_08801_));
 sky130_fd_sc_hd__xnor2_1 _16189_ (.A(_08798_),
    .B(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__clkbuf_4 _16190_ (.A(_08681_),
    .X(_08803_));
 sky130_fd_sc_hd__a31o_1 _16191_ (.A1(_07213_),
    .A2(_07185_),
    .A3(_07199_),
    .B1(_08803_),
    .X(_08804_));
 sky130_fd_sc_hd__or2_2 _16192_ (.A(_07213_),
    .B(_08682_),
    .X(_08805_));
 sky130_fd_sc_hd__and2b_1 _16193_ (.A_N(_08804_),
    .B(_08805_),
    .X(_08806_));
 sky130_fd_sc_hd__buf_2 _16194_ (.A(_08806_),
    .X(_08807_));
 sky130_fd_sc_hd__xnor2_1 _16195_ (.A(_08802_),
    .B(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__nor2_1 _16196_ (.A(_08679_),
    .B(_08685_),
    .Y(_08809_));
 sky130_fd_sc_hd__a21o_1 _16197_ (.A1(_08676_),
    .A2(_08686_),
    .B1(_08809_),
    .X(_08810_));
 sky130_fd_sc_hd__xnor2_1 _16198_ (.A(_08808_),
    .B(_08810_),
    .Y(_08811_));
 sky130_fd_sc_hd__xnor2_2 _16199_ (.A(_08797_),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__a21oi_2 _16200_ (.A1(_08671_),
    .A2(_08691_),
    .B1(_08690_),
    .Y(_08813_));
 sky130_fd_sc_hd__xor2_1 _16201_ (.A(_08812_),
    .B(_08813_),
    .X(_08814_));
 sky130_fd_sc_hd__nand2_1 _16202_ (.A(_08786_),
    .B(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__or2_1 _16203_ (.A(_08786_),
    .B(_08814_),
    .X(_08816_));
 sky130_fd_sc_hd__nand2_1 _16204_ (.A(_08815_),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__nor2_1 _16205_ (.A(_08693_),
    .B(_08695_),
    .Y(_08818_));
 sky130_fd_sc_hd__a21oi_2 _16206_ (.A1(_08660_),
    .A2(_08696_),
    .B1(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__xor2_1 _16207_ (.A(_08817_),
    .B(_08819_),
    .X(_08820_));
 sky130_fd_sc_hd__xnor2_1 _16208_ (.A(_08763_),
    .B(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__a21oi_1 _16209_ (.A1(_08636_),
    .A2(_08700_),
    .B1(_08699_),
    .Y(_08822_));
 sky130_fd_sc_hd__nor2_1 _16210_ (.A(_08821_),
    .B(_08822_),
    .Y(_08823_));
 sky130_fd_sc_hd__nand2_1 _16211_ (.A(_08821_),
    .B(_08822_),
    .Y(_08824_));
 sky130_fd_sc_hd__and2b_1 _16212_ (.A_N(_08823_),
    .B(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__xnor2_1 _16213_ (.A(_08727_),
    .B(_08825_),
    .Y(_08826_));
 sky130_fd_sc_hd__a21oi_1 _16214_ (.A1(_08702_),
    .A2(_08703_),
    .B1(_08705_),
    .Y(_08827_));
 sky130_fd_sc_hd__xor2_1 _16215_ (.A(_08826_),
    .B(_08827_),
    .X(_08828_));
 sky130_fd_sc_hd__nand2_1 _16216_ (.A(_08601_),
    .B(_08828_),
    .Y(_08829_));
 sky130_fd_sc_hd__or2_1 _16217_ (.A(_08601_),
    .B(_08828_),
    .X(_08830_));
 sky130_fd_sc_hd__nand2_2 _16218_ (.A(_08829_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__xor2_4 _16219_ (.A(_08721_),
    .B(_08831_),
    .X(_08832_));
 sky130_fd_sc_hd__o21ai_2 _16220_ (.A1(_08713_),
    .A2(_08715_),
    .B1(_08711_),
    .Y(_08833_));
 sky130_fd_sc_hd__xnor2_4 _16221_ (.A(_08832_),
    .B(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__and2_1 _16222_ (.A(_08524_),
    .B(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__nand2_1 _16223_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_08836_));
 sky130_fd_sc_hd__or2_1 _16224_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_08837_));
 sky130_fd_sc_hd__o211a_1 _16225_ (.A1(_08592_),
    .A2(_08596_),
    .B1(_08836_),
    .C1(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__inv_2 _16226_ (.A(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__a211o_1 _16227_ (.A1(_08836_),
    .A2(_08837_),
    .B1(_08592_),
    .C1(_08596_),
    .X(_08840_));
 sky130_fd_sc_hd__a31o_1 _16228_ (.A1(_08562_),
    .A2(_08839_),
    .A3(_08840_),
    .B1(_08522_),
    .X(_08841_));
 sky130_fd_sc_hd__o22a_1 _16229_ (.A1(\rbzero.wall_tracer.trackDistX[1] ),
    .A2(_08553_),
    .B1(_08835_),
    .B2(_08841_),
    .X(_00550_));
 sky130_fd_sc_hd__or2b_1 _16230_ (.A(_08762_),
    .B_N(_08728_),
    .X(_08842_));
 sky130_fd_sc_hd__o21a_1 _16231_ (.A1(_08735_),
    .A2(_08736_),
    .B1(_08739_),
    .X(_08843_));
 sky130_fd_sc_hd__a21oi_2 _16232_ (.A1(_08760_),
    .A2(_08842_),
    .B1(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__and3_1 _16233_ (.A(_08760_),
    .B(_08842_),
    .C(_08843_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _16234_ (.A(_08844_),
    .B(_08845_),
    .Y(_08846_));
 sky130_fd_sc_hd__a21o_1 _16235_ (.A1(_08741_),
    .A2(_08758_),
    .B1(_08756_),
    .X(_08847_));
 sky130_fd_sc_hd__or2b_1 _16236_ (.A(_08785_),
    .B_N(_08764_),
    .X(_08848_));
 sky130_fd_sc_hd__nor2_1 _16237_ (.A(_07972_),
    .B(_08191_),
    .Y(_08849_));
 sky130_fd_sc_hd__or4_1 _16238_ (.A(_07984_),
    .B(_07865_),
    .C(_07959_),
    .D(_08070_),
    .X(_08850_));
 sky130_fd_sc_hd__inv_2 _16239_ (.A(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__o22a_1 _16240_ (.A1(_07984_),
    .A2(_07960_),
    .B1(_08070_),
    .B2(_07865_),
    .X(_08852_));
 sky130_fd_sc_hd__nor2_1 _16241_ (.A(_08851_),
    .B(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__xnor2_1 _16242_ (.A(_08849_),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__a21oi_1 _16243_ (.A1(_08730_),
    .A2(_08734_),
    .B1(_08732_),
    .Y(_08855_));
 sky130_fd_sc_hd__nor2_1 _16244_ (.A(_08854_),
    .B(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__and2_1 _16245_ (.A(_08854_),
    .B(_08855_),
    .X(_08857_));
 sky130_fd_sc_hd__nor2_1 _16246_ (.A(_08856_),
    .B(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__and2_1 _16247_ (.A(_07856_),
    .B(_08316_),
    .X(_08859_));
 sky130_fd_sc_hd__xor2_1 _16248_ (.A(_08858_),
    .B(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__a21bo_1 _16249_ (.A1(_08746_),
    .A2(_08747_),
    .B1_N(_08745_),
    .X(_08861_));
 sky130_fd_sc_hd__clkbuf_4 _16250_ (.A(_07878_),
    .X(_08862_));
 sky130_fd_sc_hd__or3_1 _16251_ (.A(_07012_),
    .B(_08862_),
    .C(_08359_),
    .X(_08863_));
 sky130_fd_sc_hd__o31ai_1 _16252_ (.A1(_07993_),
    .A2(_07857_),
    .A3(_08769_),
    .B1(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__or2_1 _16253_ (.A(_07123_),
    .B(_07787_),
    .X(_08865_));
 sky130_fd_sc_hd__or3_1 _16254_ (.A(_07735_),
    .B(_07333_),
    .C(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__o22ai_1 _16255_ (.A1(_07993_),
    .A2(_07333_),
    .B1(_07787_),
    .B2(_08643_),
    .Y(_08867_));
 sky130_fd_sc_hd__nand2_1 _16256_ (.A(_08866_),
    .B(_08867_),
    .Y(_08868_));
 sky130_fd_sc_hd__nor2_1 _16257_ (.A(_08107_),
    .B(_08081_),
    .Y(_08869_));
 sky130_fd_sc_hd__xnor2_1 _16258_ (.A(_08868_),
    .B(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__and2_1 _16259_ (.A(_08864_),
    .B(_08870_),
    .X(_08871_));
 sky130_fd_sc_hd__nor2_1 _16260_ (.A(_08864_),
    .B(_08870_),
    .Y(_08872_));
 sky130_fd_sc_hd__nor2_1 _16261_ (.A(_08871_),
    .B(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__xnor2_1 _16262_ (.A(_08861_),
    .B(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__a21oi_1 _16263_ (.A1(_08749_),
    .A2(_08752_),
    .B1(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__and3_1 _16264_ (.A(_08749_),
    .B(_08752_),
    .C(_08874_),
    .X(_08876_));
 sky130_fd_sc_hd__nor2_1 _16265_ (.A(_08875_),
    .B(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__xnor2_1 _16266_ (.A(_08860_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__a21o_1 _16267_ (.A1(_08783_),
    .A2(_08848_),
    .B1(_08878_),
    .X(_08879_));
 sky130_fd_sc_hd__nand3_1 _16268_ (.A(_08783_),
    .B(_08848_),
    .C(_08878_),
    .Y(_08880_));
 sky130_fd_sc_hd__nand2_1 _16269_ (.A(_08879_),
    .B(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__xnor2_1 _16270_ (.A(_08847_),
    .B(_08881_),
    .Y(_08882_));
 sky130_fd_sc_hd__a21o_1 _16271_ (.A1(_08772_),
    .A2(_08781_),
    .B1(_08779_),
    .X(_08883_));
 sky130_fd_sc_hd__nand2_1 _16272_ (.A(_08787_),
    .B(_08796_),
    .Y(_08884_));
 sky130_fd_sc_hd__nor2_1 _16273_ (.A(_06858_),
    .B(_08252_),
    .Y(_08885_));
 sky130_fd_sc_hd__or4_1 _16274_ (.A(_06858_),
    .B(_07012_),
    .C(_07878_),
    .D(_08252_),
    .X(_08886_));
 sky130_fd_sc_hd__o21ai_1 _16275_ (.A1(_08768_),
    .A2(_08885_),
    .B1(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__buf_2 _16276_ (.A(_08000_),
    .X(_08888_));
 sky130_fd_sc_hd__clkbuf_4 _16277_ (.A(_07857_),
    .X(_08889_));
 sky130_fd_sc_hd__nor2_1 _16278_ (.A(_08888_),
    .B(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__xnor2_1 _16279_ (.A(_08887_),
    .B(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__or3_1 _16280_ (.A(_08229_),
    .B(_08133_),
    .C(_08773_),
    .X(_08892_));
 sky130_fd_sc_hd__o22a_1 _16281_ (.A1(_08229_),
    .A2(_08130_),
    .B1(_08133_),
    .B2(_07494_),
    .X(_08893_));
 sky130_fd_sc_hd__clkinv_2 _16282_ (.A(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__and2_1 _16283_ (.A(_08892_),
    .B(_08894_),
    .X(_08895_));
 sky130_fd_sc_hd__buf_2 _16284_ (.A(_07766_),
    .X(_08896_));
 sky130_fd_sc_hd__nor2_1 _16285_ (.A(_08108_),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__xnor2_1 _16286_ (.A(_08895_),
    .B(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__buf_2 _16287_ (.A(_08252_),
    .X(_08899_));
 sky130_fd_sc_hd__o31a_1 _16288_ (.A1(_08108_),
    .A2(_08899_),
    .A3(_08775_),
    .B1(_08774_),
    .X(_08900_));
 sky130_fd_sc_hd__nor2_1 _16289_ (.A(_08898_),
    .B(_08900_),
    .Y(_08901_));
 sky130_fd_sc_hd__and2_1 _16290_ (.A(_08898_),
    .B(_08900_),
    .X(_08902_));
 sky130_fd_sc_hd__nor2_1 _16291_ (.A(_08901_),
    .B(_08902_),
    .Y(_08903_));
 sky130_fd_sc_hd__xnor2_1 _16292_ (.A(_08891_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__a21o_1 _16293_ (.A1(_08794_),
    .A2(_08884_),
    .B1(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__nand3_1 _16294_ (.A(_08794_),
    .B(_08884_),
    .C(_08904_),
    .Y(_08906_));
 sky130_fd_sc_hd__nand2_1 _16295_ (.A(_08905_),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__xnor2_1 _16296_ (.A(_08883_),
    .B(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__a21o_1 _16297_ (.A1(_08791_),
    .A2(_08792_),
    .B1(_08789_),
    .X(_08909_));
 sky130_fd_sc_hd__a2bb2o_1 _16298_ (.A1_N(_08392_),
    .A2_N(_08799_),
    .B1(_08800_),
    .B2(_08798_),
    .X(_08910_));
 sky130_fd_sc_hd__nor2_1 _16299_ (.A(_07581_),
    .B(_07897_),
    .Y(_08911_));
 sky130_fd_sc_hd__or3b_1 _16300_ (.A(_07530_),
    .B(_08018_),
    .C_N(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__o22ai_1 _16301_ (.A1(_08245_),
    .A2(_08260_),
    .B1(_08018_),
    .B2(_08247_),
    .Y(_08913_));
 sky130_fd_sc_hd__nand2_1 _16302_ (.A(_08912_),
    .B(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__nor2_1 _16303_ (.A(_06997_),
    .B(_08134_),
    .Y(_08915_));
 sky130_fd_sc_hd__xnor2_1 _16304_ (.A(_08914_),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand2_1 _16305_ (.A(_08910_),
    .B(_08916_),
    .Y(_08917_));
 sky130_fd_sc_hd__or2_1 _16306_ (.A(_08910_),
    .B(_08916_),
    .X(_08918_));
 sky130_fd_sc_hd__and2_1 _16307_ (.A(_08917_),
    .B(_08918_),
    .X(_08919_));
 sky130_fd_sc_hd__nand2_1 _16308_ (.A(_08909_),
    .B(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__or2_1 _16309_ (.A(_08909_),
    .B(_08919_),
    .X(_08921_));
 sky130_fd_sc_hd__and2_1 _16310_ (.A(_08920_),
    .B(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__or2_1 _16311_ (.A(_07877_),
    .B(_08391_),
    .X(_08923_));
 sky130_fd_sc_hd__nor2_1 _16312_ (.A(_07662_),
    .B(_08803_),
    .Y(_08924_));
 sky130_fd_sc_hd__xor2_1 _16313_ (.A(_08799_),
    .B(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__xor2_1 _16314_ (.A(_08923_),
    .B(_08925_),
    .X(_08926_));
 sky130_fd_sc_hd__xnor2_1 _16315_ (.A(_08807_),
    .B(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__a21boi_1 _16316_ (.A1(_08802_),
    .A2(_08807_),
    .B1_N(_08805_),
    .Y(_08928_));
 sky130_fd_sc_hd__nor2_1 _16317_ (.A(_08927_),
    .B(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__and2_1 _16318_ (.A(_08927_),
    .B(_08928_),
    .X(_08930_));
 sky130_fd_sc_hd__nor2_1 _16319_ (.A(_08929_),
    .B(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__xnor2_1 _16320_ (.A(_08922_),
    .B(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__and2b_1 _16321_ (.A_N(_08808_),
    .B(_08810_),
    .X(_08933_));
 sky130_fd_sc_hd__a21oi_1 _16322_ (.A1(_08797_),
    .A2(_08811_),
    .B1(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__nor2_1 _16323_ (.A(_08932_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__and2_1 _16324_ (.A(_08932_),
    .B(_08934_),
    .X(_08936_));
 sky130_fd_sc_hd__nor2_1 _16325_ (.A(_08935_),
    .B(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__xnor2_1 _16326_ (.A(_08908_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__o21a_1 _16327_ (.A1(_08812_),
    .A2(_08813_),
    .B1(_08815_),
    .X(_08939_));
 sky130_fd_sc_hd__nor2_1 _16328_ (.A(_08938_),
    .B(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__and2_1 _16329_ (.A(_08938_),
    .B(_08939_),
    .X(_08941_));
 sky130_fd_sc_hd__nor2_1 _16330_ (.A(_08940_),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__xnor2_1 _16331_ (.A(_08882_),
    .B(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__nor2_1 _16332_ (.A(_08817_),
    .B(_08819_),
    .Y(_08944_));
 sky130_fd_sc_hd__a21oi_1 _16333_ (.A1(_08763_),
    .A2(_08820_),
    .B1(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__xor2_1 _16334_ (.A(_08943_),
    .B(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__xnor2_1 _16335_ (.A(_08846_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__a21oi_1 _16336_ (.A1(_08727_),
    .A2(_08824_),
    .B1(_08823_),
    .Y(_08948_));
 sky130_fd_sc_hd__nor2_1 _16337_ (.A(_08947_),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__nand2_1 _16338_ (.A(_08947_),
    .B(_08948_),
    .Y(_08950_));
 sky130_fd_sc_hd__and2b_1 _16339_ (.A_N(_08949_),
    .B(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__xnor2_4 _16340_ (.A(_08725_),
    .B(_08951_),
    .Y(_08952_));
 sky130_fd_sc_hd__o21a_2 _16341_ (.A1(_08826_),
    .A2(_08827_),
    .B1(_08829_),
    .X(_08953_));
 sky130_fd_sc_hd__xnor2_4 _16342_ (.A(_08952_),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__a31o_1 _16343_ (.A1(_08719_),
    .A2(_08720_),
    .A3(_08831_),
    .B1(_08711_),
    .X(_08955_));
 sky130_fd_sc_hd__or2b_1 _16344_ (.A(_08831_),
    .B_N(_08721_),
    .X(_08956_));
 sky130_fd_sc_hd__o311ai_4 _16345_ (.A1(_08713_),
    .A2(_08715_),
    .A3(_08832_),
    .B1(_08955_),
    .C1(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__xnor2_4 _16346_ (.A(_08954_),
    .B(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__and2_1 _16347_ (.A(_08524_),
    .B(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__nand2_1 _16348_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .Y(_08960_));
 sky130_fd_sc_hd__or2_1 _16349_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_08961_));
 sky130_fd_sc_hd__nand2_1 _16350_ (.A(_08836_),
    .B(_08839_),
    .Y(_08962_));
 sky130_fd_sc_hd__a21o_1 _16351_ (.A1(_08960_),
    .A2(_08961_),
    .B1(_08962_),
    .X(_08963_));
 sky130_fd_sc_hd__and3_1 _16352_ (.A(_08960_),
    .B(_08961_),
    .C(_08962_),
    .X(_08964_));
 sky130_fd_sc_hd__inv_2 _16353_ (.A(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__a31o_1 _16354_ (.A1(_08562_),
    .A2(_08963_),
    .A3(_08965_),
    .B1(_08522_),
    .X(_08966_));
 sky130_fd_sc_hd__o22a_1 _16355_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_08553_),
    .B1(_08959_),
    .B2(_08966_),
    .X(_00551_));
 sky130_fd_sc_hd__a21o_1 _16356_ (.A1(_08725_),
    .A2(_08950_),
    .B1(_08949_),
    .X(_08967_));
 sky130_fd_sc_hd__or2b_1 _16357_ (.A(_08881_),
    .B_N(_08847_),
    .X(_08968_));
 sky130_fd_sc_hd__a21oi_1 _16358_ (.A1(_08858_),
    .A2(_08859_),
    .B1(_08856_),
    .Y(_08969_));
 sky130_fd_sc_hd__a21oi_1 _16359_ (.A1(_08879_),
    .A2(_08968_),
    .B1(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__and3_1 _16360_ (.A(_08879_),
    .B(_08968_),
    .C(_08969_),
    .X(_08971_));
 sky130_fd_sc_hd__nor2_1 _16361_ (.A(_08970_),
    .B(_08971_),
    .Y(_08972_));
 sky130_fd_sc_hd__a21o_1 _16362_ (.A1(_08860_),
    .A2(_08877_),
    .B1(_08875_),
    .X(_08973_));
 sky130_fd_sc_hd__or2b_1 _16363_ (.A(_08907_),
    .B_N(_08883_),
    .X(_08974_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_07865_),
    .B(_08191_),
    .Y(_08975_));
 sky130_fd_sc_hd__or4_1 _16365_ (.A(_08107_),
    .B(_07984_),
    .C(_07960_),
    .D(_08070_),
    .X(_08976_));
 sky130_fd_sc_hd__o22ai_1 _16366_ (.A1(_08107_),
    .A2(_07960_),
    .B1(_08071_),
    .B2(_07984_),
    .Y(_08977_));
 sky130_fd_sc_hd__nand2_1 _16367_ (.A(_08976_),
    .B(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__xor2_1 _16368_ (.A(_08975_),
    .B(_08978_),
    .X(_08979_));
 sky130_fd_sc_hd__a21oi_1 _16369_ (.A1(_08849_),
    .A2(_08853_),
    .B1(_08851_),
    .Y(_08980_));
 sky130_fd_sc_hd__nor2_1 _16370_ (.A(_08979_),
    .B(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__and2_1 _16371_ (.A(_08979_),
    .B(_08980_),
    .X(_08982_));
 sky130_fd_sc_hd__nor2_1 _16372_ (.A(_08981_),
    .B(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__and2_1 _16373_ (.A(_07972_),
    .B(_08317_),
    .X(_08984_));
 sky130_fd_sc_hd__xor2_1 _16374_ (.A(_08983_),
    .B(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__a21bo_1 _16375_ (.A1(_08867_),
    .A2(_08869_),
    .B1_N(_08866_),
    .X(_08986_));
 sky130_fd_sc_hd__or2_1 _16376_ (.A(_08000_),
    .B(_07333_),
    .X(_08987_));
 sky130_fd_sc_hd__or4_1 _16377_ (.A(_08000_),
    .B(_07123_),
    .C(_07333_),
    .D(_07787_),
    .X(_08988_));
 sky130_fd_sc_hd__a21bo_1 _16378_ (.A1(_08865_),
    .A2(_08987_),
    .B1_N(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__nor2_1 _16379_ (.A(_08643_),
    .B(_08081_),
    .Y(_08990_));
 sky130_fd_sc_hd__xor2_1 _16380_ (.A(_08989_),
    .B(_08990_),
    .X(_08991_));
 sky130_fd_sc_hd__o31ai_1 _16381_ (.A1(_08888_),
    .A2(_08889_),
    .A3(_08887_),
    .B1(_08886_),
    .Y(_08992_));
 sky130_fd_sc_hd__and2b_1 _16382_ (.A_N(_08991_),
    .B(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__and2b_1 _16383_ (.A_N(_08992_),
    .B(_08991_),
    .X(_08994_));
 sky130_fd_sc_hd__nor2_1 _16384_ (.A(_08993_),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__xnor2_1 _16385_ (.A(_08986_),
    .B(_08995_),
    .Y(_08996_));
 sky130_fd_sc_hd__a21oi_1 _16386_ (.A1(_08861_),
    .A2(_08873_),
    .B1(_08871_),
    .Y(_08997_));
 sky130_fd_sc_hd__nor2_1 _16387_ (.A(_08996_),
    .B(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__and2_1 _16388_ (.A(_08996_),
    .B(_08997_),
    .X(_08999_));
 sky130_fd_sc_hd__nor2_1 _16389_ (.A(_08998_),
    .B(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__xnor2_1 _16390_ (.A(_08985_),
    .B(_09000_),
    .Y(_09001_));
 sky130_fd_sc_hd__a21o_1 _16391_ (.A1(_08905_),
    .A2(_08974_),
    .B1(_09001_),
    .X(_09002_));
 sky130_fd_sc_hd__nand3_1 _16392_ (.A(_08905_),
    .B(_08974_),
    .C(_09001_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand2_1 _16393_ (.A(_09002_),
    .B(_09003_),
    .Y(_09004_));
 sky130_fd_sc_hd__xnor2_1 _16394_ (.A(_08973_),
    .B(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__a21o_1 _16395_ (.A1(_08891_),
    .A2(_08903_),
    .B1(_08901_),
    .X(_09006_));
 sky130_fd_sc_hd__buf_2 _16396_ (.A(_07012_),
    .X(_09007_));
 sky130_fd_sc_hd__nor2_1 _16397_ (.A(_09007_),
    .B(_08896_),
    .Y(_09008_));
 sky130_fd_sc_hd__buf_2 _16398_ (.A(_06858_),
    .X(_09009_));
 sky130_fd_sc_hd__o22ai_1 _16399_ (.A1(_09007_),
    .A2(_08899_),
    .B1(_08896_),
    .B2(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__a21bo_1 _16400_ (.A1(_08885_),
    .A2(_09008_),
    .B1_N(_09010_),
    .X(_09011_));
 sky130_fd_sc_hd__nor2_1 _16401_ (.A(_08862_),
    .B(_07857_),
    .Y(_09012_));
 sky130_fd_sc_hd__xnor2_1 _16402_ (.A(_09011_),
    .B(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__buf_2 _16403_ (.A(_07494_),
    .X(_09014_));
 sky130_fd_sc_hd__or4_1 _16404_ (.A(_09014_),
    .B(_08229_),
    .C(_08133_),
    .D(_08134_),
    .X(_09015_));
 sky130_fd_sc_hd__buf_2 _16405_ (.A(_08229_),
    .X(_09016_));
 sky130_fd_sc_hd__o22ai_1 _16406_ (.A1(_09016_),
    .A2(_08133_),
    .B1(_08134_),
    .B2(_09014_),
    .Y(_09017_));
 sky130_fd_sc_hd__nand2_1 _16407_ (.A(_09015_),
    .B(_09017_),
    .Y(_09018_));
 sky130_fd_sc_hd__or2_1 _16408_ (.A(_08108_),
    .B(_08130_),
    .X(_09019_));
 sky130_fd_sc_hd__xnor2_1 _16409_ (.A(_09018_),
    .B(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__clkbuf_4 _16410_ (.A(_08108_),
    .X(_09021_));
 sky130_fd_sc_hd__o31a_1 _16411_ (.A1(_09021_),
    .A2(_08896_),
    .A3(_08893_),
    .B1(_08892_),
    .X(_09022_));
 sky130_fd_sc_hd__nor2_1 _16412_ (.A(_09020_),
    .B(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__and2_1 _16413_ (.A(_09020_),
    .B(_09022_),
    .X(_09024_));
 sky130_fd_sc_hd__nor2_1 _16414_ (.A(_09023_),
    .B(_09024_),
    .Y(_09025_));
 sky130_fd_sc_hd__xnor2_1 _16415_ (.A(_09013_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__a21o_1 _16416_ (.A1(_08917_),
    .A2(_08920_),
    .B1(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__nand3_1 _16417_ (.A(_08917_),
    .B(_08920_),
    .C(_09026_),
    .Y(_09028_));
 sky130_fd_sc_hd__nand2_1 _16418_ (.A(_09027_),
    .B(_09028_),
    .Y(_09029_));
 sky130_fd_sc_hd__xnor2_1 _16419_ (.A(_09006_),
    .B(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__a21bo_1 _16420_ (.A1(_08913_),
    .A2(_08915_),
    .B1_N(_08912_),
    .X(_09031_));
 sky130_fd_sc_hd__or3_1 _16421_ (.A(_07662_),
    .B(_08803_),
    .C(_08799_),
    .X(_09032_));
 sky130_fd_sc_hd__or2_1 _16422_ (.A(_08923_),
    .B(_08925_),
    .X(_09033_));
 sky130_fd_sc_hd__or4_1 _16423_ (.A(_08247_),
    .B(_08245_),
    .C(_08018_),
    .D(_08391_),
    .X(_09034_));
 sky130_fd_sc_hd__clkbuf_4 _16424_ (.A(_08018_),
    .X(_09035_));
 sky130_fd_sc_hd__clkbuf_4 _16425_ (.A(_08391_),
    .X(_09036_));
 sky130_fd_sc_hd__o22ai_1 _16426_ (.A1(_08245_),
    .A2(_09035_),
    .B1(_09036_),
    .B2(_08247_),
    .Y(_09037_));
 sky130_fd_sc_hd__nand2_1 _16427_ (.A(_09034_),
    .B(_09037_),
    .Y(_09038_));
 sky130_fd_sc_hd__clkbuf_4 _16428_ (.A(_08260_),
    .X(_09039_));
 sky130_fd_sc_hd__nor2_1 _16429_ (.A(_07992_),
    .B(_09039_),
    .Y(_09040_));
 sky130_fd_sc_hd__xor2_1 _16430_ (.A(_09038_),
    .B(_09040_),
    .X(_09041_));
 sky130_fd_sc_hd__a21o_1 _16431_ (.A1(_09032_),
    .A2(_09033_),
    .B1(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__nand3_1 _16432_ (.A(_09032_),
    .B(_09033_),
    .C(_09041_),
    .Y(_09043_));
 sky130_fd_sc_hd__and2_1 _16433_ (.A(_09042_),
    .B(_09043_),
    .X(_09044_));
 sky130_fd_sc_hd__xor2_2 _16434_ (.A(_09031_),
    .B(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__buf_2 _16435_ (.A(_08678_),
    .X(_09046_));
 sky130_fd_sc_hd__and2_1 _16436_ (.A(_07661_),
    .B(_07662_),
    .X(_09047_));
 sky130_fd_sc_hd__or3_2 _16437_ (.A(_07617_),
    .B(_07646_),
    .C(_08681_),
    .X(_09048_));
 sky130_fd_sc_hd__or3b_1 _16438_ (.A(_09047_),
    .B(_08803_),
    .C_N(_09048_),
    .X(_09049_));
 sky130_fd_sc_hd__or2_1 _16439_ (.A(_07877_),
    .B(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__o21ai_1 _16440_ (.A1(_07877_),
    .A2(_09046_),
    .B1(_09049_),
    .Y(_09051_));
 sky130_fd_sc_hd__o21a_1 _16441_ (.A1(_09046_),
    .A2(_09050_),
    .B1(_09051_),
    .X(_09052_));
 sky130_fd_sc_hd__xnor2_1 _16442_ (.A(_08807_),
    .B(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__a21boi_1 _16443_ (.A1(_08807_),
    .A2(_08926_),
    .B1_N(_08805_),
    .Y(_09054_));
 sky130_fd_sc_hd__nor2_1 _16444_ (.A(_09053_),
    .B(_09054_),
    .Y(_09055_));
 sky130_fd_sc_hd__and2_1 _16445_ (.A(_09053_),
    .B(_09054_),
    .X(_09056_));
 sky130_fd_sc_hd__nor2_1 _16446_ (.A(_09055_),
    .B(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__xnor2_2 _16447_ (.A(_09045_),
    .B(_09057_),
    .Y(_09058_));
 sky130_fd_sc_hd__a21o_1 _16448_ (.A1(_08922_),
    .A2(_08931_),
    .B1(_08929_),
    .X(_09059_));
 sky130_fd_sc_hd__xnor2_1 _16449_ (.A(_09058_),
    .B(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__xnor2_1 _16450_ (.A(_09030_),
    .B(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__a21oi_1 _16451_ (.A1(_08908_),
    .A2(_08937_),
    .B1(_08935_),
    .Y(_09062_));
 sky130_fd_sc_hd__nor2_1 _16452_ (.A(_09061_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_1 _16453_ (.A(_09061_),
    .B(_09062_),
    .Y(_09064_));
 sky130_fd_sc_hd__and2b_1 _16454_ (.A_N(_09063_),
    .B(_09064_),
    .X(_09065_));
 sky130_fd_sc_hd__xnor2_1 _16455_ (.A(_09005_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__a21oi_1 _16456_ (.A1(_08882_),
    .A2(_08942_),
    .B1(_08940_),
    .Y(_09067_));
 sky130_fd_sc_hd__nor2_1 _16457_ (.A(_09066_),
    .B(_09067_),
    .Y(_09068_));
 sky130_fd_sc_hd__and2_1 _16458_ (.A(_09066_),
    .B(_09067_),
    .X(_09069_));
 sky130_fd_sc_hd__nor2_1 _16459_ (.A(_09068_),
    .B(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__xnor2_2 _16460_ (.A(_08972_),
    .B(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__nor2_1 _16461_ (.A(_08943_),
    .B(_08945_),
    .Y(_09072_));
 sky130_fd_sc_hd__a21oi_2 _16462_ (.A1(_08846_),
    .A2(_08946_),
    .B1(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__xor2_2 _16463_ (.A(_09071_),
    .B(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__xnor2_2 _16464_ (.A(_08844_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__xor2_2 _16465_ (.A(_08967_),
    .B(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__nand2_1 _16466_ (.A(_08952_),
    .B(_08953_),
    .Y(_09077_));
 sky130_fd_sc_hd__nor2_1 _16467_ (.A(_08952_),
    .B(_08953_),
    .Y(_09078_));
 sky130_fd_sc_hd__a21oi_2 _16468_ (.A1(_09077_),
    .A2(_08957_),
    .B1(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__o21ai_1 _16469_ (.A1(_09076_),
    .A2(_09079_),
    .B1(_08485_),
    .Y(_09080_));
 sky130_fd_sc_hd__a21oi_4 _16470_ (.A1(_09076_),
    .A2(_09079_),
    .B1(_09080_),
    .Y(_09081_));
 sky130_fd_sc_hd__nand2_1 _16471_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_09082_));
 sky130_fd_sc_hd__or2_1 _16472_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_09083_));
 sky130_fd_sc_hd__nand2_1 _16473_ (.A(_08960_),
    .B(_08965_),
    .Y(_09084_));
 sky130_fd_sc_hd__and3_1 _16474_ (.A(_09082_),
    .B(_09083_),
    .C(_09084_),
    .X(_09085_));
 sky130_fd_sc_hd__inv_2 _16475_ (.A(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__a21o_1 _16476_ (.A1(_09082_),
    .A2(_09083_),
    .B1(_09084_),
    .X(_09087_));
 sky130_fd_sc_hd__a31o_1 _16477_ (.A1(_08562_),
    .A2(_09086_),
    .A3(_09087_),
    .B1(_08487_),
    .X(_09088_));
 sky130_fd_sc_hd__o22a_1 _16478_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_08553_),
    .B1(_09081_),
    .B2(_09088_),
    .X(_00552_));
 sky130_fd_sc_hd__or2b_1 _16479_ (.A(_08967_),
    .B_N(_09075_),
    .X(_09089_));
 sky130_fd_sc_hd__nor2_1 _16480_ (.A(_08954_),
    .B(_09076_),
    .Y(_09090_));
 sky130_fd_sc_hd__and2b_1 _16481_ (.A_N(_09075_),
    .B(_08967_),
    .X(_09091_));
 sky130_fd_sc_hd__a221o_1 _16482_ (.A1(_09078_),
    .A2(_09089_),
    .B1(_09090_),
    .B2(_08957_),
    .C1(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__or2b_1 _16483_ (.A(_09004_),
    .B_N(_08973_),
    .X(_09093_));
 sky130_fd_sc_hd__a21oi_1 _16484_ (.A1(_08983_),
    .A2(_08984_),
    .B1(_08981_),
    .Y(_09094_));
 sky130_fd_sc_hd__a21oi_2 _16485_ (.A1(_09002_),
    .A2(_09093_),
    .B1(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__and3_1 _16486_ (.A(_09002_),
    .B(_09093_),
    .C(_09094_),
    .X(_09096_));
 sky130_fd_sc_hd__nor2_1 _16487_ (.A(_09095_),
    .B(_09096_),
    .Y(_09097_));
 sky130_fd_sc_hd__a21o_1 _16488_ (.A1(_08985_),
    .A2(_09000_),
    .B1(_08998_),
    .X(_09098_));
 sky130_fd_sc_hd__or2b_1 _16489_ (.A(_09029_),
    .B_N(_09006_),
    .X(_09099_));
 sky130_fd_sc_hd__nor2_1 _16490_ (.A(_07984_),
    .B(_08191_),
    .Y(_09100_));
 sky130_fd_sc_hd__or4_1 _16491_ (.A(_08643_),
    .B(_08107_),
    .C(_07960_),
    .D(_08070_),
    .X(_09101_));
 sky130_fd_sc_hd__inv_2 _16492_ (.A(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__o22a_1 _16493_ (.A1(_08643_),
    .A2(_07960_),
    .B1(_08071_),
    .B2(_08107_),
    .X(_09103_));
 sky130_fd_sc_hd__nor2_1 _16494_ (.A(_09102_),
    .B(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__xnor2_1 _16495_ (.A(_09100_),
    .B(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__o31a_1 _16496_ (.A1(_07865_),
    .A2(_08333_),
    .A3(_08978_),
    .B1(_08976_),
    .X(_09106_));
 sky130_fd_sc_hd__xnor2_1 _16497_ (.A(_09105_),
    .B(_09106_),
    .Y(_09107_));
 sky130_fd_sc_hd__and2_1 _16498_ (.A(_07865_),
    .B(_08317_),
    .X(_09108_));
 sky130_fd_sc_hd__xnor2_1 _16499_ (.A(_09107_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__clkbuf_4 _16500_ (.A(_08081_),
    .X(_09110_));
 sky130_fd_sc_hd__o31ai_1 _16501_ (.A1(_08643_),
    .A2(_09110_),
    .A3(_08989_),
    .B1(_08988_),
    .Y(_09111_));
 sky130_fd_sc_hd__a22o_1 _16502_ (.A1(_08885_),
    .A2(_09008_),
    .B1(_09010_),
    .B2(_09012_),
    .X(_09112_));
 sky130_fd_sc_hd__or3_1 _16503_ (.A(_07878_),
    .B(_07787_),
    .C(_08987_),
    .X(_09113_));
 sky130_fd_sc_hd__a2bb2o_1 _16504_ (.A1_N(_07878_),
    .A2_N(_07333_),
    .B1(_07784_),
    .B2(_08767_),
    .X(_09114_));
 sky130_fd_sc_hd__and2_1 _16505_ (.A(_09113_),
    .B(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__nor2_1 _16506_ (.A(_07993_),
    .B(_08081_),
    .Y(_09116_));
 sky130_fd_sc_hd__xor2_1 _16507_ (.A(_09115_),
    .B(_09116_),
    .X(_09117_));
 sky130_fd_sc_hd__and2_1 _16508_ (.A(_09112_),
    .B(_09117_),
    .X(_09118_));
 sky130_fd_sc_hd__nor2_1 _16509_ (.A(_09112_),
    .B(_09117_),
    .Y(_09119_));
 sky130_fd_sc_hd__nor2_1 _16510_ (.A(_09118_),
    .B(_09119_),
    .Y(_09120_));
 sky130_fd_sc_hd__xnor2_1 _16511_ (.A(_09111_),
    .B(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__a21oi_1 _16512_ (.A1(_08986_),
    .A2(_08995_),
    .B1(_08993_),
    .Y(_09122_));
 sky130_fd_sc_hd__nor2_1 _16513_ (.A(_09121_),
    .B(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__and2_1 _16514_ (.A(_09121_),
    .B(_09122_),
    .X(_09124_));
 sky130_fd_sc_hd__nor2_1 _16515_ (.A(_09123_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__xnor2_1 _16516_ (.A(_09109_),
    .B(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__a21o_1 _16517_ (.A1(_09027_),
    .A2(_09099_),
    .B1(_09126_),
    .X(_09127_));
 sky130_fd_sc_hd__nand3_1 _16518_ (.A(_09027_),
    .B(_09099_),
    .C(_09126_),
    .Y(_09128_));
 sky130_fd_sc_hd__nand2_1 _16519_ (.A(_09127_),
    .B(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__xnor2_1 _16520_ (.A(_09098_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__a21o_1 _16521_ (.A1(_09013_),
    .A2(_09025_),
    .B1(_09023_),
    .X(_09131_));
 sky130_fd_sc_hd__nand2_1 _16522_ (.A(_09031_),
    .B(_09044_),
    .Y(_09132_));
 sky130_fd_sc_hd__buf_2 _16523_ (.A(_08130_),
    .X(_09133_));
 sky130_fd_sc_hd__or4_1 _16524_ (.A(_06858_),
    .B(_07012_),
    .C(_07766_),
    .D(_09133_),
    .X(_09134_));
 sky130_fd_sc_hd__o21bai_1 _16525_ (.A1(_09009_),
    .A2(_09133_),
    .B1_N(_09008_),
    .Y(_09135_));
 sky130_fd_sc_hd__nand2_1 _16526_ (.A(_09134_),
    .B(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__nor2_1 _16527_ (.A(_08899_),
    .B(_07857_),
    .Y(_09137_));
 sky130_fd_sc_hd__xnor2_1 _16528_ (.A(_09136_),
    .B(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__or4_1 _16529_ (.A(_09014_),
    .B(_09016_),
    .C(_08134_),
    .D(_08260_),
    .X(_09139_));
 sky130_fd_sc_hd__o22ai_1 _16530_ (.A1(_09016_),
    .A2(_08134_),
    .B1(_09039_),
    .B2(_09014_),
    .Y(_09140_));
 sky130_fd_sc_hd__nand2_1 _16531_ (.A(_09139_),
    .B(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__buf_2 _16532_ (.A(_08133_),
    .X(_09142_));
 sky130_fd_sc_hd__nor2_1 _16533_ (.A(_08108_),
    .B(_09142_),
    .Y(_09143_));
 sky130_fd_sc_hd__xor2_1 _16534_ (.A(_09141_),
    .B(_09143_),
    .X(_09144_));
 sky130_fd_sc_hd__o31a_1 _16535_ (.A1(_09021_),
    .A2(_09133_),
    .A3(_09018_),
    .B1(_09015_),
    .X(_09145_));
 sky130_fd_sc_hd__nor2_1 _16536_ (.A(_09144_),
    .B(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__nand2_1 _16537_ (.A(_09144_),
    .B(_09145_),
    .Y(_09147_));
 sky130_fd_sc_hd__and2b_1 _16538_ (.A_N(_09146_),
    .B(_09147_),
    .X(_09148_));
 sky130_fd_sc_hd__xnor2_1 _16539_ (.A(_09138_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__a21o_1 _16540_ (.A1(_09042_),
    .A2(_09132_),
    .B1(_09149_),
    .X(_09150_));
 sky130_fd_sc_hd__nand3_1 _16541_ (.A(_09042_),
    .B(_09132_),
    .C(_09149_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_1 _16542_ (.A(_09150_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__xnor2_2 _16543_ (.A(_09131_),
    .B(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__a21bo_1 _16544_ (.A1(_09037_),
    .A2(_09040_),
    .B1_N(_09034_),
    .X(_09154_));
 sky130_fd_sc_hd__or2_1 _16545_ (.A(_09046_),
    .B(_09050_),
    .X(_09155_));
 sky130_fd_sc_hd__nor4_1 _16546_ (.A(_08247_),
    .B(_08245_),
    .C(_09036_),
    .D(_08678_),
    .Y(_09156_));
 sky130_fd_sc_hd__o22a_1 _16547_ (.A1(_08245_),
    .A2(_08391_),
    .B1(_08678_),
    .B2(_08247_),
    .X(_09157_));
 sky130_fd_sc_hd__nor2_1 _16548_ (.A(_09156_),
    .B(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__nor2_1 _16549_ (.A(_07992_),
    .B(_09035_),
    .Y(_09159_));
 sky130_fd_sc_hd__xnor2_1 _16550_ (.A(_09158_),
    .B(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__a21o_1 _16551_ (.A1(_09048_),
    .A2(_09155_),
    .B1(_09160_),
    .X(_09161_));
 sky130_fd_sc_hd__nand3_1 _16552_ (.A(_09048_),
    .B(_09155_),
    .C(_09160_),
    .Y(_09162_));
 sky130_fd_sc_hd__and2_1 _16553_ (.A(_09161_),
    .B(_09162_),
    .X(_09163_));
 sky130_fd_sc_hd__xor2_2 _16554_ (.A(_09154_),
    .B(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__nand2_1 _16555_ (.A(_08807_),
    .B(_09052_),
    .Y(_09165_));
 sky130_fd_sc_hd__o21ai_1 _16556_ (.A1(_07877_),
    .A2(_08803_),
    .B1(_09049_),
    .Y(_09166_));
 sky130_fd_sc_hd__and2_1 _16557_ (.A(_09050_),
    .B(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__xnor2_1 _16558_ (.A(_08807_),
    .B(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__a21oi_1 _16559_ (.A1(_08805_),
    .A2(_09165_),
    .B1(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__and3_1 _16560_ (.A(_08805_),
    .B(_09165_),
    .C(_09168_),
    .X(_09170_));
 sky130_fd_sc_hd__nor2_1 _16561_ (.A(_09169_),
    .B(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__xnor2_2 _16562_ (.A(_09164_),
    .B(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__a21oi_2 _16563_ (.A1(_09045_),
    .A2(_09057_),
    .B1(_09055_),
    .Y(_09173_));
 sky130_fd_sc_hd__xor2_2 _16564_ (.A(_09172_),
    .B(_09173_),
    .X(_09174_));
 sky130_fd_sc_hd__xnor2_2 _16565_ (.A(_09153_),
    .B(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__and2b_1 _16566_ (.A_N(_09058_),
    .B(_09059_),
    .X(_09176_));
 sky130_fd_sc_hd__a21oi_1 _16567_ (.A1(_09030_),
    .A2(_09060_),
    .B1(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__nor2_1 _16568_ (.A(_09175_),
    .B(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__and2_1 _16569_ (.A(_09175_),
    .B(_09177_),
    .X(_09179_));
 sky130_fd_sc_hd__nor2_1 _16570_ (.A(_09178_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__xnor2_1 _16571_ (.A(_09130_),
    .B(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__a21oi_1 _16572_ (.A1(_09005_),
    .A2(_09064_),
    .B1(_09063_),
    .Y(_09182_));
 sky130_fd_sc_hd__nor2_1 _16573_ (.A(_09181_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_1 _16574_ (.A(_09181_),
    .B(_09182_),
    .Y(_09184_));
 sky130_fd_sc_hd__and2b_1 _16575_ (.A_N(_09183_),
    .B(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__xnor2_1 _16576_ (.A(_09097_),
    .B(_09185_),
    .Y(_09186_));
 sky130_fd_sc_hd__a21oi_1 _16577_ (.A1(_08972_),
    .A2(_09070_),
    .B1(_09068_),
    .Y(_09187_));
 sky130_fd_sc_hd__xor2_1 _16578_ (.A(_09186_),
    .B(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__nand2_1 _16579_ (.A(_08970_),
    .B(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__or2_1 _16580_ (.A(_08970_),
    .B(_09188_),
    .X(_09190_));
 sky130_fd_sc_hd__nand2_1 _16581_ (.A(_09189_),
    .B(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__nor2_1 _16582_ (.A(_09071_),
    .B(_09073_),
    .Y(_09192_));
 sky130_fd_sc_hd__a21oi_1 _16583_ (.A1(_08844_),
    .A2(_09074_),
    .B1(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__xnor2_1 _16584_ (.A(_09191_),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__or2b_1 _16585_ (.A(_09092_),
    .B_N(_09194_),
    .X(_09195_));
 sky130_fd_sc_hd__or2b_1 _16586_ (.A(_09194_),
    .B_N(_09092_),
    .X(_09196_));
 sky130_fd_sc_hd__and3_2 _16587_ (.A(_08485_),
    .B(_09195_),
    .C(_09196_),
    .X(_09197_));
 sky130_fd_sc_hd__nand2_1 _16588_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_09198_));
 sky130_fd_sc_hd__or2_1 _16589_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_09199_));
 sky130_fd_sc_hd__nand2_1 _16590_ (.A(_09198_),
    .B(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__nand2_1 _16591_ (.A(_09082_),
    .B(_09086_),
    .Y(_09201_));
 sky130_fd_sc_hd__xnor2_1 _16592_ (.A(_09200_),
    .B(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__a21o_1 _16593_ (.A1(_08512_),
    .A2(_09202_),
    .B1(_08489_),
    .X(_09203_));
 sky130_fd_sc_hd__o22a_1 _16594_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(_08553_),
    .B1(_09197_),
    .B2(_09203_),
    .X(_00553_));
 sky130_fd_sc_hd__or2_1 _16595_ (.A(_09186_),
    .B(_09187_),
    .X(_09204_));
 sky130_fd_sc_hd__or2b_1 _16596_ (.A(_09129_),
    .B_N(_09098_),
    .X(_09205_));
 sky130_fd_sc_hd__or2b_1 _16597_ (.A(_09107_),
    .B_N(_09108_),
    .X(_09206_));
 sky130_fd_sc_hd__o21a_1 _16598_ (.A1(_09105_),
    .A2(_09106_),
    .B1(_09206_),
    .X(_09207_));
 sky130_fd_sc_hd__a21oi_1 _16599_ (.A1(_09127_),
    .A2(_09205_),
    .B1(_09207_),
    .Y(_09208_));
 sky130_fd_sc_hd__and3_1 _16600_ (.A(_09127_),
    .B(_09205_),
    .C(_09207_),
    .X(_09209_));
 sky130_fd_sc_hd__nor2_1 _16601_ (.A(_09208_),
    .B(_09209_),
    .Y(_09210_));
 sky130_fd_sc_hd__a21o_1 _16602_ (.A1(_09109_),
    .A2(_09125_),
    .B1(_09123_),
    .X(_09211_));
 sky130_fd_sc_hd__or2b_1 _16603_ (.A(_09152_),
    .B_N(_09131_),
    .X(_09212_));
 sky130_fd_sc_hd__nand2_2 _16604_ (.A(_09150_),
    .B(_09212_),
    .Y(_09213_));
 sky130_fd_sc_hd__nor2_1 _16605_ (.A(_08107_),
    .B(_08191_),
    .Y(_09214_));
 sky130_fd_sc_hd__nor2_1 _16606_ (.A(_07123_),
    .B(_08070_),
    .Y(_09215_));
 sky130_fd_sc_hd__or3b_1 _16607_ (.A(_08643_),
    .B(_07960_),
    .C_N(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__inv_2 _16608_ (.A(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__o22a_1 _16609_ (.A1(_07993_),
    .A2(_07960_),
    .B1(_08071_),
    .B2(_08643_),
    .X(_09218_));
 sky130_fd_sc_hd__nor2_1 _16610_ (.A(_09217_),
    .B(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__xnor2_1 _16611_ (.A(_09214_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__a21oi_1 _16612_ (.A1(_09100_),
    .A2(_09104_),
    .B1(_09102_),
    .Y(_09221_));
 sky130_fd_sc_hd__xnor2_1 _16613_ (.A(_09220_),
    .B(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand2_1 _16614_ (.A(_07984_),
    .B(_08316_),
    .Y(_09223_));
 sky130_fd_sc_hd__nor2_1 _16615_ (.A(_09222_),
    .B(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__and2_1 _16616_ (.A(_09222_),
    .B(_09223_),
    .X(_09225_));
 sky130_fd_sc_hd__or2_1 _16617_ (.A(_09224_),
    .B(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__a21bo_1 _16618_ (.A1(_09114_),
    .A2(_09116_),
    .B1_N(_09113_),
    .X(_09227_));
 sky130_fd_sc_hd__a21bo_1 _16619_ (.A1(_09135_),
    .A2(_09137_),
    .B1_N(_09134_),
    .X(_09228_));
 sky130_fd_sc_hd__buf_2 _16620_ (.A(_07787_),
    .X(_09229_));
 sky130_fd_sc_hd__nor2_1 _16621_ (.A(_08862_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__buf_2 _16622_ (.A(_07333_),
    .X(_09231_));
 sky130_fd_sc_hd__nor2_1 _16623_ (.A(_08252_),
    .B(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__or4_1 _16624_ (.A(_07878_),
    .B(_08252_),
    .C(_09231_),
    .D(_09229_),
    .X(_09233_));
 sky130_fd_sc_hd__o21ai_1 _16625_ (.A1(_09230_),
    .A2(_09232_),
    .B1(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__nor2_1 _16626_ (.A(_08888_),
    .B(_09110_),
    .Y(_09235_));
 sky130_fd_sc_hd__xnor2_1 _16627_ (.A(_09234_),
    .B(_09235_),
    .Y(_09236_));
 sky130_fd_sc_hd__and2_1 _16628_ (.A(_09228_),
    .B(_09236_),
    .X(_09237_));
 sky130_fd_sc_hd__nor2_1 _16629_ (.A(_09228_),
    .B(_09236_),
    .Y(_09238_));
 sky130_fd_sc_hd__nor2_1 _16630_ (.A(_09237_),
    .B(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__xnor2_1 _16631_ (.A(_09227_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__a21oi_1 _16632_ (.A1(_09111_),
    .A2(_09120_),
    .B1(_09118_),
    .Y(_09241_));
 sky130_fd_sc_hd__xor2_1 _16633_ (.A(_09240_),
    .B(_09241_),
    .X(_09242_));
 sky130_fd_sc_hd__xnor2_1 _16634_ (.A(_09226_),
    .B(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__xnor2_1 _16635_ (.A(_09213_),
    .B(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__xnor2_1 _16636_ (.A(_09211_),
    .B(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__a21o_1 _16637_ (.A1(_09138_),
    .A2(_09147_),
    .B1(_09146_),
    .X(_09246_));
 sky130_fd_sc_hd__nand2_1 _16638_ (.A(_09154_),
    .B(_09163_),
    .Y(_09247_));
 sky130_fd_sc_hd__or4_1 _16639_ (.A(_06858_),
    .B(_07012_),
    .C(_08130_),
    .D(_09142_),
    .X(_09248_));
 sky130_fd_sc_hd__a2bb2o_1 _16640_ (.A1_N(_07012_),
    .A2_N(_08130_),
    .B1(_07173_),
    .B2(_08766_),
    .X(_09249_));
 sky130_fd_sc_hd__nand2_1 _16641_ (.A(_09248_),
    .B(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__nor2_1 _16642_ (.A(_08896_),
    .B(_08889_),
    .Y(_09251_));
 sky130_fd_sc_hd__xnor2_1 _16643_ (.A(_09250_),
    .B(_09251_),
    .Y(_09252_));
 sky130_fd_sc_hd__or4_1 _16644_ (.A(_07494_),
    .B(_08229_),
    .C(_08260_),
    .D(_08018_),
    .X(_09253_));
 sky130_fd_sc_hd__o22ai_1 _16645_ (.A1(_09016_),
    .A2(_08260_),
    .B1(_09035_),
    .B2(_09014_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand2_1 _16646_ (.A(_09253_),
    .B(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__buf_2 _16647_ (.A(_08134_),
    .X(_09256_));
 sky130_fd_sc_hd__nor2_1 _16648_ (.A(_08108_),
    .B(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__xnor2_1 _16649_ (.A(_09255_),
    .B(_09257_),
    .Y(_09258_));
 sky130_fd_sc_hd__a21bo_1 _16650_ (.A1(_09140_),
    .A2(_09143_),
    .B1_N(_09139_),
    .X(_09259_));
 sky130_fd_sc_hd__xor2_1 _16651_ (.A(_09258_),
    .B(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__and2_1 _16652_ (.A(_09252_),
    .B(_09260_),
    .X(_09261_));
 sky130_fd_sc_hd__nor2_1 _16653_ (.A(_09252_),
    .B(_09260_),
    .Y(_09262_));
 sky130_fd_sc_hd__or2_1 _16654_ (.A(_09261_),
    .B(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__a21o_1 _16655_ (.A1(_09161_),
    .A2(_09247_),
    .B1(_09263_),
    .X(_09264_));
 sky130_fd_sc_hd__nand3_1 _16656_ (.A(_09161_),
    .B(_09247_),
    .C(_09263_),
    .Y(_09265_));
 sky130_fd_sc_hd__nand2_1 _16657_ (.A(_09264_),
    .B(_09265_),
    .Y(_09266_));
 sky130_fd_sc_hd__xnor2_2 _16658_ (.A(_09246_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__a21o_1 _16659_ (.A1(_09158_),
    .A2(_09159_),
    .B1(_09156_),
    .X(_09268_));
 sky130_fd_sc_hd__nand2_2 _16660_ (.A(_09048_),
    .B(_09050_),
    .Y(_09269_));
 sky130_fd_sc_hd__nor2_1 _16661_ (.A(_08245_),
    .B(_08678_),
    .Y(_09270_));
 sky130_fd_sc_hd__nor2_1 _16662_ (.A(_08247_),
    .B(_08681_),
    .Y(_09271_));
 sky130_fd_sc_hd__xnor2_1 _16663_ (.A(_09270_),
    .B(_09271_),
    .Y(_09272_));
 sky130_fd_sc_hd__or3_1 _16664_ (.A(_07992_),
    .B(_08391_),
    .C(_09272_),
    .X(_09273_));
 sky130_fd_sc_hd__o21ai_1 _16665_ (.A1(_07992_),
    .A2(_09036_),
    .B1(_09272_),
    .Y(_09274_));
 sky130_fd_sc_hd__and2_1 _16666_ (.A(_09273_),
    .B(_09274_),
    .X(_09275_));
 sky130_fd_sc_hd__xor2_1 _16667_ (.A(_09269_),
    .B(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__nand2_1 _16668_ (.A(_09268_),
    .B(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__or2_1 _16669_ (.A(_09268_),
    .B(_09276_),
    .X(_09278_));
 sky130_fd_sc_hd__and2_1 _16670_ (.A(_09277_),
    .B(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__or2b_2 _16671_ (.A(_08805_),
    .B_N(_09167_),
    .X(_09280_));
 sky130_fd_sc_hd__or2b_1 _16672_ (.A(_09167_),
    .B_N(_08804_),
    .X(_09281_));
 sky130_fd_sc_hd__and2_1 _16673_ (.A(_09280_),
    .B(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__buf_2 _16674_ (.A(_09282_),
    .X(_09283_));
 sky130_fd_sc_hd__xnor2_1 _16675_ (.A(_09279_),
    .B(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__a21oi_2 _16676_ (.A1(_09164_),
    .A2(_09171_),
    .B1(_09169_),
    .Y(_09285_));
 sky130_fd_sc_hd__nor2_1 _16677_ (.A(_09284_),
    .B(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__and2_1 _16678_ (.A(_09284_),
    .B(_09285_),
    .X(_09287_));
 sky130_fd_sc_hd__nor2_1 _16679_ (.A(_09286_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__xnor2_2 _16680_ (.A(_09267_),
    .B(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nor2_1 _16681_ (.A(_09172_),
    .B(_09173_),
    .Y(_09290_));
 sky130_fd_sc_hd__a21oi_2 _16682_ (.A1(_09153_),
    .A2(_09174_),
    .B1(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__xor2_1 _16683_ (.A(_09289_),
    .B(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__xnor2_1 _16684_ (.A(_09245_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__a21oi_1 _16685_ (.A1(_09130_),
    .A2(_09180_),
    .B1(_09178_),
    .Y(_09294_));
 sky130_fd_sc_hd__nor2_1 _16686_ (.A(_09293_),
    .B(_09294_),
    .Y(_09295_));
 sky130_fd_sc_hd__and2_1 _16687_ (.A(_09293_),
    .B(_09294_),
    .X(_09296_));
 sky130_fd_sc_hd__nor2_1 _16688_ (.A(_09295_),
    .B(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__xnor2_1 _16689_ (.A(_09210_),
    .B(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__a21oi_1 _16690_ (.A1(_09097_),
    .A2(_09184_),
    .B1(_09183_),
    .Y(_09299_));
 sky130_fd_sc_hd__xor2_1 _16691_ (.A(_09298_),
    .B(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__xnor2_1 _16692_ (.A(_09095_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__and3_1 _16693_ (.A(_09204_),
    .B(_09189_),
    .C(_09301_),
    .X(_09302_));
 sky130_fd_sc_hd__a21o_1 _16694_ (.A1(_09204_),
    .A2(_09189_),
    .B1(_09301_),
    .X(_09303_));
 sky130_fd_sc_hd__or2b_1 _16695_ (.A(_09302_),
    .B_N(_09303_),
    .X(_09304_));
 sky130_fd_sc_hd__or2_1 _16696_ (.A(_09191_),
    .B(_09193_),
    .X(_09305_));
 sky130_fd_sc_hd__and2_1 _16697_ (.A(_09305_),
    .B(_09196_),
    .X(_09306_));
 sky130_fd_sc_hd__o21ai_1 _16698_ (.A1(_09304_),
    .A2(_09306_),
    .B1(_08485_),
    .Y(_09307_));
 sky130_fd_sc_hd__a21oi_4 _16699_ (.A1(_09304_),
    .A2(_09306_),
    .B1(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__nor2_1 _16700_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_09309_));
 sky130_fd_sc_hd__and2_1 _16701_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_09310_));
 sky130_fd_sc_hd__a21boi_1 _16702_ (.A1(_09199_),
    .A2(_09201_),
    .B1_N(_09198_),
    .Y(_09311_));
 sky130_fd_sc_hd__or3_1 _16703_ (.A(_09309_),
    .B(_09310_),
    .C(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__o21ai_1 _16704_ (.A1(_09309_),
    .A2(_09310_),
    .B1(_09311_),
    .Y(_09313_));
 sky130_fd_sc_hd__a31o_1 _16705_ (.A1(_08562_),
    .A2(_09312_),
    .A3(_09313_),
    .B1(_08487_),
    .X(_09314_));
 sky130_fd_sc_hd__o22a_1 _16706_ (.A1(\rbzero.wall_tracer.trackDistX[5] ),
    .A2(_08553_),
    .B1(_09308_),
    .B2(_09314_),
    .X(_00554_));
 sky130_fd_sc_hd__nand2_1 _16707_ (.A(_09213_),
    .B(_09243_),
    .Y(_09315_));
 sky130_fd_sc_hd__or2b_1 _16708_ (.A(_09244_),
    .B_N(_09211_),
    .X(_09316_));
 sky130_fd_sc_hd__o21ba_1 _16709_ (.A1(_09220_),
    .A2(_09221_),
    .B1_N(_09224_),
    .X(_09317_));
 sky130_fd_sc_hd__a21oi_2 _16710_ (.A1(_09315_),
    .A2(_09316_),
    .B1(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__and3_1 _16711_ (.A(_09315_),
    .B(_09316_),
    .C(_09317_),
    .X(_09319_));
 sky130_fd_sc_hd__nor2_1 _16712_ (.A(_09318_),
    .B(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__or2b_1 _16713_ (.A(_09226_),
    .B_N(_09242_),
    .X(_09321_));
 sky130_fd_sc_hd__o21ai_1 _16714_ (.A1(_09240_),
    .A2(_09241_),
    .B1(_09321_),
    .Y(_09322_));
 sky130_fd_sc_hd__or2b_1 _16715_ (.A(_09266_),
    .B_N(_09246_),
    .X(_09323_));
 sky130_fd_sc_hd__nor2_1 _16716_ (.A(_08643_),
    .B(_08191_),
    .Y(_09324_));
 sky130_fd_sc_hd__nor2_1 _16717_ (.A(_08888_),
    .B(_07961_),
    .Y(_09325_));
 sky130_fd_sc_hd__or4_1 _16718_ (.A(_08000_),
    .B(_07993_),
    .C(_07960_),
    .D(_08070_),
    .X(_09326_));
 sky130_fd_sc_hd__o21a_1 _16719_ (.A1(_09215_),
    .A2(_09325_),
    .B1(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__xnor2_1 _16720_ (.A(_09324_),
    .B(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__a21oi_1 _16721_ (.A1(_09214_),
    .A2(_09219_),
    .B1(_09217_),
    .Y(_09329_));
 sky130_fd_sc_hd__nor2_1 _16722_ (.A(_09328_),
    .B(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__and2_1 _16723_ (.A(_09328_),
    .B(_09329_),
    .X(_09331_));
 sky130_fd_sc_hd__nor2_1 _16724_ (.A(_09330_),
    .B(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__and2_1 _16725_ (.A(_08107_),
    .B(_08317_),
    .X(_09333_));
 sky130_fd_sc_hd__xor2_1 _16726_ (.A(_09332_),
    .B(_09333_),
    .X(_09334_));
 sky130_fd_sc_hd__o31ai_2 _16727_ (.A1(_08888_),
    .A2(_09110_),
    .A3(_09234_),
    .B1(_09233_),
    .Y(_09335_));
 sky130_fd_sc_hd__o31a_1 _16728_ (.A1(_08896_),
    .A2(_08889_),
    .A3(_09250_),
    .B1(_09248_),
    .X(_09336_));
 sky130_fd_sc_hd__nor2_1 _16729_ (.A(_07766_),
    .B(_09229_),
    .Y(_09337_));
 sky130_fd_sc_hd__o22ai_1 _16730_ (.A1(_07766_),
    .A2(_09231_),
    .B1(_09229_),
    .B2(_08899_),
    .Y(_09338_));
 sky130_fd_sc_hd__a21bo_1 _16731_ (.A1(_09232_),
    .A2(_09337_),
    .B1_N(_09338_),
    .X(_09339_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_08862_),
    .B(_09110_),
    .Y(_09340_));
 sky130_fd_sc_hd__xnor2_1 _16733_ (.A(_09339_),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__and2b_1 _16734_ (.A_N(_09336_),
    .B(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__and2b_1 _16735_ (.A_N(_09341_),
    .B(_09336_),
    .X(_09343_));
 sky130_fd_sc_hd__nor2_1 _16736_ (.A(_09342_),
    .B(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__xnor2_1 _16737_ (.A(_09335_),
    .B(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__a21oi_1 _16738_ (.A1(_09227_),
    .A2(_09239_),
    .B1(_09237_),
    .Y(_09346_));
 sky130_fd_sc_hd__xor2_1 _16739_ (.A(_09345_),
    .B(_09346_),
    .X(_09347_));
 sky130_fd_sc_hd__nand2_1 _16740_ (.A(_09334_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__or2_1 _16741_ (.A(_09334_),
    .B(_09347_),
    .X(_09349_));
 sky130_fd_sc_hd__nand2_1 _16742_ (.A(_09348_),
    .B(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__a21o_1 _16743_ (.A1(_09264_),
    .A2(_09323_),
    .B1(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__nand3_1 _16744_ (.A(_09264_),
    .B(_09323_),
    .C(_09350_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_1 _16745_ (.A(_09351_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__xnor2_1 _16746_ (.A(_09322_),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__a21o_1 _16747_ (.A1(_09258_),
    .A2(_09259_),
    .B1(_09261_),
    .X(_09355_));
 sky130_fd_sc_hd__nand2_1 _16748_ (.A(_09269_),
    .B(_09275_),
    .Y(_09356_));
 sky130_fd_sc_hd__or4_1 _16749_ (.A(_09009_),
    .B(_09007_),
    .C(_09142_),
    .D(_08134_),
    .X(_09357_));
 sky130_fd_sc_hd__o22ai_1 _16750_ (.A1(_09007_),
    .A2(_09142_),
    .B1(_09256_),
    .B2(_09009_),
    .Y(_09358_));
 sky130_fd_sc_hd__nand2_1 _16751_ (.A(_09357_),
    .B(_09358_),
    .Y(_09359_));
 sky130_fd_sc_hd__nor2_1 _16752_ (.A(_09133_),
    .B(_08889_),
    .Y(_09360_));
 sky130_fd_sc_hd__xnor2_1 _16753_ (.A(_09359_),
    .B(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__or4_1 _16754_ (.A(_09014_),
    .B(_09016_),
    .C(_09035_),
    .D(_09036_),
    .X(_09362_));
 sky130_fd_sc_hd__o22ai_1 _16755_ (.A1(_09016_),
    .A2(_09035_),
    .B1(_09036_),
    .B2(_09014_),
    .Y(_09363_));
 sky130_fd_sc_hd__nand2_1 _16756_ (.A(_09362_),
    .B(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__nor2_1 _16757_ (.A(_09021_),
    .B(_09039_),
    .Y(_09365_));
 sky130_fd_sc_hd__xor2_1 _16758_ (.A(_09364_),
    .B(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__o31a_1 _16759_ (.A1(_09021_),
    .A2(_09256_),
    .A3(_09255_),
    .B1(_09253_),
    .X(_09367_));
 sky130_fd_sc_hd__nor2_1 _16760_ (.A(_09366_),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__and2_1 _16761_ (.A(_09366_),
    .B(_09367_),
    .X(_09369_));
 sky130_fd_sc_hd__nor2_1 _16762_ (.A(_09368_),
    .B(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__xnor2_1 _16763_ (.A(_09361_),
    .B(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__a21o_1 _16764_ (.A1(_09356_),
    .A2(_09277_),
    .B1(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__nand3_1 _16765_ (.A(_09356_),
    .B(_09277_),
    .C(_09371_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand2_1 _16766_ (.A(_09372_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__xnor2_1 _16767_ (.A(_09355_),
    .B(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__a21bo_1 _16768_ (.A1(_09270_),
    .A2(_09271_),
    .B1_N(_09273_),
    .X(_09376_));
 sky130_fd_sc_hd__or3_1 _16769_ (.A(_08247_),
    .B(_07530_),
    .C(_08681_),
    .X(_09377_));
 sky130_fd_sc_hd__a21oi_1 _16770_ (.A1(_08247_),
    .A2(_08245_),
    .B1(_08803_),
    .Y(_09378_));
 sky130_fd_sc_hd__and2_1 _16771_ (.A(_09377_),
    .B(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__nor2_1 _16772_ (.A(_07992_),
    .B(_09046_),
    .Y(_09380_));
 sky130_fd_sc_hd__or2b_1 _16773_ (.A(_07992_),
    .B_N(_09379_),
    .X(_09381_));
 sky130_fd_sc_hd__or2_1 _16774_ (.A(_09046_),
    .B(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__o21a_1 _16775_ (.A1(_09379_),
    .A2(_09380_),
    .B1(_09382_),
    .X(_09383_));
 sky130_fd_sc_hd__xnor2_1 _16776_ (.A(_09269_),
    .B(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__xnor2_1 _16777_ (.A(_09376_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__xnor2_1 _16778_ (.A(_09283_),
    .B(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__a21boi_1 _16779_ (.A1(_09279_),
    .A2(_09283_),
    .B1_N(_09280_),
    .Y(_09387_));
 sky130_fd_sc_hd__or2_1 _16780_ (.A(_09386_),
    .B(_09387_),
    .X(_09388_));
 sky130_fd_sc_hd__nand2_1 _16781_ (.A(_09386_),
    .B(_09387_),
    .Y(_09389_));
 sky130_fd_sc_hd__and2_1 _16782_ (.A(_09388_),
    .B(_09389_),
    .X(_09390_));
 sky130_fd_sc_hd__nand2_1 _16783_ (.A(_09375_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__or2_1 _16784_ (.A(_09375_),
    .B(_09390_),
    .X(_09392_));
 sky130_fd_sc_hd__nand2_1 _16785_ (.A(_09391_),
    .B(_09392_),
    .Y(_09393_));
 sky130_fd_sc_hd__a21oi_2 _16786_ (.A1(_09267_),
    .A2(_09288_),
    .B1(_09286_),
    .Y(_09394_));
 sky130_fd_sc_hd__xor2_2 _16787_ (.A(_09393_),
    .B(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__xnor2_2 _16788_ (.A(_09354_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__nor2_1 _16789_ (.A(_09289_),
    .B(_09291_),
    .Y(_09397_));
 sky130_fd_sc_hd__a21oi_1 _16790_ (.A1(_09245_),
    .A2(_09292_),
    .B1(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__xor2_1 _16791_ (.A(_09396_),
    .B(_09398_),
    .X(_09399_));
 sky130_fd_sc_hd__xnor2_1 _16792_ (.A(_09320_),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__a21o_1 _16793_ (.A1(_09210_),
    .A2(_09297_),
    .B1(_09295_),
    .X(_09401_));
 sky130_fd_sc_hd__xnor2_1 _16794_ (.A(_09400_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__nand2_1 _16795_ (.A(_09208_),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__or2_1 _16796_ (.A(_09208_),
    .B(_09402_),
    .X(_09404_));
 sky130_fd_sc_hd__nand2_1 _16797_ (.A(_09403_),
    .B(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__nor2_1 _16798_ (.A(_09298_),
    .B(_09299_),
    .Y(_09406_));
 sky130_fd_sc_hd__a21oi_1 _16799_ (.A1(_09095_),
    .A2(_09300_),
    .B1(_09406_),
    .Y(_09407_));
 sky130_fd_sc_hd__or2_1 _16800_ (.A(_09405_),
    .B(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__nand2_1 _16801_ (.A(_09405_),
    .B(_09407_),
    .Y(_09409_));
 sky130_fd_sc_hd__nand2_1 _16802_ (.A(_09408_),
    .B(_09409_),
    .Y(_09410_));
 sky130_fd_sc_hd__nor2_1 _16803_ (.A(_09194_),
    .B(_09304_),
    .Y(_09411_));
 sky130_fd_sc_hd__a21oi_1 _16804_ (.A1(_09305_),
    .A2(_09303_),
    .B1(_09302_),
    .Y(_09412_));
 sky130_fd_sc_hd__a21oi_1 _16805_ (.A1(_09092_),
    .A2(_09411_),
    .B1(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(_09410_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__or2_1 _16807_ (.A(_09410_),
    .B(_09413_),
    .X(_09415_));
 sky130_fd_sc_hd__and3_2 _16808_ (.A(_08485_),
    .B(_09414_),
    .C(_09415_),
    .X(_09416_));
 sky130_fd_sc_hd__nor2_1 _16809_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_09417_));
 sky130_fd_sc_hd__and2_1 _16810_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .X(_09418_));
 sky130_fd_sc_hd__o21ba_1 _16811_ (.A1(_09309_),
    .A2(_09311_),
    .B1_N(_09310_),
    .X(_09419_));
 sky130_fd_sc_hd__or3_1 _16812_ (.A(_09417_),
    .B(_09418_),
    .C(_09419_),
    .X(_09420_));
 sky130_fd_sc_hd__o21ai_1 _16813_ (.A1(_09417_),
    .A2(_09418_),
    .B1(_09419_),
    .Y(_09421_));
 sky130_fd_sc_hd__a31o_1 _16814_ (.A1(_08562_),
    .A2(_09420_),
    .A3(_09421_),
    .B1(_08487_),
    .X(_09422_));
 sky130_fd_sc_hd__o22a_1 _16815_ (.A1(\rbzero.wall_tracer.trackDistX[6] ),
    .A2(_08553_),
    .B1(_09416_),
    .B2(_09422_),
    .X(_00555_));
 sky130_fd_sc_hd__or2b_1 _16816_ (.A(_09400_),
    .B_N(_09401_),
    .X(_09423_));
 sky130_fd_sc_hd__or2b_1 _16817_ (.A(_09353_),
    .B_N(_09322_),
    .X(_09424_));
 sky130_fd_sc_hd__a21oi_1 _16818_ (.A1(_09332_),
    .A2(_09333_),
    .B1(_09330_),
    .Y(_09425_));
 sky130_fd_sc_hd__a21oi_1 _16819_ (.A1(_09351_),
    .A2(_09424_),
    .B1(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__and3_1 _16820_ (.A(_09351_),
    .B(_09424_),
    .C(_09425_),
    .X(_09427_));
 sky130_fd_sc_hd__nor2_1 _16821_ (.A(_09426_),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__nor2_1 _16822_ (.A(_09393_),
    .B(_09394_),
    .Y(_09429_));
 sky130_fd_sc_hd__and2_1 _16823_ (.A(_09354_),
    .B(_09395_),
    .X(_09430_));
 sky130_fd_sc_hd__or2b_1 _16824_ (.A(_09374_),
    .B_N(_09355_),
    .X(_09431_));
 sky130_fd_sc_hd__nand2_1 _16825_ (.A(_09372_),
    .B(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__nor2_1 _16826_ (.A(_08862_),
    .B(_08071_),
    .Y(_09433_));
 sky130_fd_sc_hd__o22a_1 _16827_ (.A1(_08862_),
    .A2(_07961_),
    .B1(_08071_),
    .B2(_08888_),
    .X(_09434_));
 sky130_fd_sc_hd__a21oi_1 _16828_ (.A1(_09325_),
    .A2(_09433_),
    .B1(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__nor2_1 _16829_ (.A(_07993_),
    .B(_08333_),
    .Y(_09436_));
 sky130_fd_sc_hd__xnor2_1 _16830_ (.A(_09435_),
    .B(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__a21boi_1 _16831_ (.A1(_09324_),
    .A2(_09327_),
    .B1_N(_09326_),
    .Y(_09438_));
 sky130_fd_sc_hd__xor2_1 _16832_ (.A(_09437_),
    .B(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__and2_1 _16833_ (.A(_08643_),
    .B(_08317_),
    .X(_09440_));
 sky130_fd_sc_hd__nand2_1 _16834_ (.A(_09439_),
    .B(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__or2_1 _16835_ (.A(_09439_),
    .B(_09440_),
    .X(_09442_));
 sky130_fd_sc_hd__and2_1 _16836_ (.A(_09441_),
    .B(_09442_),
    .X(_09443_));
 sky130_fd_sc_hd__a22o_1 _16837_ (.A1(_09232_),
    .A2(_09337_),
    .B1(_09338_),
    .B2(_09340_),
    .X(_09444_));
 sky130_fd_sc_hd__a21bo_1 _16838_ (.A1(_09358_),
    .A2(_09360_),
    .B1_N(_09357_),
    .X(_09445_));
 sky130_fd_sc_hd__or4_1 _16839_ (.A(_07766_),
    .B(_08130_),
    .C(_09231_),
    .D(_09229_),
    .X(_09446_));
 sky130_fd_sc_hd__o21bai_1 _16840_ (.A1(_09133_),
    .A2(_09231_),
    .B1_N(_09337_),
    .Y(_09447_));
 sky130_fd_sc_hd__nand2_1 _16841_ (.A(_09446_),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__nor2_1 _16842_ (.A(_08899_),
    .B(_09110_),
    .Y(_09449_));
 sky130_fd_sc_hd__xnor2_1 _16843_ (.A(_09448_),
    .B(_09449_),
    .Y(_09450_));
 sky130_fd_sc_hd__xor2_1 _16844_ (.A(_09445_),
    .B(_09450_),
    .X(_09451_));
 sky130_fd_sc_hd__and2_1 _16845_ (.A(_09444_),
    .B(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__nor2_1 _16846_ (.A(_09444_),
    .B(_09451_),
    .Y(_09453_));
 sky130_fd_sc_hd__or2_1 _16847_ (.A(_09452_),
    .B(_09453_),
    .X(_09454_));
 sky130_fd_sc_hd__a21oi_1 _16848_ (.A1(_09335_),
    .A2(_09344_),
    .B1(_09342_),
    .Y(_09455_));
 sky130_fd_sc_hd__nor2_1 _16849_ (.A(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__and2_1 _16850_ (.A(_09454_),
    .B(_09455_),
    .X(_09457_));
 sky130_fd_sc_hd__nor2_1 _16851_ (.A(_09456_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__xnor2_1 _16852_ (.A(_09443_),
    .B(_09458_),
    .Y(_09459_));
 sky130_fd_sc_hd__xor2_1 _16853_ (.A(_09432_),
    .B(_09459_),
    .X(_09460_));
 sky130_fd_sc_hd__o21ai_1 _16854_ (.A1(_09345_),
    .A2(_09346_),
    .B1(_09348_),
    .Y(_09461_));
 sky130_fd_sc_hd__or2b_1 _16855_ (.A(_09460_),
    .B_N(_09461_),
    .X(_09462_));
 sky130_fd_sc_hd__or2b_1 _16856_ (.A(_09461_),
    .B_N(_09460_),
    .X(_09463_));
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(_09462_),
    .B(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand2_1 _16858_ (.A(_09377_),
    .B(_09382_),
    .Y(_09465_));
 sky130_fd_sc_hd__nor2_1 _16859_ (.A(_07992_),
    .B(_08803_),
    .Y(_09466_));
 sky130_fd_sc_hd__o21a_1 _16860_ (.A1(_09379_),
    .A2(_09466_),
    .B1(_09381_),
    .X(_09467_));
 sky130_fd_sc_hd__nand2_1 _16861_ (.A(_09269_),
    .B(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__or2_1 _16862_ (.A(_09269_),
    .B(_09467_),
    .X(_09469_));
 sky130_fd_sc_hd__nand2_2 _16863_ (.A(_09468_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__xnor2_1 _16864_ (.A(_09465_),
    .B(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__xnor2_1 _16865_ (.A(_09283_),
    .B(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__a21boi_1 _16866_ (.A1(_09283_),
    .A2(_09385_),
    .B1_N(_09280_),
    .Y(_09473_));
 sky130_fd_sc_hd__nor2_1 _16867_ (.A(_09472_),
    .B(_09473_),
    .Y(_09474_));
 sky130_fd_sc_hd__and2_1 _16868_ (.A(_09472_),
    .B(_09473_),
    .X(_09475_));
 sky130_fd_sc_hd__nor2_1 _16869_ (.A(_09474_),
    .B(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__a21o_1 _16870_ (.A1(_09361_),
    .A2(_09370_),
    .B1(_09368_),
    .X(_09477_));
 sky130_fd_sc_hd__nand2_1 _16871_ (.A(_09269_),
    .B(_09383_),
    .Y(_09478_));
 sky130_fd_sc_hd__or2b_1 _16872_ (.A(_09384_),
    .B_N(_09376_),
    .X(_09479_));
 sky130_fd_sc_hd__nor4_1 _16873_ (.A(_09009_),
    .B(_09007_),
    .C(_09256_),
    .D(_09039_),
    .Y(_09480_));
 sky130_fd_sc_hd__o22a_1 _16874_ (.A1(_09007_),
    .A2(_09256_),
    .B1(_09039_),
    .B2(_09009_),
    .X(_09481_));
 sky130_fd_sc_hd__or2_1 _16875_ (.A(_09480_),
    .B(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__nor2_1 _16876_ (.A(_09142_),
    .B(_08889_),
    .Y(_09483_));
 sky130_fd_sc_hd__xnor2_1 _16877_ (.A(_09482_),
    .B(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__or2_1 _16878_ (.A(_09016_),
    .B(_08678_),
    .X(_09485_));
 sky130_fd_sc_hd__nor3_1 _16879_ (.A(_09014_),
    .B(_09036_),
    .C(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__o22a_1 _16880_ (.A1(_09016_),
    .A2(_09036_),
    .B1(_09046_),
    .B2(_09014_),
    .X(_09487_));
 sky130_fd_sc_hd__nor2_1 _16881_ (.A(_09486_),
    .B(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__nor2_1 _16882_ (.A(_09021_),
    .B(_09035_),
    .Y(_09489_));
 sky130_fd_sc_hd__xnor2_2 _16883_ (.A(_09488_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__o31a_1 _16884_ (.A1(_09021_),
    .A2(_09039_),
    .A3(_09364_),
    .B1(_09362_),
    .X(_09491_));
 sky130_fd_sc_hd__xor2_1 _16885_ (.A(_09490_),
    .B(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__nand2_1 _16886_ (.A(_09484_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__or2_1 _16887_ (.A(_09484_),
    .B(_09492_),
    .X(_09494_));
 sky130_fd_sc_hd__nand2_1 _16888_ (.A(_09493_),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__a21o_1 _16889_ (.A1(_09478_),
    .A2(_09479_),
    .B1(_09495_),
    .X(_09496_));
 sky130_fd_sc_hd__nand3_1 _16890_ (.A(_09478_),
    .B(_09479_),
    .C(_09495_),
    .Y(_09497_));
 sky130_fd_sc_hd__nand2_1 _16891_ (.A(_09496_),
    .B(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__xnor2_1 _16892_ (.A(_09477_),
    .B(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__xnor2_1 _16893_ (.A(_09476_),
    .B(_09499_),
    .Y(_09500_));
 sky130_fd_sc_hd__a21oi_1 _16894_ (.A1(_09388_),
    .A2(_09391_),
    .B1(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__and3_1 _16895_ (.A(_09388_),
    .B(_09391_),
    .C(_09500_),
    .X(_09502_));
 sky130_fd_sc_hd__nor2_1 _16896_ (.A(_09501_),
    .B(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__xnor2_1 _16897_ (.A(_09464_),
    .B(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__o21ai_1 _16898_ (.A1(_09429_),
    .A2(_09430_),
    .B1(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__or3_1 _16899_ (.A(_09429_),
    .B(_09430_),
    .C(_09504_),
    .X(_09506_));
 sky130_fd_sc_hd__nand2_1 _16900_ (.A(_09505_),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__xor2_2 _16901_ (.A(_09428_),
    .B(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__nor2_1 _16902_ (.A(_09396_),
    .B(_09398_),
    .Y(_09509_));
 sky130_fd_sc_hd__a21oi_1 _16903_ (.A1(_09320_),
    .A2(_09399_),
    .B1(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__nor2_1 _16904_ (.A(_09508_),
    .B(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__and2_1 _16905_ (.A(_09508_),
    .B(_09510_),
    .X(_09512_));
 sky130_fd_sc_hd__nor2_1 _16906_ (.A(_09511_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__xnor2_1 _16907_ (.A(_09318_),
    .B(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__a21oi_1 _16908_ (.A1(_09423_),
    .A2(_09403_),
    .B1(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand3_1 _16909_ (.A(_09423_),
    .B(_09403_),
    .C(_09514_),
    .Y(_09516_));
 sky130_fd_sc_hd__and2b_1 _16910_ (.A_N(_09515_),
    .B(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__nand2_1 _16911_ (.A(_09408_),
    .B(_09415_),
    .Y(_09518_));
 sky130_fd_sc_hd__a21oi_1 _16912_ (.A1(_09517_),
    .A2(_09518_),
    .B1(_08509_),
    .Y(_09519_));
 sky130_fd_sc_hd__o21ai_2 _16913_ (.A1(_09517_),
    .A2(_09518_),
    .B1(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__nor2_1 _16914_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_09521_));
 sky130_fd_sc_hd__nand2_1 _16915_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_09522_));
 sky130_fd_sc_hd__and2b_1 _16916_ (.A_N(_09521_),
    .B(_09522_),
    .X(_09523_));
 sky130_fd_sc_hd__o21ba_1 _16917_ (.A1(_09417_),
    .A2(_09419_),
    .B1_N(_09418_),
    .X(_09524_));
 sky130_fd_sc_hd__xnor2_1 _16918_ (.A(_09523_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__a21oi_1 _16919_ (.A1(_08512_),
    .A2(_09525_),
    .B1(_08489_),
    .Y(_09526_));
 sky130_fd_sc_hd__o2bb2a_1 _16920_ (.A1_N(_09520_),
    .A2_N(_09526_),
    .B1(\rbzero.wall_tracer.trackDistX[7] ),
    .B2(_08508_),
    .X(_00556_));
 sky130_fd_sc_hd__a21o_1 _16921_ (.A1(_09372_),
    .A2(_09431_),
    .B1(_09459_),
    .X(_09527_));
 sky130_fd_sc_hd__o21a_1 _16922_ (.A1(_09437_),
    .A2(_09438_),
    .B1(_09441_),
    .X(_09528_));
 sky130_fd_sc_hd__a21oi_2 _16923_ (.A1(_09527_),
    .A2(_09462_),
    .B1(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__and3_1 _16924_ (.A(_09527_),
    .B(_09462_),
    .C(_09528_),
    .X(_09530_));
 sky130_fd_sc_hd__nor2_1 _16925_ (.A(_09529_),
    .B(_09530_),
    .Y(_09531_));
 sky130_fd_sc_hd__a21bo_1 _16926_ (.A1(_09283_),
    .A2(_09471_),
    .B1_N(_09280_),
    .X(_09532_));
 sky130_fd_sc_hd__and2_1 _16927_ (.A(_09377_),
    .B(_09381_),
    .X(_09533_));
 sky130_fd_sc_hd__xor2_2 _16928_ (.A(_09470_),
    .B(_09533_),
    .X(_09534_));
 sky130_fd_sc_hd__xor2_1 _16929_ (.A(_09283_),
    .B(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__xnor2_1 _16930_ (.A(_09532_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__o21ai_2 _16931_ (.A1(_09490_),
    .A2(_09491_),
    .B1(_09493_),
    .Y(_09537_));
 sky130_fd_sc_hd__or2b_1 _16932_ (.A(_09470_),
    .B_N(_09465_),
    .X(_09538_));
 sky130_fd_sc_hd__nand2_1 _16933_ (.A(_09468_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__nor2_1 _16934_ (.A(_09007_),
    .B(_09039_),
    .Y(_09540_));
 sky130_fd_sc_hd__nor2_1 _16935_ (.A(_09009_),
    .B(_09035_),
    .Y(_09541_));
 sky130_fd_sc_hd__or4_1 _16936_ (.A(_09009_),
    .B(_09007_),
    .C(_09039_),
    .D(_09035_),
    .X(_09542_));
 sky130_fd_sc_hd__o21ai_2 _16937_ (.A1(_09540_),
    .A2(_09541_),
    .B1(_09542_),
    .Y(_09543_));
 sky130_fd_sc_hd__nor2_1 _16938_ (.A(_08889_),
    .B(_09256_),
    .Y(_09544_));
 sky130_fd_sc_hd__xnor2_2 _16939_ (.A(_09543_),
    .B(_09544_),
    .Y(_09545_));
 sky130_fd_sc_hd__or2_1 _16940_ (.A(_07494_),
    .B(_08803_),
    .X(_09546_));
 sky130_fd_sc_hd__or2_1 _16941_ (.A(_09016_),
    .B(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__nor2_1 _16942_ (.A(_09046_),
    .B(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__a21oi_1 _16943_ (.A1(_09485_),
    .A2(_09546_),
    .B1(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__nor2_1 _16944_ (.A(_09021_),
    .B(_09036_),
    .Y(_09550_));
 sky130_fd_sc_hd__and2_1 _16945_ (.A(_09549_),
    .B(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__nor2_1 _16946_ (.A(_09549_),
    .B(_09550_),
    .Y(_09552_));
 sky130_fd_sc_hd__or2_1 _16947_ (.A(_09551_),
    .B(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__a21oi_1 _16948_ (.A1(_09488_),
    .A2(_09489_),
    .B1(_09486_),
    .Y(_09554_));
 sky130_fd_sc_hd__nor2_1 _16949_ (.A(_09553_),
    .B(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__nand2_1 _16950_ (.A(_09553_),
    .B(_09554_),
    .Y(_09556_));
 sky130_fd_sc_hd__and2b_1 _16951_ (.A_N(_09555_),
    .B(_09556_),
    .X(_09557_));
 sky130_fd_sc_hd__xor2_1 _16952_ (.A(_09545_),
    .B(_09557_),
    .X(_09558_));
 sky130_fd_sc_hd__xnor2_1 _16953_ (.A(_09539_),
    .B(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__xnor2_2 _16954_ (.A(_09537_),
    .B(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__xor2_2 _16955_ (.A(_09536_),
    .B(_09560_),
    .X(_09561_));
 sky130_fd_sc_hd__a21oi_1 _16956_ (.A1(_09476_),
    .A2(_09499_),
    .B1(_09474_),
    .Y(_09562_));
 sky130_fd_sc_hd__xor2_1 _16957_ (.A(_09561_),
    .B(_09562_),
    .X(_09563_));
 sky130_fd_sc_hd__a21o_1 _16958_ (.A1(_09443_),
    .A2(_09458_),
    .B1(_09456_),
    .X(_09564_));
 sky130_fd_sc_hd__or2b_1 _16959_ (.A(_09498_),
    .B_N(_09477_),
    .X(_09565_));
 sky130_fd_sc_hd__nor2_1 _16960_ (.A(_08899_),
    .B(_07961_),
    .Y(_09566_));
 sky130_fd_sc_hd__or4_1 _16961_ (.A(_08862_),
    .B(_08899_),
    .C(_07961_),
    .D(_08071_),
    .X(_09567_));
 sky130_fd_sc_hd__o21ai_1 _16962_ (.A1(_09433_),
    .A2(_09566_),
    .B1(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__nor2_1 _16963_ (.A(_08888_),
    .B(_08333_),
    .Y(_09569_));
 sky130_fd_sc_hd__xor2_1 _16964_ (.A(_09568_),
    .B(_09569_),
    .X(_09570_));
 sky130_fd_sc_hd__nand2_1 _16965_ (.A(_09325_),
    .B(_09433_),
    .Y(_09571_));
 sky130_fd_sc_hd__o31a_1 _16966_ (.A1(_07993_),
    .A2(_08333_),
    .A3(_09434_),
    .B1(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__nor2_1 _16967_ (.A(_09570_),
    .B(_09572_),
    .Y(_09573_));
 sky130_fd_sc_hd__and2_1 _16968_ (.A(_09570_),
    .B(_09572_),
    .X(_09574_));
 sky130_fd_sc_hd__nor2_1 _16969_ (.A(_09573_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__and2_1 _16970_ (.A(_07993_),
    .B(_08317_),
    .X(_09576_));
 sky130_fd_sc_hd__xor2_1 _16971_ (.A(_09575_),
    .B(_09576_),
    .X(_09577_));
 sky130_fd_sc_hd__a21bo_1 _16972_ (.A1(_09447_),
    .A2(_09449_),
    .B1_N(_09446_),
    .X(_09578_));
 sky130_fd_sc_hd__inv_2 _16973_ (.A(_09481_),
    .Y(_09579_));
 sky130_fd_sc_hd__a21o_1 _16974_ (.A1(_09579_),
    .A2(_09483_),
    .B1(_09480_),
    .X(_09580_));
 sky130_fd_sc_hd__or4_1 _16975_ (.A(_09133_),
    .B(_09142_),
    .C(_09231_),
    .D(_09229_),
    .X(_09581_));
 sky130_fd_sc_hd__o22ai_1 _16976_ (.A1(_09142_),
    .A2(_09231_),
    .B1(_09229_),
    .B2(_09133_),
    .Y(_09582_));
 sky130_fd_sc_hd__nand2_1 _16977_ (.A(_09581_),
    .B(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__nor2_1 _16978_ (.A(_08896_),
    .B(_09110_),
    .Y(_09584_));
 sky130_fd_sc_hd__xnor2_1 _16979_ (.A(_09583_),
    .B(_09584_),
    .Y(_09585_));
 sky130_fd_sc_hd__and2_1 _16980_ (.A(_09580_),
    .B(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__nor2_1 _16981_ (.A(_09580_),
    .B(_09585_),
    .Y(_09587_));
 sky130_fd_sc_hd__nor2_1 _16982_ (.A(_09586_),
    .B(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__xnor2_1 _16983_ (.A(_09578_),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__a21oi_1 _16984_ (.A1(_09445_),
    .A2(_09450_),
    .B1(_09452_),
    .Y(_09590_));
 sky130_fd_sc_hd__xor2_1 _16985_ (.A(_09589_),
    .B(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__nand2_1 _16986_ (.A(_09577_),
    .B(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__or2_1 _16987_ (.A(_09577_),
    .B(_09591_),
    .X(_09593_));
 sky130_fd_sc_hd__nand2_1 _16988_ (.A(_09592_),
    .B(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__a21oi_1 _16989_ (.A1(_09496_),
    .A2(_09565_),
    .B1(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__and3_1 _16990_ (.A(_09496_),
    .B(_09565_),
    .C(_09594_),
    .X(_09596_));
 sky130_fd_sc_hd__or2_1 _16991_ (.A(_09595_),
    .B(_09596_),
    .X(_09597_));
 sky130_fd_sc_hd__xnor2_1 _16992_ (.A(_09564_),
    .B(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand2_1 _16993_ (.A(_09563_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__or2_1 _16994_ (.A(_09563_),
    .B(_09598_),
    .X(_09600_));
 sky130_fd_sc_hd__nand2_1 _16995_ (.A(_09599_),
    .B(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__o21ba_1 _16996_ (.A1(_09464_),
    .A2(_09502_),
    .B1_N(_09501_),
    .X(_09602_));
 sky130_fd_sc_hd__xor2_1 _16997_ (.A(_09601_),
    .B(_09602_),
    .X(_09603_));
 sky130_fd_sc_hd__nand2_1 _16998_ (.A(_09531_),
    .B(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__or2_1 _16999_ (.A(_09531_),
    .B(_09603_),
    .X(_09605_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_09604_),
    .B(_09605_),
    .Y(_09606_));
 sky130_fd_sc_hd__a21boi_1 _17001_ (.A1(_09428_),
    .A2(_09506_),
    .B1_N(_09505_),
    .Y(_09607_));
 sky130_fd_sc_hd__xor2_1 _17002_ (.A(_09606_),
    .B(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__nand2_1 _17003_ (.A(_09426_),
    .B(_09608_),
    .Y(_09609_));
 sky130_fd_sc_hd__or2_1 _17004_ (.A(_09426_),
    .B(_09608_),
    .X(_09610_));
 sky130_fd_sc_hd__nand2_1 _17005_ (.A(_09609_),
    .B(_09610_),
    .Y(_09611_));
 sky130_fd_sc_hd__a21oi_1 _17006_ (.A1(_09318_),
    .A2(_09513_),
    .B1(_09511_),
    .Y(_09612_));
 sky130_fd_sc_hd__nor2_1 _17007_ (.A(_09611_),
    .B(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__and2_1 _17008_ (.A(_09611_),
    .B(_09612_),
    .X(_09614_));
 sky130_fd_sc_hd__nor2_2 _17009_ (.A(_09613_),
    .B(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__a21o_1 _17010_ (.A1(_09092_),
    .A2(_09411_),
    .B1(_09412_),
    .X(_09616_));
 sky130_fd_sc_hd__inv_2 _17011_ (.A(_09408_),
    .Y(_09617_));
 sky130_fd_sc_hd__a21o_1 _17012_ (.A1(_09617_),
    .A2(_09516_),
    .B1(_09515_),
    .X(_09618_));
 sky130_fd_sc_hd__a41o_2 _17013_ (.A1(_09408_),
    .A2(_09409_),
    .A3(_09616_),
    .A4(_09517_),
    .B1(_09618_),
    .X(_09619_));
 sky130_fd_sc_hd__buf_6 _17014_ (.A(\rbzero.wall_tracer.state[1] ),
    .X(_09620_));
 sky130_fd_sc_hd__a21oi_1 _17015_ (.A1(_09615_),
    .A2(_09619_),
    .B1(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__o21ai_2 _17016_ (.A1(_09615_),
    .A2(_09619_),
    .B1(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__or2_1 _17017_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .X(_09623_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_09624_));
 sky130_fd_sc_hd__o21ai_1 _17019_ (.A1(_09521_),
    .A2(_09524_),
    .B1(_09522_),
    .Y(_09625_));
 sky130_fd_sc_hd__a21oi_1 _17020_ (.A1(_09623_),
    .A2(_09624_),
    .B1(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__a31o_1 _17021_ (.A1(_09623_),
    .A2(_09624_),
    .A3(_09625_),
    .B1(_04946_),
    .X(_09627_));
 sky130_fd_sc_hd__o21a_1 _17022_ (.A1(_09626_),
    .A2(_09627_),
    .B1(_08507_),
    .X(_09628_));
 sky130_fd_sc_hd__o2bb2a_1 _17023_ (.A1_N(_09622_),
    .A2_N(_09628_),
    .B1(\rbzero.wall_tracer.trackDistX[8] ),
    .B2(_08508_),
    .X(_00557_));
 sky130_fd_sc_hd__or2_1 _17024_ (.A(_09606_),
    .B(_09607_),
    .X(_09629_));
 sky130_fd_sc_hd__or2_1 _17025_ (.A(_09601_),
    .B(_09602_),
    .X(_09630_));
 sky130_fd_sc_hd__and2b_1 _17026_ (.A_N(_09536_),
    .B(_09560_),
    .X(_09631_));
 sky130_fd_sc_hd__a21o_1 _17027_ (.A1(_09532_),
    .A2(_09535_),
    .B1(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__nor2_1 _17028_ (.A(_09281_),
    .B(_09534_),
    .Y(_09633_));
 sky130_fd_sc_hd__inv_2 _17029_ (.A(_09534_),
    .Y(_09634_));
 sky130_fd_sc_hd__a21o_1 _17030_ (.A1(_09545_),
    .A2(_09556_),
    .B1(_09555_),
    .X(_09635_));
 sky130_fd_sc_hd__o21a_1 _17031_ (.A1(_09470_),
    .A2(_09533_),
    .B1(_09468_),
    .X(_09636_));
 sky130_fd_sc_hd__nor2_1 _17032_ (.A(_09007_),
    .B(_09036_),
    .Y(_09637_));
 sky130_fd_sc_hd__o22ai_1 _17033_ (.A1(_09007_),
    .A2(_09035_),
    .B1(_09036_),
    .B2(_09009_),
    .Y(_09638_));
 sky130_fd_sc_hd__a21bo_1 _17034_ (.A1(_09541_),
    .A2(_09637_),
    .B1_N(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__nor2_1 _17035_ (.A(_08889_),
    .B(_09039_),
    .Y(_09640_));
 sky130_fd_sc_hd__xor2_2 _17036_ (.A(_09639_),
    .B(_09640_),
    .X(_09641_));
 sky130_fd_sc_hd__a21oi_1 _17037_ (.A1(_09014_),
    .A2(_09016_),
    .B1(_08803_),
    .Y(_09642_));
 sky130_fd_sc_hd__nand2_1 _17038_ (.A(_09547_),
    .B(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__nor2_1 _17039_ (.A(_09021_),
    .B(_09046_),
    .Y(_09644_));
 sky130_fd_sc_hd__xnor2_1 _17040_ (.A(_09643_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__o21a_1 _17041_ (.A1(_09548_),
    .A2(_09551_),
    .B1(_09645_),
    .X(_09646_));
 sky130_fd_sc_hd__nor3_1 _17042_ (.A(_09548_),
    .B(_09551_),
    .C(_09645_),
    .Y(_09647_));
 sky130_fd_sc_hd__nor2_1 _17043_ (.A(_09646_),
    .B(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__xnor2_1 _17044_ (.A(_09641_),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__xnor2_1 _17045_ (.A(_09636_),
    .B(_09649_),
    .Y(_09650_));
 sky130_fd_sc_hd__and2_1 _17046_ (.A(_09635_),
    .B(_09650_),
    .X(_09651_));
 sky130_fd_sc_hd__nor2_1 _17047_ (.A(_09635_),
    .B(_09650_),
    .Y(_09652_));
 sky130_fd_sc_hd__nor2_1 _17048_ (.A(_09651_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__o21ai_1 _17049_ (.A1(_09280_),
    .A2(_09634_),
    .B1(_09653_),
    .Y(_09654_));
 sky130_fd_sc_hd__o21ba_1 _17050_ (.A1(_09280_),
    .A2(_09634_),
    .B1_N(_09633_),
    .X(_09655_));
 sky130_fd_sc_hd__o22a_1 _17051_ (.A1(_09633_),
    .A2(_09654_),
    .B1(_09655_),
    .B2(_09653_),
    .X(_09656_));
 sky130_fd_sc_hd__xnor2_1 _17052_ (.A(_09632_),
    .B(_09656_),
    .Y(_09657_));
 sky130_fd_sc_hd__o21ai_1 _17053_ (.A1(_09589_),
    .A2(_09590_),
    .B1(_09592_),
    .Y(_09658_));
 sky130_fd_sc_hd__or2b_1 _17054_ (.A(_09559_),
    .B_N(_09537_),
    .X(_09659_));
 sky130_fd_sc_hd__a21bo_1 _17055_ (.A1(_09539_),
    .A2(_09558_),
    .B1_N(_09659_),
    .X(_09660_));
 sky130_fd_sc_hd__or2_1 _17056_ (.A(_08899_),
    .B(_07961_),
    .X(_09661_));
 sky130_fd_sc_hd__or2_1 _17057_ (.A(_08896_),
    .B(_08071_),
    .X(_09662_));
 sky130_fd_sc_hd__o22a_1 _17058_ (.A1(_08896_),
    .A2(_07961_),
    .B1(_08071_),
    .B2(_08899_),
    .X(_09663_));
 sky130_fd_sc_hd__o21ba_1 _17059_ (.A1(_09661_),
    .A2(_09662_),
    .B1_N(_09663_),
    .X(_09664_));
 sky130_fd_sc_hd__nor2_1 _17060_ (.A(_08862_),
    .B(_08333_),
    .Y(_09665_));
 sky130_fd_sc_hd__xnor2_1 _17061_ (.A(_09664_),
    .B(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__o31a_1 _17062_ (.A1(_08888_),
    .A2(_08333_),
    .A3(_09568_),
    .B1(_09567_),
    .X(_09667_));
 sky130_fd_sc_hd__nor2_1 _17063_ (.A(_09666_),
    .B(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__and2_1 _17064_ (.A(_09666_),
    .B(_09667_),
    .X(_09669_));
 sky130_fd_sc_hd__nor2_1 _17065_ (.A(_09668_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__nand2_1 _17066_ (.A(_08888_),
    .B(_08317_),
    .Y(_09671_));
 sky130_fd_sc_hd__xnor2_2 _17067_ (.A(_09670_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__o31a_1 _17068_ (.A1(_08896_),
    .A2(_09110_),
    .A3(_09583_),
    .B1(_09581_),
    .X(_09673_));
 sky130_fd_sc_hd__o31ai_1 _17069_ (.A1(_08889_),
    .A2(_09256_),
    .A3(_09543_),
    .B1(_09542_),
    .Y(_09674_));
 sky130_fd_sc_hd__nor2_1 _17070_ (.A(_09256_),
    .B(_09229_),
    .Y(_09675_));
 sky130_fd_sc_hd__o22a_1 _17071_ (.A1(_09231_),
    .A2(_09256_),
    .B1(_09229_),
    .B2(_09142_),
    .X(_09676_));
 sky130_fd_sc_hd__a41o_1 _17072_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_07256_),
    .A3(_07173_),
    .A4(_09675_),
    .B1(_09676_),
    .X(_09677_));
 sky130_fd_sc_hd__nor2_1 _17073_ (.A(_09133_),
    .B(_09110_),
    .Y(_09678_));
 sky130_fd_sc_hd__xnor2_1 _17074_ (.A(_09677_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__xor2_1 _17075_ (.A(_09674_),
    .B(_09679_),
    .X(_09680_));
 sky130_fd_sc_hd__and2b_1 _17076_ (.A_N(_09673_),
    .B(_09680_),
    .X(_09681_));
 sky130_fd_sc_hd__and2b_1 _17077_ (.A_N(_09680_),
    .B(_09673_),
    .X(_09682_));
 sky130_fd_sc_hd__or2_1 _17078_ (.A(_09681_),
    .B(_09682_),
    .X(_09683_));
 sky130_fd_sc_hd__a21o_1 _17079_ (.A1(_09578_),
    .A2(_09588_),
    .B1(_09586_),
    .X(_09684_));
 sky130_fd_sc_hd__xnor2_1 _17080_ (.A(_09683_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__xor2_1 _17081_ (.A(_09672_),
    .B(_09685_),
    .X(_09686_));
 sky130_fd_sc_hd__nand2_1 _17082_ (.A(_09660_),
    .B(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__or2_1 _17083_ (.A(_09660_),
    .B(_09686_),
    .X(_09688_));
 sky130_fd_sc_hd__and2_1 _17084_ (.A(_09687_),
    .B(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__xor2_1 _17085_ (.A(_09658_),
    .B(_09689_),
    .X(_09690_));
 sky130_fd_sc_hd__xor2_1 _17086_ (.A(_09657_),
    .B(_09690_),
    .X(_09691_));
 sky130_fd_sc_hd__o21a_1 _17087_ (.A1(_09561_),
    .A2(_09562_),
    .B1(_09599_),
    .X(_09692_));
 sky130_fd_sc_hd__xnor2_1 _17088_ (.A(_09691_),
    .B(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__and2b_1 _17089_ (.A_N(_09597_),
    .B(_09564_),
    .X(_09694_));
 sky130_fd_sc_hd__a21oi_1 _17090_ (.A1(_09575_),
    .A2(_09576_),
    .B1(_09573_),
    .Y(_09695_));
 sky130_fd_sc_hd__o21ba_1 _17091_ (.A1(_09595_),
    .A2(_09694_),
    .B1_N(_09695_),
    .X(_09696_));
 sky130_fd_sc_hd__or3b_1 _17092_ (.A(_09595_),
    .B(_09694_),
    .C_N(_09695_),
    .X(_09697_));
 sky130_fd_sc_hd__and2b_1 _17093_ (.A_N(_09696_),
    .B(_09697_),
    .X(_09698_));
 sky130_fd_sc_hd__xor2_1 _17094_ (.A(_09693_),
    .B(_09698_),
    .X(_09699_));
 sky130_fd_sc_hd__a21oi_1 _17095_ (.A1(_09630_),
    .A2(_09604_),
    .B1(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__and3_1 _17096_ (.A(_09630_),
    .B(_09604_),
    .C(_09699_),
    .X(_09701_));
 sky130_fd_sc_hd__nor2_1 _17097_ (.A(_09700_),
    .B(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__xnor2_1 _17098_ (.A(_09529_),
    .B(_09702_),
    .Y(_09703_));
 sky130_fd_sc_hd__a21o_1 _17099_ (.A1(_09629_),
    .A2(_09609_),
    .B1(_09703_),
    .X(_09704_));
 sky130_fd_sc_hd__nand3_1 _17100_ (.A(_09629_),
    .B(_09609_),
    .C(_09703_),
    .Y(_09705_));
 sky130_fd_sc_hd__and2_1 _17101_ (.A(_09704_),
    .B(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__a21o_1 _17102_ (.A1(_09615_),
    .A2(_09619_),
    .B1(_09613_),
    .X(_09707_));
 sky130_fd_sc_hd__a21oi_1 _17103_ (.A1(_09706_),
    .A2(_09707_),
    .B1(_08509_),
    .Y(_09708_));
 sky130_fd_sc_hd__o21ai_2 _17104_ (.A1(_09706_),
    .A2(_09707_),
    .B1(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__nand2_1 _17105_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_09710_));
 sky130_fd_sc_hd__or2_1 _17106_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_09711_));
 sky130_fd_sc_hd__a21bo_1 _17107_ (.A1(_09623_),
    .A2(_09625_),
    .B1_N(_09624_),
    .X(_09712_));
 sky130_fd_sc_hd__a21oi_1 _17108_ (.A1(_09710_),
    .A2(_09711_),
    .B1(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__a31o_1 _17109_ (.A1(_09710_),
    .A2(_09711_),
    .A3(_09712_),
    .B1(_04946_),
    .X(_09714_));
 sky130_fd_sc_hd__o21a_1 _17110_ (.A1(_09713_),
    .A2(_09714_),
    .B1(_08507_),
    .X(_09715_));
 sky130_fd_sc_hd__o2bb2a_1 _17111_ (.A1_N(_09709_),
    .A2_N(_09715_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_08508_),
    .X(_00558_));
 sky130_fd_sc_hd__a21bo_1 _17112_ (.A1(_09613_),
    .A2(_09705_),
    .B1_N(_09704_),
    .X(_09716_));
 sky130_fd_sc_hd__a31o_1 _17113_ (.A1(_09615_),
    .A2(_09619_),
    .A3(_09706_),
    .B1(_09716_),
    .X(_01457_));
 sky130_fd_sc_hd__a21oi_2 _17114_ (.A1(_09529_),
    .A2(_09702_),
    .B1(_09700_),
    .Y(_01458_));
 sky130_fd_sc_hd__or2b_1 _17115_ (.A(_09693_),
    .B_N(_09698_),
    .X(_01459_));
 sky130_fd_sc_hd__o21a_1 _17116_ (.A1(_09691_),
    .A2(_09692_),
    .B1(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__or2b_1 _17117_ (.A(_09633_),
    .B_N(_09654_),
    .X(_01461_));
 sky130_fd_sc_hd__inv_2 _17118_ (.A(_09649_),
    .Y(_01462_));
 sky130_fd_sc_hd__o21ba_1 _17119_ (.A1(_09636_),
    .A2(_01462_),
    .B1_N(_09651_),
    .X(_01463_));
 sky130_fd_sc_hd__nand2_1 _17120_ (.A(_08862_),
    .B(_08317_),
    .Y(_01464_));
 sky130_fd_sc_hd__xor2_1 _17121_ (.A(_09636_),
    .B(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__xnor2_1 _17122_ (.A(_01463_),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__nor2_1 _17123_ (.A(_08899_),
    .B(_08333_),
    .Y(_01467_));
 sky130_fd_sc_hd__a31o_1 _17124_ (.A1(_08888_),
    .A2(_08317_),
    .A3(_09670_),
    .B1(_09668_),
    .X(_01468_));
 sky130_fd_sc_hd__or4_1 _17125_ (.A(_09142_),
    .B(_09231_),
    .C(_09256_),
    .D(_09229_),
    .X(_01469_));
 sky130_fd_sc_hd__o31a_1 _17126_ (.A1(_09133_),
    .A2(_09110_),
    .A3(_09676_),
    .B1(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__xor2_1 _17127_ (.A(_01468_),
    .B(_01470_),
    .X(_01471_));
 sky130_fd_sc_hd__xnor2_2 _17128_ (.A(_01467_),
    .B(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__xnor2_1 _17129_ (.A(_01466_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__xnor2_2 _17130_ (.A(_01461_),
    .B(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__and2b_1 _17131_ (.A_N(_09657_),
    .B(_09690_),
    .X(_01475_));
 sky130_fd_sc_hd__a21oi_1 _17132_ (.A1(_09632_),
    .A2(_09656_),
    .B1(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__a21bo_1 _17133_ (.A1(_09658_),
    .A2(_09689_),
    .B1_N(_09687_),
    .X(_01477_));
 sky130_fd_sc_hd__and2b_1 _17134_ (.A_N(_09683_),
    .B(_09684_),
    .X(_01478_));
 sky130_fd_sc_hd__a21o_1 _17135_ (.A1(_09672_),
    .A2(_09685_),
    .B1(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__o32a_1 _17136_ (.A1(_08862_),
    .A2(_08333_),
    .A3(_09663_),
    .B1(_09662_),
    .B2(_09661_),
    .X(_01480_));
 sky130_fd_sc_hd__xnor2_1 _17137_ (.A(_01479_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__a22o_1 _17138_ (.A1(_09541_),
    .A2(_09637_),
    .B1(_09638_),
    .B2(_09640_),
    .X(_01482_));
 sky130_fd_sc_hd__nor2_1 _17139_ (.A(_09009_),
    .B(_09046_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _17140_ (.A(_09133_),
    .B(_07961_),
    .Y(_01484_));
 sky130_fd_sc_hd__xnor2_2 _17141_ (.A(_09662_),
    .B(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__xnor2_1 _17142_ (.A(_09637_),
    .B(_01485_),
    .Y(_01486_));
 sky130_fd_sc_hd__xnor2_1 _17143_ (.A(_01483_),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__xnor2_1 _17144_ (.A(_01482_),
    .B(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__or2_1 _17145_ (.A(_09231_),
    .B(_09039_),
    .X(_01489_));
 sky130_fd_sc_hd__inv_2 _17146_ (.A(_09641_),
    .Y(_01490_));
 sky130_fd_sc_hd__a21oi_1 _17147_ (.A1(_01490_),
    .A2(_09648_),
    .B1(_09646_),
    .Y(_01491_));
 sky130_fd_sc_hd__xnor2_1 _17148_ (.A(_01489_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__xnor2_1 _17149_ (.A(_01488_),
    .B(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__xnor2_1 _17150_ (.A(_01481_),
    .B(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__a21oi_1 _17151_ (.A1(_09674_),
    .A2(_09679_),
    .B1(_09681_),
    .Y(_01495_));
 sky130_fd_sc_hd__o21ai_1 _17152_ (.A1(_09021_),
    .A2(_09046_),
    .B1(_09642_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_1 _17153_ (.A(_09547_),
    .B(_01496_),
    .Y(_01497_));
 sky130_fd_sc_hd__nor2_1 _17154_ (.A(_09142_),
    .B(_09110_),
    .Y(_01498_));
 sky130_fd_sc_hd__or2_1 _17155_ (.A(_09021_),
    .B(_08803_),
    .X(_01499_));
 sky130_fd_sc_hd__nor2_1 _17156_ (.A(_08889_),
    .B(_09035_),
    .Y(_01500_));
 sky130_fd_sc_hd__xnor2_1 _17157_ (.A(_09675_),
    .B(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__xnor2_1 _17158_ (.A(_01499_),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__xnor2_1 _17159_ (.A(_01498_),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__xnor2_1 _17160_ (.A(_01497_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__xnor2_1 _17161_ (.A(_01495_),
    .B(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__xnor2_1 _17162_ (.A(_01494_),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__xnor2_1 _17163_ (.A(_01477_),
    .B(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__xnor2_1 _17164_ (.A(_09696_),
    .B(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__xnor2_1 _17165_ (.A(_01476_),
    .B(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__xnor2_2 _17166_ (.A(_01474_),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__xnor2_4 _17167_ (.A(_01460_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__xnor2_4 _17168_ (.A(_01458_),
    .B(_01511_),
    .Y(_01512_));
 sky130_fd_sc_hd__a21oi_1 _17169_ (.A1(_01457_),
    .A2(_01512_),
    .B1(_08509_),
    .Y(_01513_));
 sky130_fd_sc_hd__o21ai_2 _17170_ (.A1(_01457_),
    .A2(_01512_),
    .B1(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__a21bo_1 _17171_ (.A1(_09711_),
    .A2(_09712_),
    .B1_N(_09710_),
    .X(_01515_));
 sky130_fd_sc_hd__or2_1 _17172_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .X(_01516_));
 sky130_fd_sc_hd__nand2_1 _17173_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_01517_));
 sky130_fd_sc_hd__and3_1 _17174_ (.A(_01515_),
    .B(_01516_),
    .C(_01517_),
    .X(_01518_));
 sky130_fd_sc_hd__a21oi_1 _17175_ (.A1(_01516_),
    .A2(_01517_),
    .B1(_01515_),
    .Y(_01519_));
 sky130_fd_sc_hd__o31a_1 _17176_ (.A1(_08524_),
    .A2(_01518_),
    .A3(_01519_),
    .B1(_08507_),
    .X(_01520_));
 sky130_fd_sc_hd__o2bb2a_1 _17177_ (.A1_N(_01514_),
    .A2_N(_01520_),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_08508_),
    .X(_00559_));
 sky130_fd_sc_hd__and3_1 _17178_ (.A(_03483_),
    .B(_03458_),
    .C(_05005_),
    .X(_01521_));
 sky130_fd_sc_hd__o21a_2 _17179_ (.A1(\rbzero.wall_tracer.state[1] ),
    .A2(_03493_),
    .B1(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__clkbuf_4 _17180_ (.A(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_01524_));
 sky130_fd_sc_hd__or2_1 _17182_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_01525_));
 sky130_fd_sc_hd__o21ai_4 _17183_ (.A1(\rbzero.wall_tracer.state[1] ),
    .A2(_03493_),
    .B1(_01521_),
    .Y(_01526_));
 sky130_fd_sc_hd__buf_4 _17184_ (.A(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__a31o_1 _17185_ (.A1(_08562_),
    .A2(_01524_),
    .A3(_01525_),
    .B1(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__o22a_1 _17186_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(_01523_),
    .B1(_01528_),
    .B2(_08511_),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _17187_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_01529_));
 sky130_fd_sc_hd__nand2_1 _17188_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_01530_));
 sky130_fd_sc_hd__nand3b_1 _17189_ (.A_N(_01524_),
    .B(_01529_),
    .C(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__a21bo_1 _17190_ (.A1(_01529_),
    .A2(_01530_),
    .B1_N(_01524_),
    .X(_01532_));
 sky130_fd_sc_hd__a31o_1 _17191_ (.A1(_08562_),
    .A2(_01531_),
    .A3(_01532_),
    .B1(_01527_),
    .X(_01533_));
 sky130_fd_sc_hd__o22a_1 _17192_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(_01523_),
    .B1(_01533_),
    .B2(_08517_),
    .X(_00561_));
 sky130_fd_sc_hd__clkbuf_4 _17193_ (.A(_08509_),
    .X(_01534_));
 sky130_fd_sc_hd__and2_1 _17194_ (.A(_01530_),
    .B(_01531_),
    .X(_01535_));
 sky130_fd_sc_hd__nor2_1 _17195_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_01536_));
 sky130_fd_sc_hd__and2_1 _17196_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_01537_));
 sky130_fd_sc_hd__or3_1 _17197_ (.A(_01535_),
    .B(_01536_),
    .C(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__o21ai_1 _17198_ (.A1(_01536_),
    .A2(_01537_),
    .B1(_01535_),
    .Y(_01539_));
 sky130_fd_sc_hd__a31o_1 _17199_ (.A1(_01534_),
    .A2(_01538_),
    .A3(_01539_),
    .B1(_01527_),
    .X(_01540_));
 sky130_fd_sc_hd__o22a_1 _17200_ (.A1(\rbzero.wall_tracer.trackDistY[-9] ),
    .A2(_01523_),
    .B1(_01540_),
    .B2(_08525_),
    .X(_00562_));
 sky130_fd_sc_hd__or2_1 _17201_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_01541_));
 sky130_fd_sc_hd__nand2_1 _17202_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .Y(_01542_));
 sky130_fd_sc_hd__o21bai_1 _17203_ (.A1(_01535_),
    .A2(_01536_),
    .B1_N(_01537_),
    .Y(_01543_));
 sky130_fd_sc_hd__nand3_1 _17204_ (.A(_01541_),
    .B(_01542_),
    .C(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21o_1 _17205_ (.A1(_01541_),
    .A2(_01542_),
    .B1(_01543_),
    .X(_01545_));
 sky130_fd_sc_hd__a31o_1 _17206_ (.A1(_01534_),
    .A2(_01544_),
    .A3(_01545_),
    .B1(_01527_),
    .X(_01546_));
 sky130_fd_sc_hd__o22a_1 _17207_ (.A1(\rbzero.wall_tracer.trackDistY[-8] ),
    .A2(_01523_),
    .B1(_01546_),
    .B2(_08532_),
    .X(_00563_));
 sky130_fd_sc_hd__nor2_1 _17208_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_01547_));
 sky130_fd_sc_hd__and2_1 _17209_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .X(_01548_));
 sky130_fd_sc_hd__a21boi_1 _17210_ (.A1(_01541_),
    .A2(_01543_),
    .B1_N(_01542_),
    .Y(_01549_));
 sky130_fd_sc_hd__or3_1 _17211_ (.A(_01547_),
    .B(_01548_),
    .C(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__o21ai_1 _17212_ (.A1(_01547_),
    .A2(_01548_),
    .B1(_01549_),
    .Y(_01551_));
 sky130_fd_sc_hd__a31o_1 _17213_ (.A1(_01534_),
    .A2(_01550_),
    .A3(_01551_),
    .B1(_01526_),
    .X(_01552_));
 sky130_fd_sc_hd__o22a_1 _17214_ (.A1(\rbzero.wall_tracer.trackDistY[-7] ),
    .A2(_01523_),
    .B1(_01552_),
    .B2(_08539_),
    .X(_00564_));
 sky130_fd_sc_hd__or2_1 _17215_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_01553_));
 sky130_fd_sc_hd__nand2_1 _17216_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .Y(_01554_));
 sky130_fd_sc_hd__o21bai_1 _17217_ (.A1(_01547_),
    .A2(_01549_),
    .B1_N(_01548_),
    .Y(_01555_));
 sky130_fd_sc_hd__a21oi_1 _17218_ (.A1(_01553_),
    .A2(_01554_),
    .B1(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__a31o_1 _17219_ (.A1(_01553_),
    .A2(_01554_),
    .A3(_01555_),
    .B1(_04946_),
    .X(_01557_));
 sky130_fd_sc_hd__clkbuf_4 _17220_ (.A(_01522_),
    .X(_01558_));
 sky130_fd_sc_hd__o21ai_1 _17221_ (.A1(_01556_),
    .A2(_01557_),
    .B1(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__o22a_1 _17222_ (.A1(\rbzero.wall_tracer.trackDistY[-6] ),
    .A2(_01523_),
    .B1(_01559_),
    .B2(_08546_),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _17223_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_01560_));
 sky130_fd_sc_hd__and2_1 _17224_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .X(_01561_));
 sky130_fd_sc_hd__a21boi_1 _17225_ (.A1(_01553_),
    .A2(_01555_),
    .B1_N(_01554_),
    .Y(_01562_));
 sky130_fd_sc_hd__or3_1 _17226_ (.A(_01560_),
    .B(_01561_),
    .C(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__o21ai_1 _17227_ (.A1(_01560_),
    .A2(_01561_),
    .B1(_01562_),
    .Y(_01564_));
 sky130_fd_sc_hd__a31o_1 _17228_ (.A1(_01534_),
    .A2(_01563_),
    .A3(_01564_),
    .B1(_01526_),
    .X(_01565_));
 sky130_fd_sc_hd__o22a_1 _17229_ (.A1(\rbzero.wall_tracer.trackDistY[-5] ),
    .A2(_01523_),
    .B1(_01565_),
    .B2(_08554_),
    .X(_00566_));
 sky130_fd_sc_hd__or2_1 _17230_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(_01566_));
 sky130_fd_sc_hd__nand2_1 _17231_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_01567_));
 sky130_fd_sc_hd__o21bai_1 _17232_ (.A1(_01560_),
    .A2(_01562_),
    .B1_N(_01561_),
    .Y(_01568_));
 sky130_fd_sc_hd__a21oi_1 _17233_ (.A1(_01566_),
    .A2(_01567_),
    .B1(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__a31o_1 _17234_ (.A1(_01566_),
    .A2(_01567_),
    .A3(_01568_),
    .B1(_04946_),
    .X(_01570_));
 sky130_fd_sc_hd__o21ai_1 _17235_ (.A1(_01569_),
    .A2(_01570_),
    .B1(_01558_),
    .Y(_01571_));
 sky130_fd_sc_hd__o22a_1 _17236_ (.A1(\rbzero.wall_tracer.trackDistY[-4] ),
    .A2(_01558_),
    .B1(_01571_),
    .B2(_08561_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _17237_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_01572_));
 sky130_fd_sc_hd__and2_1 _17238_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .X(_01573_));
 sky130_fd_sc_hd__a21boi_1 _17239_ (.A1(_01566_),
    .A2(_01568_),
    .B1_N(_01567_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor3_1 _17240_ (.A(_01572_),
    .B(_01573_),
    .C(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__o21a_1 _17241_ (.A1(_01572_),
    .A2(_01573_),
    .B1(_01574_),
    .X(_01576_));
 sky130_fd_sc_hd__o311a_1 _17242_ (.A1(_08485_),
    .A2(_01575_),
    .A3(_01576_),
    .B1(_08575_),
    .C1(_01522_),
    .X(_01577_));
 sky130_fd_sc_hd__a21oi_1 _17243_ (.A1(_04986_),
    .A2(_01527_),
    .B1(_01577_),
    .Y(_00568_));
 sky130_fd_sc_hd__or2_1 _17244_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_01578_));
 sky130_fd_sc_hd__nand2_1 _17245_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_01579_));
 sky130_fd_sc_hd__o21bai_1 _17246_ (.A1(_01572_),
    .A2(_01574_),
    .B1_N(_01573_),
    .Y(_01580_));
 sky130_fd_sc_hd__nand3_1 _17247_ (.A(_01578_),
    .B(_01579_),
    .C(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__a21o_1 _17248_ (.A1(_01578_),
    .A2(_01579_),
    .B1(_01580_),
    .X(_01582_));
 sky130_fd_sc_hd__a31o_1 _17249_ (.A1(_01534_),
    .A2(_01581_),
    .A3(_01582_),
    .B1(_01526_),
    .X(_01583_));
 sky130_fd_sc_hd__o22a_1 _17250_ (.A1(\rbzero.wall_tracer.trackDistY[-2] ),
    .A2(_01558_),
    .B1(_01583_),
    .B2(_08577_),
    .X(_00569_));
 sky130_fd_sc_hd__nor2_1 _17251_ (.A(_04964_),
    .B(_07115_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _17252_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_01585_));
 sky130_fd_sc_hd__a21boi_1 _17253_ (.A1(_01578_),
    .A2(_01580_),
    .B1_N(_01579_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor3_1 _17254_ (.A(_01584_),
    .B(_01585_),
    .C(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__o21a_1 _17255_ (.A1(_01584_),
    .A2(_01585_),
    .B1(_01586_),
    .X(_01588_));
 sky130_fd_sc_hd__o311a_1 _17256_ (.A1(_08485_),
    .A2(_01587_),
    .A3(_01588_),
    .B1(_08584_),
    .C1(_01522_),
    .X(_01589_));
 sky130_fd_sc_hd__a21oi_1 _17257_ (.A1(_04964_),
    .A2(_01527_),
    .B1(_01589_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _17258_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_01590_));
 sky130_fd_sc_hd__or2_1 _17259_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .X(_01591_));
 sky130_fd_sc_hd__o211a_1 _17260_ (.A1(_01584_),
    .A2(_01587_),
    .B1(_01590_),
    .C1(_01591_),
    .X(_01592_));
 sky130_fd_sc_hd__a211oi_1 _17261_ (.A1(_01590_),
    .A2(_01591_),
    .B1(_01584_),
    .C1(_01587_),
    .Y(_01593_));
 sky130_fd_sc_hd__o311a_1 _17262_ (.A1(_04946_),
    .A2(_01592_),
    .A3(_01593_),
    .B1(_08717_),
    .C1(_01522_),
    .X(_01594_));
 sky130_fd_sc_hd__a21oi_1 _17263_ (.A1(_04963_),
    .A2(_01527_),
    .B1(_01594_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _17264_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_01595_));
 sky130_fd_sc_hd__or2_1 _17265_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_01596_));
 sky130_fd_sc_hd__a21o_1 _17266_ (.A1(\rbzero.wall_tracer.trackDistY[0] ),
    .A2(\rbzero.wall_tracer.stepDistY[0] ),
    .B1(_01592_),
    .X(_01597_));
 sky130_fd_sc_hd__and3_1 _17267_ (.A(_01595_),
    .B(_01596_),
    .C(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__inv_2 _17268_ (.A(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__a21o_1 _17269_ (.A1(_01595_),
    .A2(_01596_),
    .B1(_01597_),
    .X(_01600_));
 sky130_fd_sc_hd__a31o_1 _17270_ (.A1(_01534_),
    .A2(_01599_),
    .A3(_01600_),
    .B1(_01526_),
    .X(_01601_));
 sky130_fd_sc_hd__o22a_1 _17271_ (.A1(\rbzero.wall_tracer.trackDistY[1] ),
    .A2(_01558_),
    .B1(_01601_),
    .B2(_08835_),
    .X(_00572_));
 sky130_fd_sc_hd__nand2_1 _17272_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_01602_));
 sky130_fd_sc_hd__or2_1 _17273_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_01603_));
 sky130_fd_sc_hd__nand2_1 _17274_ (.A(_01595_),
    .B(_01599_),
    .Y(_01604_));
 sky130_fd_sc_hd__a21o_1 _17275_ (.A1(_01602_),
    .A2(_01603_),
    .B1(_01604_),
    .X(_01605_));
 sky130_fd_sc_hd__and3_1 _17276_ (.A(_01602_),
    .B(_01603_),
    .C(_01604_),
    .X(_01606_));
 sky130_fd_sc_hd__inv_2 _17277_ (.A(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__a31o_1 _17278_ (.A1(_01534_),
    .A2(_01605_),
    .A3(_01607_),
    .B1(_01526_),
    .X(_01608_));
 sky130_fd_sc_hd__o22a_1 _17279_ (.A1(\rbzero.wall_tracer.trackDistY[2] ),
    .A2(_01558_),
    .B1(_01608_),
    .B2(_08959_),
    .X(_00573_));
 sky130_fd_sc_hd__nand2_1 _17280_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_01609_));
 sky130_fd_sc_hd__or2_1 _17281_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_01610_));
 sky130_fd_sc_hd__nand2_1 _17282_ (.A(_01602_),
    .B(_01607_),
    .Y(_01611_));
 sky130_fd_sc_hd__and3_1 _17283_ (.A(_01609_),
    .B(_01610_),
    .C(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__inv_2 _17284_ (.A(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hd__a21o_1 _17285_ (.A1(_01609_),
    .A2(_01610_),
    .B1(_01611_),
    .X(_01614_));
 sky130_fd_sc_hd__a31o_1 _17286_ (.A1(_01534_),
    .A2(_01613_),
    .A3(_01614_),
    .B1(_01526_),
    .X(_01615_));
 sky130_fd_sc_hd__o22a_1 _17287_ (.A1(\rbzero.wall_tracer.trackDistY[3] ),
    .A2(_01558_),
    .B1(_01615_),
    .B2(_09081_),
    .X(_00574_));
 sky130_fd_sc_hd__nand2_1 _17288_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .Y(_01616_));
 sky130_fd_sc_hd__or2_1 _17289_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_01617_));
 sky130_fd_sc_hd__nand2_1 _17290_ (.A(_01616_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _17291_ (.A(_01609_),
    .B(_01613_),
    .Y(_01619_));
 sky130_fd_sc_hd__xnor2_1 _17292_ (.A(_01618_),
    .B(_01619_),
    .Y(_01620_));
 sky130_fd_sc_hd__a21o_1 _17293_ (.A1(_08512_),
    .A2(_01620_),
    .B1(_01527_),
    .X(_01621_));
 sky130_fd_sc_hd__o22a_1 _17294_ (.A1(\rbzero.wall_tracer.trackDistY[4] ),
    .A2(_01558_),
    .B1(_01621_),
    .B2(_09197_),
    .X(_00575_));
 sky130_fd_sc_hd__nor2_1 _17295_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_01622_));
 sky130_fd_sc_hd__and2_1 _17296_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_01623_));
 sky130_fd_sc_hd__a21boi_2 _17297_ (.A1(_01617_),
    .A2(_01619_),
    .B1_N(_01616_),
    .Y(_01624_));
 sky130_fd_sc_hd__or3_1 _17298_ (.A(_01622_),
    .B(_01623_),
    .C(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__o21ai_1 _17299_ (.A1(_01622_),
    .A2(_01623_),
    .B1(_01624_),
    .Y(_01626_));
 sky130_fd_sc_hd__a31o_1 _17300_ (.A1(_01534_),
    .A2(_01625_),
    .A3(_01626_),
    .B1(_01526_),
    .X(_01627_));
 sky130_fd_sc_hd__o22a_1 _17301_ (.A1(\rbzero.wall_tracer.trackDistY[5] ),
    .A2(_01558_),
    .B1(_01627_),
    .B2(_09308_),
    .X(_00576_));
 sky130_fd_sc_hd__nor2_1 _17302_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_01628_));
 sky130_fd_sc_hd__and2_1 _17303_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .X(_01629_));
 sky130_fd_sc_hd__o21ba_1 _17304_ (.A1(_01622_),
    .A2(_01624_),
    .B1_N(_01623_),
    .X(_01630_));
 sky130_fd_sc_hd__or3_1 _17305_ (.A(_01628_),
    .B(_01629_),
    .C(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__o21ai_1 _17306_ (.A1(_01628_),
    .A2(_01629_),
    .B1(_01630_),
    .Y(_01632_));
 sky130_fd_sc_hd__a31o_1 _17307_ (.A1(_01534_),
    .A2(_01631_),
    .A3(_01632_),
    .B1(_01526_),
    .X(_01633_));
 sky130_fd_sc_hd__o22a_1 _17308_ (.A1(\rbzero.wall_tracer.trackDistY[6] ),
    .A2(_01558_),
    .B1(_01633_),
    .B2(_09416_),
    .X(_00577_));
 sky130_fd_sc_hd__nor2_1 _17309_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_01634_));
 sky130_fd_sc_hd__nand2_1 _17310_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_01635_));
 sky130_fd_sc_hd__and2b_1 _17311_ (.A_N(_01634_),
    .B(_01635_),
    .X(_01636_));
 sky130_fd_sc_hd__o21ba_1 _17312_ (.A1(_01628_),
    .A2(_01630_),
    .B1_N(_01629_),
    .X(_01637_));
 sky130_fd_sc_hd__xnor2_1 _17313_ (.A(_01636_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__a21oi_1 _17314_ (.A1(_08512_),
    .A2(_01638_),
    .B1(_01527_),
    .Y(_01639_));
 sky130_fd_sc_hd__o2bb2a_1 _17315_ (.A1_N(_01639_),
    .A2_N(_09520_),
    .B1(\rbzero.wall_tracer.trackDistY[7] ),
    .B2(_01523_),
    .X(_00578_));
 sky130_fd_sc_hd__or2_1 _17316_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .X(_01640_));
 sky130_fd_sc_hd__nand2_1 _17317_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_01641_));
 sky130_fd_sc_hd__o21ai_1 _17318_ (.A1(_01634_),
    .A2(_01637_),
    .B1(_01635_),
    .Y(_01642_));
 sky130_fd_sc_hd__a21oi_1 _17319_ (.A1(_01640_),
    .A2(_01641_),
    .B1(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__a31o_1 _17320_ (.A1(_01640_),
    .A2(_01641_),
    .A3(_01642_),
    .B1(_03341_),
    .X(_01644_));
 sky130_fd_sc_hd__o211a_1 _17321_ (.A1(_01643_),
    .A2(_01644_),
    .B1(_09622_),
    .C1(_01522_),
    .X(_01645_));
 sky130_fd_sc_hd__a21oi_1 _17322_ (.A1(_04956_),
    .A2(_01527_),
    .B1(_01645_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _17323_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_01646_));
 sky130_fd_sc_hd__or2_1 _17324_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_01647_));
 sky130_fd_sc_hd__a21bo_1 _17325_ (.A1(_01640_),
    .A2(_01642_),
    .B1_N(_01641_),
    .X(_01648_));
 sky130_fd_sc_hd__a21oi_1 _17326_ (.A1(_01646_),
    .A2(_01647_),
    .B1(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__a31o_1 _17327_ (.A1(_01646_),
    .A2(_01647_),
    .A3(_01648_),
    .B1(_03341_),
    .X(_01650_));
 sky130_fd_sc_hd__o21a_1 _17328_ (.A1(_01649_),
    .A2(_01650_),
    .B1(_01522_),
    .X(_01651_));
 sky130_fd_sc_hd__o2bb2a_1 _17329_ (.A1_N(_01651_),
    .A2_N(_09709_),
    .B1(\rbzero.wall_tracer.trackDistY[9] ),
    .B2(_01523_),
    .X(_00580_));
 sky130_fd_sc_hd__a21bo_1 _17330_ (.A1(_01647_),
    .A2(_01648_),
    .B1_N(_01646_),
    .X(_01652_));
 sky130_fd_sc_hd__or2_1 _17331_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .X(_01653_));
 sky130_fd_sc_hd__nand2_1 _17332_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .Y(_01654_));
 sky130_fd_sc_hd__and3_1 _17333_ (.A(_01652_),
    .B(_01653_),
    .C(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__a21oi_1 _17334_ (.A1(_01653_),
    .A2(_01654_),
    .B1(_01652_),
    .Y(_01656_));
 sky130_fd_sc_hd__o31a_1 _17335_ (.A1(_08485_),
    .A2(_01655_),
    .A3(_01656_),
    .B1(_01522_),
    .X(_01657_));
 sky130_fd_sc_hd__o2bb2a_1 _17336_ (.A1_N(_01657_),
    .A2_N(_01514_),
    .B1(\rbzero.wall_tracer.trackDistY[10] ),
    .B2(_01523_),
    .X(_00581_));
 sky130_fd_sc_hd__inv_2 _17337_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .Y(_01658_));
 sky130_fd_sc_hd__or4b_2 _17338_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_01658_),
    .C(\rbzero.spi_registers.spi_cmd[3] ),
    .D_N(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_01659_));
 sky130_fd_sc_hd__inv_2 _17339_ (.A(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__and3_1 _17340_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02907_),
    .C(_01660_),
    .X(_01661_));
 sky130_fd_sc_hd__buf_2 _17341_ (.A(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__clkbuf_4 _17342_ (.A(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _17343_ (.A0(\rbzero.spi_registers.new_mapd[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__clkbuf_1 _17344_ (.A(_01664_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _17345_ (.A0(\rbzero.spi_registers.new_mapd[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_01663_),
    .X(_01665_));
 sky130_fd_sc_hd__clkbuf_1 _17346_ (.A(_01665_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _17347_ (.A0(\rbzero.spi_registers.new_mapd[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_01663_),
    .X(_01666_));
 sky130_fd_sc_hd__clkbuf_1 _17348_ (.A(_01666_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _17349_ (.A0(\rbzero.spi_registers.new_mapd[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_01663_),
    .X(_01667_));
 sky130_fd_sc_hd__clkbuf_1 _17350_ (.A(_01667_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _17351_ (.A0(\rbzero.spi_registers.new_mapd[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_01663_),
    .X(_01668_));
 sky130_fd_sc_hd__clkbuf_1 _17352_ (.A(_01668_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _17353_ (.A0(\rbzero.spi_registers.new_mapd[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_01663_),
    .X(_01669_));
 sky130_fd_sc_hd__clkbuf_1 _17354_ (.A(_01669_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _17355_ (.A0(\rbzero.spi_registers.new_mapd[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_01663_),
    .X(_01670_));
 sky130_fd_sc_hd__clkbuf_1 _17356_ (.A(_01670_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _17357_ (.A0(\rbzero.spi_registers.new_mapd[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_01663_),
    .X(_01671_));
 sky130_fd_sc_hd__clkbuf_1 _17358_ (.A(_01671_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _17359_ (.A0(\rbzero.spi_registers.new_mapd[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_01663_),
    .X(_01672_));
 sky130_fd_sc_hd__clkbuf_1 _17360_ (.A(_01672_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _17361_ (.A0(\rbzero.spi_registers.new_mapd[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_01662_),
    .X(_01673_));
 sky130_fd_sc_hd__clkbuf_1 _17362_ (.A(_01673_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _17363_ (.A0(\rbzero.spi_registers.new_mapd[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_01662_),
    .X(_01674_));
 sky130_fd_sc_hd__clkbuf_1 _17364_ (.A(_01674_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _17365_ (.A0(\rbzero.spi_registers.new_mapd[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_01662_),
    .X(_01675_));
 sky130_fd_sc_hd__clkbuf_1 _17366_ (.A(_01675_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _17367_ (.A0(\rbzero.spi_registers.new_mapd[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_01662_),
    .X(_01676_));
 sky130_fd_sc_hd__clkbuf_1 _17368_ (.A(_01676_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _17369_ (.A0(\rbzero.spi_registers.new_mapd[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_01662_),
    .X(_01677_));
 sky130_fd_sc_hd__clkbuf_1 _17370_ (.A(_01677_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _17371_ (.A0(\rbzero.spi_registers.new_mapd[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_01662_),
    .X(_01678_));
 sky130_fd_sc_hd__clkbuf_1 _17372_ (.A(_01678_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _17373_ (.A0(\rbzero.spi_registers.new_mapd[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_01662_),
    .X(_01679_));
 sky130_fd_sc_hd__clkbuf_1 _17374_ (.A(_01679_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _17375_ (.A0(\rbzero.debug_overlay.playerX[0] ),
    .A1(_03373_),
    .S(_09620_),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _17376_ (.A0(_03395_),
    .A1(_01680_),
    .S(_08507_),
    .X(_01681_));
 sky130_fd_sc_hd__clkbuf_1 _17377_ (.A(_01681_),
    .X(_00598_));
 sky130_fd_sc_hd__or2_1 _17378_ (.A(_03395_),
    .B(_08472_),
    .X(_01682_));
 sky130_fd_sc_hd__nor2_1 _17379_ (.A(_03342_),
    .B(_09620_),
    .Y(_01683_));
 sky130_fd_sc_hd__a31o_1 _17380_ (.A1(_08509_),
    .A2(_08473_),
    .A3(_01682_),
    .B1(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _17381_ (.A0(_03343_),
    .A1(_01684_),
    .S(_08507_),
    .X(_01685_));
 sky130_fd_sc_hd__clkbuf_1 _17382_ (.A(_01685_),
    .X(_00599_));
 sky130_fd_sc_hd__xor2_1 _17383_ (.A(_08474_),
    .B(_08477_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _17384_ (.A0(\rbzero.debug_overlay.playerX[2] ),
    .A1(_01686_),
    .S(_09620_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _17385_ (.A0(_03353_),
    .A1(_01687_),
    .S(_08506_),
    .X(_01688_));
 sky130_fd_sc_hd__clkbuf_1 _17386_ (.A(_01688_),
    .X(_00600_));
 sky130_fd_sc_hd__xnor2_1 _17387_ (.A(_03369_),
    .B(_07826_),
    .Y(_01689_));
 sky130_fd_sc_hd__xnor2_1 _17388_ (.A(_08478_),
    .B(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__mux2_1 _17389_ (.A0(\rbzero.debug_overlay.playerX[3] ),
    .A1(_01690_),
    .S(_09620_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _17390_ (.A0(_03369_),
    .A1(_01691_),
    .S(_08506_),
    .X(_01692_));
 sky130_fd_sc_hd__clkbuf_1 _17391_ (.A(_01692_),
    .X(_00601_));
 sky130_fd_sc_hd__xor2_1 _17392_ (.A(_08471_),
    .B(_08480_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _17393_ (.A0(\rbzero.debug_overlay.playerX[4] ),
    .A1(_01693_),
    .S(\rbzero.wall_tracer.state[1] ),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _17394_ (.A0(\rbzero.map_rom.i_col[4] ),
    .A1(_01694_),
    .S(_08506_),
    .X(_01695_));
 sky130_fd_sc_hd__clkbuf_1 _17395_ (.A(_01695_),
    .X(_00602_));
 sky130_fd_sc_hd__a21oi_1 _17396_ (.A1(_08471_),
    .A2(_08480_),
    .B1(_08469_),
    .Y(_01696_));
 sky130_fd_sc_hd__xnor2_1 _17397_ (.A(_08468_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__mux2_1 _17398_ (.A0(\rbzero.debug_overlay.playerX[5] ),
    .A1(_01697_),
    .S(\rbzero.wall_tracer.state[1] ),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _17399_ (.A0(\rbzero.wall_tracer.mapX[5] ),
    .A1(_01698_),
    .S(_08506_),
    .X(_01699_));
 sky130_fd_sc_hd__clkbuf_1 _17400_ (.A(_01699_),
    .X(_00603_));
 sky130_fd_sc_hd__nor2_1 _17401_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_01700_));
 sky130_fd_sc_hd__nand2_1 _17402_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_01701_));
 sky130_fd_sc_hd__and2b_1 _17403_ (.A_N(_01700_),
    .B(_01701_),
    .X(_01702_));
 sky130_fd_sc_hd__or2_1 _17404_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .X(_01703_));
 sky130_fd_sc_hd__nor2_1 _17405_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _17406_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .Y(_01705_));
 sky130_fd_sc_hd__nor2_1 _17407_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_01706_));
 sky130_fd_sc_hd__and2_1 _17408_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_01707_));
 sky130_fd_sc_hd__o21ba_1 _17409_ (.A1(_01705_),
    .A2(_01706_),
    .B1_N(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__nand2_1 _17410_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_01709_));
 sky130_fd_sc_hd__o21ai_1 _17411_ (.A1(_01704_),
    .A2(_01708_),
    .B1(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand2_1 _17412_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .Y(_01711_));
 sky130_fd_sc_hd__a21boi_1 _17413_ (.A1(_01703_),
    .A2(_01710_),
    .B1_N(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__xnor2_1 _17414_ (.A(_01702_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__clkbuf_4 _17415_ (.A(_03340_),
    .X(_01714_));
 sky130_fd_sc_hd__a22o_1 _17416_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_01714_),
    .B1(_08448_),
    .B2(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(_01715_));
 sky130_fd_sc_hd__a21o_1 _17417_ (.A1(_08453_),
    .A2(_01713_),
    .B1(_01715_),
    .X(_00604_));
 sky130_fd_sc_hd__nor2_1 _17418_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .Y(_01716_));
 sky130_fd_sc_hd__and2_1 _17419_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_01717_));
 sky130_fd_sc_hd__o21ai_1 _17420_ (.A1(_01700_),
    .A2(_01712_),
    .B1(_01701_),
    .Y(_01718_));
 sky130_fd_sc_hd__or3_1 _17421_ (.A(_01716_),
    .B(_01717_),
    .C(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__o21ai_1 _17422_ (.A1(_01716_),
    .A2(_01717_),
    .B1(_01718_),
    .Y(_01720_));
 sky130_fd_sc_hd__a21oi_1 _17423_ (.A1(_01719_),
    .A2(_01720_),
    .B1(_03486_),
    .Y(_01721_));
 sky130_fd_sc_hd__clkbuf_4 _17424_ (.A(_03340_),
    .X(_01722_));
 sky130_fd_sc_hd__or2_1 _17425_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_01723_));
 sky130_fd_sc_hd__nand2_1 _17426_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_01724_));
 sky130_fd_sc_hd__a31o_1 _17427_ (.A1(_01722_),
    .A2(_01723_),
    .A3(_01724_),
    .B1(_08460_),
    .X(_01725_));
 sky130_fd_sc_hd__o22a_1 _17428_ (.A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_00013_),
    .B1(_01721_),
    .B2(_01725_),
    .X(_00605_));
 sky130_fd_sc_hd__nor2_1 _17429_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_01726_));
 sky130_fd_sc_hd__and2_1 _17430_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .X(_01727_));
 sky130_fd_sc_hd__or2_1 _17431_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_01728_));
 sky130_fd_sc_hd__a21oi_1 _17432_ (.A1(_01728_),
    .A2(_01718_),
    .B1(_01717_),
    .Y(_01729_));
 sky130_fd_sc_hd__o21ai_1 _17433_ (.A1(_01726_),
    .A2(_01727_),
    .B1(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__o311a_1 _17434_ (.A1(_01726_),
    .A2(_01727_),
    .A3(_01729_),
    .B1(_01730_),
    .C1(_03497_),
    .X(_01731_));
 sky130_fd_sc_hd__or2_1 _17435_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_01723_),
    .X(_01732_));
 sky130_fd_sc_hd__nand2_1 _17436_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_01723_),
    .Y(_01733_));
 sky130_fd_sc_hd__a31o_1 _17437_ (.A1(_01722_),
    .A2(_01732_),
    .A3(_01733_),
    .B1(_08460_),
    .X(_01734_));
 sky130_fd_sc_hd__o22a_1 _17438_ (.A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A2(_00013_),
    .B1(_01731_),
    .B2(_01734_),
    .X(_00606_));
 sky130_fd_sc_hd__nor2_1 _17439_ (.A(_04109_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_01735_));
 sky130_fd_sc_hd__and2_1 _17440_ (.A(_04109_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_01736_));
 sky130_fd_sc_hd__nand2_1 _17441_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_01737_));
 sky130_fd_sc_hd__o21ai_1 _17442_ (.A1(_01726_),
    .A2(_01729_),
    .B1(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__or3_1 _17443_ (.A(_01735_),
    .B(_01736_),
    .C(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__o21ai_1 _17444_ (.A1(_01735_),
    .A2(_01736_),
    .B1(_01738_),
    .Y(_01740_));
 sky130_fd_sc_hd__a21oi_1 _17445_ (.A1(_01739_),
    .A2(_01740_),
    .B1(_03486_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _17446_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_01732_),
    .Y(_01742_));
 sky130_fd_sc_hd__or2_1 _17447_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_01732_),
    .X(_01743_));
 sky130_fd_sc_hd__a31o_1 _17448_ (.A1(_01722_),
    .A2(_01742_),
    .A3(_01743_),
    .B1(_08460_),
    .X(_01744_));
 sky130_fd_sc_hd__o22a_1 _17449_ (.A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A2(_00013_),
    .B1(_01741_),
    .B2(_01744_),
    .X(_00607_));
 sky130_fd_sc_hd__buf_4 _17450_ (.A(_08452_),
    .X(_01745_));
 sky130_fd_sc_hd__or2_1 _17451_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_01746_));
 sky130_fd_sc_hd__nand2_1 _17452_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_01747_));
 sky130_fd_sc_hd__or2_1 _17453_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_01748_));
 sky130_fd_sc_hd__a21o_1 _17454_ (.A1(_01748_),
    .A2(_01738_),
    .B1(_01736_),
    .X(_01749_));
 sky130_fd_sc_hd__nand3_1 _17455_ (.A(_01746_),
    .B(_01747_),
    .C(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__a21o_1 _17456_ (.A1(_01746_),
    .A2(_01747_),
    .B1(_01749_),
    .X(_01751_));
 sky130_fd_sc_hd__inv_2 _17457_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_01752_));
 sky130_fd_sc_hd__o31a_1 _17458_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(\rbzero.debug_overlay.vplaneY[-7] ),
    .A3(\rbzero.debug_overlay.vplaneY[-8] ),
    .B1(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__xor2_1 _17459_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__a22o_1 _17460_ (.A1(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A2(_08447_),
    .B1(_01754_),
    .B2(_01714_),
    .X(_01755_));
 sky130_fd_sc_hd__a31o_1 _17461_ (.A1(_01745_),
    .A2(_01750_),
    .A3(_01751_),
    .B1(_01755_),
    .X(_00608_));
 sky130_fd_sc_hd__a21bo_1 _17462_ (.A1(_01746_),
    .A2(_01749_),
    .B1_N(_01747_),
    .X(_01756_));
 sky130_fd_sc_hd__clkbuf_4 _17463_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_01757_));
 sky130_fd_sc_hd__nor2_1 _17464_ (.A(_01757_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_01758_));
 sky130_fd_sc_hd__and2_1 _17465_ (.A(_01757_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_01759_));
 sky130_fd_sc_hd__or2_1 _17466_ (.A(_01758_),
    .B(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__xnor2_1 _17467_ (.A(_01756_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__or2_1 _17468_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_01762_));
 sky130_fd_sc_hd__nand2_1 _17469_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _17470_ (.A(_01762_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_1 _17471_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_01765_));
 sky130_fd_sc_hd__or2_1 _17472_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(_01743_),
    .X(_01766_));
 sky130_fd_sc_hd__and3_1 _17473_ (.A(_01764_),
    .B(_01765_),
    .C(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__a21o_1 _17474_ (.A1(_01765_),
    .A2(_01766_),
    .B1(_01764_),
    .X(_01768_));
 sky130_fd_sc_hd__nand2_1 _17475_ (.A(_03339_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__o22a_1 _17476_ (.A1(_03340_),
    .A2(_01761_),
    .B1(_01767_),
    .B2(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _17477_ (.A0(\rbzero.wall_tracer.rayAddendY[0] ),
    .A1(_01770_),
    .S(_03509_),
    .X(_01771_));
 sky130_fd_sc_hd__clkbuf_1 _17478_ (.A(_01771_),
    .X(_00609_));
 sky130_fd_sc_hd__nand2_1 _17479_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_01772_));
 sky130_fd_sc_hd__or2_1 _17480_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_01773_));
 sky130_fd_sc_hd__o21a_1 _17481_ (.A1(_01757_),
    .A2(\rbzero.wall_tracer.rayAddendY[0] ),
    .B1(_01756_),
    .X(_01774_));
 sky130_fd_sc_hd__a211o_1 _17482_ (.A1(_01772_),
    .A2(_01773_),
    .B1(_01774_),
    .C1(_01759_),
    .X(_01775_));
 sky130_fd_sc_hd__o211ai_2 _17483_ (.A1(_01759_),
    .A2(_01774_),
    .B1(_01773_),
    .C1(_01772_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor2_1 _17484_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_01777_));
 sky130_fd_sc_hd__and2_1 _17485_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(_01778_));
 sky130_fd_sc_hd__nor2_1 _17486_ (.A(_01777_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__xnor2_1 _17487_ (.A(_01762_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__a21bo_1 _17488_ (.A1(_01764_),
    .A2(_01766_),
    .B1_N(_01765_),
    .X(_01781_));
 sky130_fd_sc_hd__xnor2_1 _17489_ (.A(_01780_),
    .B(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__a22o_1 _17490_ (.A1(\rbzero.wall_tracer.rayAddendY[1] ),
    .A2(_08447_),
    .B1(_01782_),
    .B2(_01714_),
    .X(_01783_));
 sky130_fd_sc_hd__a31o_1 _17491_ (.A1(_01745_),
    .A2(_01775_),
    .A3(_01776_),
    .B1(_01783_),
    .X(_00610_));
 sky130_fd_sc_hd__buf_2 _17492_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_01784_));
 sky130_fd_sc_hd__clkbuf_4 _17493_ (.A(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__clkbuf_4 _17494_ (.A(_01785_),
    .X(_01786_));
 sky130_fd_sc_hd__xnor2_1 _17495_ (.A(_01786_),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_01787_));
 sky130_fd_sc_hd__a21oi_1 _17496_ (.A1(_01772_),
    .A2(_01776_),
    .B1(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__a311oi_1 _17497_ (.A1(_01772_),
    .A2(_01776_),
    .A3(_01787_),
    .B1(_01788_),
    .C1(_03486_),
    .Y(_01789_));
 sky130_fd_sc_hd__xor2_1 _17498_ (.A(_04109_),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_01790_));
 sky130_fd_sc_hd__nor2_1 _17499_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_01791_));
 sky130_fd_sc_hd__and2b_1 _17500_ (.A_N(_01781_),
    .B(_01780_),
    .X(_01792_));
 sky130_fd_sc_hd__a21o_1 _17501_ (.A1(_01791_),
    .A2(_01779_),
    .B1(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__xnor2_1 _17502_ (.A(_01790_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__xnor2_1 _17503_ (.A(_01777_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21o_1 _17504_ (.A1(_01714_),
    .A2(_01795_),
    .B1(_08448_),
    .X(_01796_));
 sky130_fd_sc_hd__o22a_1 _17505_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(_00013_),
    .B1(_01789_),
    .B2(_01796_),
    .X(_00611_));
 sky130_fd_sc_hd__o21ai_1 _17506_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(_01784_),
    .Y(_01797_));
 sky130_fd_sc_hd__o21bai_1 _17507_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1_N(_01776_),
    .Y(_01798_));
 sky130_fd_sc_hd__and2_1 _17508_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_01799_));
 sky130_fd_sc_hd__nor2_1 _17509_ (.A(_01784_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_01800_));
 sky130_fd_sc_hd__a211o_1 _17510_ (.A1(_01797_),
    .A2(_01798_),
    .B1(_01799_),
    .C1(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__o211ai_1 _17511_ (.A1(_01799_),
    .A2(_01800_),
    .B1(_01797_),
    .C1(_01798_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand2_1 _17512_ (.A(_01790_),
    .B(_01793_),
    .Y(_01803_));
 sky130_fd_sc_hd__o21ai_1 _17513_ (.A1(_01792_),
    .A2(_01790_),
    .B1(_01777_),
    .Y(_01804_));
 sky130_fd_sc_hd__or2_1 _17514_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_01805_));
 sky130_fd_sc_hd__nand2_1 _17515_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _17516_ (.A(_01805_),
    .B(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__or3_1 _17517_ (.A(_04109_),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .C(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__o21ai_1 _17518_ (.A1(_04109_),
    .A2(\rbzero.debug_overlay.vplaneY[-6] ),
    .B1(_01807_),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_1 _17519_ (.A(_01808_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__a21o_1 _17520_ (.A1(_01803_),
    .A2(_01804_),
    .B1(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__nand3_1 _17521_ (.A(_01803_),
    .B(_01810_),
    .C(_01804_),
    .Y(_01812_));
 sky130_fd_sc_hd__a32o_1 _17522_ (.A1(_01722_),
    .A2(_01811_),
    .A3(_01812_),
    .B1(_08448_),
    .B2(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_01813_));
 sky130_fd_sc_hd__a31o_1 _17523_ (.A1(_01745_),
    .A2(_01801_),
    .A3(_01802_),
    .B1(_01813_),
    .X(_00612_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(_01786_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_01814_));
 sky130_fd_sc_hd__xor2_1 _17525_ (.A(_01784_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_01815_));
 sky130_fd_sc_hd__a21oi_1 _17526_ (.A1(_01814_),
    .A2(_01801_),
    .B1(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__a31o_1 _17527_ (.A1(_01814_),
    .A2(_01801_),
    .A3(_01815_),
    .B1(_03339_),
    .X(_01817_));
 sky130_fd_sc_hd__or2_1 _17528_ (.A(_01757_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_01818_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_01757_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _17530_ (.A(_01818_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__a21o_1 _17531_ (.A1(_01808_),
    .A2(_01811_),
    .B1(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__nand3_1 _17532_ (.A(_01808_),
    .B(_01811_),
    .C(_01820_),
    .Y(_01822_));
 sky130_fd_sc_hd__and2_1 _17533_ (.A(_01821_),
    .B(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__xnor2_1 _17534_ (.A(_01805_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__o22a_1 _17535_ (.A1(_01816_),
    .A2(_01817_),
    .B1(_01824_),
    .B2(_03484_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _17536_ (.A0(\rbzero.wall_tracer.rayAddendY[4] ),
    .A1(_01825_),
    .S(_03509_),
    .X(_01826_));
 sky130_fd_sc_hd__clkbuf_1 _17537_ (.A(_01826_),
    .X(_00613_));
 sky130_fd_sc_hd__nand2_1 _17538_ (.A(_01784_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_01827_));
 sky130_fd_sc_hd__or2_1 _17539_ (.A(_01784_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_01828_));
 sky130_fd_sc_hd__nand2_1 _17540_ (.A(_01827_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__or2b_1 _17541_ (.A(_01801_),
    .B_N(_01815_),
    .X(_01830_));
 sky130_fd_sc_hd__o21ai_1 _17542_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_01786_),
    .Y(_01831_));
 sky130_fd_sc_hd__nand3_1 _17543_ (.A(_01829_),
    .B(_01830_),
    .C(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__a21o_1 _17544_ (.A1(_01830_),
    .A2(_01831_),
    .B1(_01829_),
    .X(_01833_));
 sky130_fd_sc_hd__nor2_1 _17545_ (.A(_01784_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .Y(_01834_));
 sky130_fd_sc_hd__and2_1 _17546_ (.A(_01784_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_01835_));
 sky130_fd_sc_hd__o21a_1 _17547_ (.A1(_01834_),
    .A2(_01835_),
    .B1(_01818_),
    .X(_01836_));
 sky130_fd_sc_hd__nor3_1 _17548_ (.A(_01818_),
    .B(_01834_),
    .C(_01835_),
    .Y(_01837_));
 sky130_fd_sc_hd__nor2_1 _17549_ (.A(_01836_),
    .B(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__a22o_1 _17550_ (.A1(_01811_),
    .A2(_01820_),
    .B1(_01821_),
    .B2(_01805_),
    .X(_01839_));
 sky130_fd_sc_hd__xnor2_1 _17551_ (.A(_01838_),
    .B(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__a22o_1 _17552_ (.A1(\rbzero.wall_tracer.rayAddendY[5] ),
    .A2(_08447_),
    .B1(_01840_),
    .B2(_01714_),
    .X(_01841_));
 sky130_fd_sc_hd__a31o_1 _17553_ (.A1(_01745_),
    .A2(_01832_),
    .A3(_01833_),
    .B1(_01841_),
    .X(_00614_));
 sky130_fd_sc_hd__xnor2_1 _17554_ (.A(_01785_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_01842_));
 sky130_fd_sc_hd__nand3_1 _17555_ (.A(_01827_),
    .B(_01833_),
    .C(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21o_1 _17556_ (.A1(_01827_),
    .A2(_01833_),
    .B1(_01842_),
    .X(_01844_));
 sky130_fd_sc_hd__or2_1 _17557_ (.A(_01784_),
    .B(_04109_),
    .X(_01845_));
 sky130_fd_sc_hd__nand2_1 _17558_ (.A(_01785_),
    .B(_04109_),
    .Y(_01846_));
 sky130_fd_sc_hd__a21o_1 _17559_ (.A1(_01845_),
    .A2(_01846_),
    .B1(_01834_),
    .X(_01847_));
 sky130_fd_sc_hd__nand2_1 _17560_ (.A(_04109_),
    .B(_01834_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _17561_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__o21bai_1 _17562_ (.A1(_01836_),
    .A2(_01839_),
    .B1_N(_01837_),
    .Y(_01850_));
 sky130_fd_sc_hd__xnor2_1 _17563_ (.A(_01849_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__a22o_1 _17564_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(_08447_),
    .B1(_01851_),
    .B2(_01714_),
    .X(_01852_));
 sky130_fd_sc_hd__a31o_1 _17565_ (.A1(_08458_),
    .A2(_01843_),
    .A3(_01844_),
    .B1(_01852_),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_1 _17566_ (.A(_01785_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_01853_));
 sky130_fd_sc_hd__or2_1 _17567_ (.A(_01785_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_01854_));
 sky130_fd_sc_hd__nor3_1 _17568_ (.A(_01829_),
    .B(_01830_),
    .C(_01842_),
    .Y(_01855_));
 sky130_fd_sc_hd__o41a_1 _17569_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .A3(\rbzero.wall_tracer.rayAddendY[4] ),
    .A4(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_01785_),
    .X(_01856_));
 sky130_fd_sc_hd__a211o_1 _17570_ (.A1(_01853_),
    .A2(_01854_),
    .B1(_01855_),
    .C1(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__o211ai_2 _17571_ (.A1(_01855_),
    .A2(_01856_),
    .B1(_01853_),
    .C1(_01854_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _17572_ (.A(_01785_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .Y(_01859_));
 sky130_fd_sc_hd__and2_1 _17573_ (.A(_01784_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_01860_));
 sky130_fd_sc_hd__o21ai_1 _17574_ (.A1(_01859_),
    .A2(_01860_),
    .B1(_01845_),
    .Y(_01861_));
 sky130_fd_sc_hd__or3_1 _17575_ (.A(_01845_),
    .B(_01859_),
    .C(_01860_),
    .X(_01862_));
 sky130_fd_sc_hd__nand2_1 _17576_ (.A(_01861_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__a21boi_1 _17577_ (.A1(_01847_),
    .A2(_01850_),
    .B1_N(_01848_),
    .Y(_01864_));
 sky130_fd_sc_hd__xor2_1 _17578_ (.A(_01863_),
    .B(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__a22o_1 _17579_ (.A1(\rbzero.wall_tracer.rayAddendY[7] ),
    .A2(_08447_),
    .B1(_01865_),
    .B2(_01714_),
    .X(_01866_));
 sky130_fd_sc_hd__a31o_1 _17580_ (.A1(_08458_),
    .A2(_01857_),
    .A3(_01858_),
    .B1(_01866_),
    .X(_00616_));
 sky130_fd_sc_hd__xnor2_1 _17581_ (.A(_01785_),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_01867_));
 sky130_fd_sc_hd__a21oi_1 _17582_ (.A1(_01853_),
    .A2(_01858_),
    .B1(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__a31o_1 _17583_ (.A1(_01853_),
    .A2(_01858_),
    .A3(_01867_),
    .B1(_03339_),
    .X(_01869_));
 sky130_fd_sc_hd__or2_1 _17584_ (.A(_01863_),
    .B(_01864_),
    .X(_01870_));
 sky130_fd_sc_hd__inv_2 _17585_ (.A(_01757_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21oi_1 _17586_ (.A1(_01757_),
    .A2(\rbzero.debug_overlay.vplaneY[-1] ),
    .B1(_01785_),
    .Y(_01872_));
 sky130_fd_sc_hd__a21oi_1 _17587_ (.A1(_01786_),
    .A2(_01757_),
    .B1(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__a21oi_1 _17588_ (.A1(_01871_),
    .A2(_01859_),
    .B1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__a21o_1 _17589_ (.A1(_01862_),
    .A2(_01870_),
    .B1(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__nand2_1 _17590_ (.A(_03339_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__a31o_1 _17591_ (.A1(_01862_),
    .A2(_01870_),
    .A3(_01874_),
    .B1(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__o21ai_1 _17592_ (.A1(_01868_),
    .A2(_01869_),
    .B1(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__mux2_1 _17593_ (.A0(\rbzero.wall_tracer.rayAddendY[8] ),
    .A1(_01878_),
    .S(_03509_),
    .X(_01879_));
 sky130_fd_sc_hd__clkbuf_1 _17594_ (.A(_01879_),
    .X(_00617_));
 sky130_fd_sc_hd__or2_1 _17595_ (.A(_01786_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_01880_));
 sky130_fd_sc_hd__nand2_1 _17596_ (.A(_01786_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_1 _17597_ (.A(_01880_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__o21ai_1 _17598_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(\rbzero.wall_tracer.rayAddendY[7] ),
    .B1(_01785_),
    .Y(_01883_));
 sky130_fd_sc_hd__o21ai_1 _17599_ (.A1(_01858_),
    .A2(_01867_),
    .B1(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__xnor2_1 _17600_ (.A(_01882_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__o21ba_1 _17601_ (.A1(_01786_),
    .A2(_01757_),
    .B1_N(_01875_),
    .X(_01886_));
 sky130_fd_sc_hd__a211o_1 _17602_ (.A1(_01872_),
    .A2(_01875_),
    .B1(_01886_),
    .C1(_03497_),
    .X(_01887_));
 sky130_fd_sc_hd__o221a_1 _17603_ (.A1(\rbzero.wall_tracer.rayAddendY[9] ),
    .A2(_00013_),
    .B1(_08464_),
    .B2(_01885_),
    .C1(_01887_),
    .X(_00618_));
 sky130_fd_sc_hd__o21ai_1 _17604_ (.A1(_01757_),
    .A2(_01875_),
    .B1(_03339_),
    .Y(_01888_));
 sky130_fd_sc_hd__a21bo_1 _17605_ (.A1(_01880_),
    .A2(_01884_),
    .B1_N(_01881_),
    .X(_01889_));
 sky130_fd_sc_hd__xnor2_1 _17606_ (.A(_01786_),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_01890_));
 sky130_fd_sc_hd__xnor2_1 _17607_ (.A(_01889_),
    .B(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__a2bb2o_1 _17608_ (.A1_N(_01786_),
    .A2_N(_01888_),
    .B1(_01891_),
    .B2(_03484_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _17609_ (.A0(\rbzero.wall_tracer.rayAddendY[10] ),
    .A1(_01892_),
    .S(_03509_),
    .X(_01893_));
 sky130_fd_sc_hd__clkbuf_1 _17610_ (.A(_01893_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _17611_ (.A0(\rbzero.debug_overlay.playerY[0] ),
    .A1(_03352_),
    .S(_09620_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _17612_ (.A0(_01894_),
    .A1(_03390_),
    .S(_05009_),
    .X(_01895_));
 sky130_fd_sc_hd__clkbuf_1 _17613_ (.A(_01895_),
    .X(_00620_));
 sky130_fd_sc_hd__or2_1 _17614_ (.A(_03390_),
    .B(_04934_),
    .X(_01896_));
 sky130_fd_sc_hd__nor2_1 _17615_ (.A(_03357_),
    .B(_09620_),
    .Y(_01897_));
 sky130_fd_sc_hd__a31o_1 _17616_ (.A1(_08509_),
    .A2(_04935_),
    .A3(_01896_),
    .B1(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _17617_ (.A0(_01898_),
    .A1(_03358_),
    .S(_05009_),
    .X(_01899_));
 sky130_fd_sc_hd__clkbuf_1 _17618_ (.A(_01899_),
    .X(_00621_));
 sky130_fd_sc_hd__xor2_1 _17619_ (.A(_04936_),
    .B(_04939_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _17620_ (.A0(\rbzero.debug_overlay.playerY[2] ),
    .A1(_01900_),
    .S(_09620_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _17621_ (.A0(_01901_),
    .A1(_03345_),
    .S(_05009_),
    .X(_01902_));
 sky130_fd_sc_hd__clkbuf_1 _17622_ (.A(_01902_),
    .X(_00622_));
 sky130_fd_sc_hd__inv_2 _17623_ (.A(_04933_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _17624_ (.A(_04941_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__xnor2_1 _17625_ (.A(_04940_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__mux2_1 _17626_ (.A0(\rbzero.debug_overlay.playerY[3] ),
    .A1(_01905_),
    .S(_09620_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _17627_ (.A0(_01906_),
    .A1(\rbzero.map_rom.a6 ),
    .S(_05009_),
    .X(_01907_));
 sky130_fd_sc_hd__clkbuf_1 _17628_ (.A(_01907_),
    .X(_00623_));
 sky130_fd_sc_hd__or2_1 _17629_ (.A(_04932_),
    .B(_04942_),
    .X(_01908_));
 sky130_fd_sc_hd__nor2_1 _17630_ (.A(_03341_),
    .B(_04943_),
    .Y(_01909_));
 sky130_fd_sc_hd__a22o_1 _17631_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_03341_),
    .B1(_01908_),
    .B2(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _17632_ (.A0(_01910_),
    .A1(\rbzero.map_rom.i_row[4] ),
    .S(_05009_),
    .X(_01911_));
 sky130_fd_sc_hd__clkbuf_1 _17633_ (.A(_01911_),
    .X(_00624_));
 sky130_fd_sc_hd__a21oi_1 _17634_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(_04923_),
    .B1(_04943_),
    .Y(_01912_));
 sky130_fd_sc_hd__xnor2_1 _17635_ (.A(_04931_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__mux2_1 _17636_ (.A0(\rbzero.debug_overlay.playerY[5] ),
    .A1(_01913_),
    .S(_09620_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _17637_ (.A0(_01914_),
    .A1(\rbzero.wall_tracer.mapY[5] ),
    .S(_05006_),
    .X(_01915_));
 sky130_fd_sc_hd__clkbuf_1 _17638_ (.A(_01915_),
    .X(_00625_));
 sky130_fd_sc_hd__nor2_1 _17639_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_1 _17640_ (.A(_04100_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_01917_));
 sky130_fd_sc_hd__and2b_1 _17641_ (.A_N(_01916_),
    .B(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__or2_1 _17642_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .X(_01919_));
 sky130_fd_sc_hd__nor2_1 _17643_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_01920_));
 sky130_fd_sc_hd__nand2_1 _17644_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .Y(_01921_));
 sky130_fd_sc_hd__nand2_1 _17645_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_01922_));
 sky130_fd_sc_hd__or2_1 _17646_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_01923_));
 sky130_fd_sc_hd__nand2_1 _17647_ (.A(_01922_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__o21a_1 _17648_ (.A1(_01921_),
    .A2(_01924_),
    .B1(_01922_),
    .X(_01925_));
 sky130_fd_sc_hd__nand2_1 _17649_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_01926_));
 sky130_fd_sc_hd__o21ai_1 _17650_ (.A1(_01920_),
    .A2(_01925_),
    .B1(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__nand2_1 _17651_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .Y(_01928_));
 sky130_fd_sc_hd__a21boi_1 _17652_ (.A1(_01919_),
    .A2(_01927_),
    .B1_N(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__xnor2_1 _17653_ (.A(_01918_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__mux2_1 _17654_ (.A0(\rbzero.debug_overlay.vplaneX[-9] ),
    .A1(_01930_),
    .S(_03484_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _17655_ (.A0(\rbzero.wall_tracer.rayAddendX[-5] ),
    .A1(_01931_),
    .S(_03509_),
    .X(_01932_));
 sky130_fd_sc_hd__clkbuf_1 _17656_ (.A(_01932_),
    .X(_00626_));
 sky130_fd_sc_hd__or2_1 _17657_ (.A(_04102_),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_01933_));
 sky130_fd_sc_hd__nand2_1 _17658_ (.A(_04102_),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .Y(_01934_));
 sky130_fd_sc_hd__o21ai_1 _17659_ (.A1(_01916_),
    .A2(_01929_),
    .B1(_01917_),
    .Y(_01935_));
 sky130_fd_sc_hd__and3_1 _17660_ (.A(_01933_),
    .B(_01934_),
    .C(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__a21oi_1 _17661_ (.A1(_01933_),
    .A2(_01934_),
    .B1(_01935_),
    .Y(_01937_));
 sky130_fd_sc_hd__o21ai_1 _17662_ (.A1(_01936_),
    .A2(_01937_),
    .B1(_03485_),
    .Y(_01938_));
 sky130_fd_sc_hd__or2_1 _17663_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_01939_));
 sky130_fd_sc_hd__nand2_1 _17664_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_01940_));
 sky130_fd_sc_hd__a31o_1 _17665_ (.A1(_01722_),
    .A2(_01939_),
    .A3(_01940_),
    .B1(_08452_),
    .X(_01941_));
 sky130_fd_sc_hd__a22o_1 _17666_ (.A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_08463_),
    .B1(_01938_),
    .B2(_01941_),
    .X(_00627_));
 sky130_fd_sc_hd__nor2_1 _17667_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_01942_));
 sky130_fd_sc_hd__and2_1 _17668_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .X(_01943_));
 sky130_fd_sc_hd__a21o_1 _17669_ (.A1(_04102_),
    .A2(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B1(_01935_),
    .X(_01944_));
 sky130_fd_sc_hd__o21ai_1 _17670_ (.A1(_04102_),
    .A2(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B1(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__o21ai_1 _17671_ (.A1(_01942_),
    .A2(_01943_),
    .B1(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__o311a_1 _17672_ (.A1(_01942_),
    .A2(_01943_),
    .A3(_01945_),
    .B1(_01946_),
    .C1(_03497_),
    .X(_01947_));
 sky130_fd_sc_hd__or2_1 _17673_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_01939_),
    .X(_01948_));
 sky130_fd_sc_hd__nand2_1 _17674_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_01939_),
    .Y(_01949_));
 sky130_fd_sc_hd__a31o_1 _17675_ (.A1(_01722_),
    .A2(_01948_),
    .A3(_01949_),
    .B1(_08460_),
    .X(_01950_));
 sky130_fd_sc_hd__o22a_1 _17676_ (.A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A2(_00013_),
    .B1(_01947_),
    .B2(_01950_),
    .X(_00628_));
 sky130_fd_sc_hd__nor2_1 _17677_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_01951_));
 sky130_fd_sc_hd__and2_1 _17678_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_01952_));
 sky130_fd_sc_hd__nand2_1 _17679_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_01953_));
 sky130_fd_sc_hd__o21ai_1 _17680_ (.A1(_01942_),
    .A2(_01945_),
    .B1(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__or3_1 _17681_ (.A(_01951_),
    .B(_01952_),
    .C(_01954_),
    .X(_01955_));
 sky130_fd_sc_hd__o21ai_1 _17682_ (.A1(_01951_),
    .A2(_01952_),
    .B1(_01954_),
    .Y(_01956_));
 sky130_fd_sc_hd__a21oi_1 _17683_ (.A1(_01955_),
    .A2(_01956_),
    .B1(_03486_),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _17684_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_01948_),
    .Y(_01958_));
 sky130_fd_sc_hd__or2_1 _17685_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_01948_),
    .X(_01959_));
 sky130_fd_sc_hd__a31o_1 _17686_ (.A1(_01722_),
    .A2(_01958_),
    .A3(_01959_),
    .B1(_08460_),
    .X(_01960_));
 sky130_fd_sc_hd__o22a_1 _17687_ (.A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A2(_00013_),
    .B1(_01957_),
    .B2(_01960_),
    .X(_00629_));
 sky130_fd_sc_hd__or2_1 _17688_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_01961_));
 sky130_fd_sc_hd__nand2_1 _17689_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _17690_ (.A(_01952_),
    .B(_01954_),
    .Y(_01963_));
 sky130_fd_sc_hd__nor2_1 _17691_ (.A(_01951_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand3_1 _17692_ (.A(_01961_),
    .B(_01962_),
    .C(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__a21o_1 _17693_ (.A1(_01961_),
    .A2(_01962_),
    .B1(_01964_),
    .X(_01966_));
 sky130_fd_sc_hd__inv_2 _17694_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_01967_));
 sky130_fd_sc_hd__o31a_1 _17695_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(\rbzero.debug_overlay.vplaneX[-7] ),
    .A3(\rbzero.debug_overlay.vplaneX[-8] ),
    .B1(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__xor2_1 _17696_ (.A(_04100_),
    .B(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__a22o_1 _17697_ (.A1(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A2(_08447_),
    .B1(_01969_),
    .B2(_01714_),
    .X(_01970_));
 sky130_fd_sc_hd__a31o_1 _17698_ (.A1(_08458_),
    .A2(_01965_),
    .A3(_01966_),
    .B1(_01970_),
    .X(_00630_));
 sky130_fd_sc_hd__a21bo_1 _17699_ (.A1(_01961_),
    .A2(_01964_),
    .B1_N(_01962_),
    .X(_01971_));
 sky130_fd_sc_hd__buf_2 _17700_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_01972_));
 sky130_fd_sc_hd__nor2_1 _17701_ (.A(_01972_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_01973_));
 sky130_fd_sc_hd__and2_1 _17702_ (.A(_01972_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_01974_));
 sky130_fd_sc_hd__or2_1 _17703_ (.A(_01973_),
    .B(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_01971_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__or2_1 _17705_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_01977_));
 sky130_fd_sc_hd__nand2_1 _17706_ (.A(_04102_),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _17707_ (.A(_01977_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _17708_ (.A(_04100_),
    .B(_01959_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21oi_1 _17709_ (.A1(_04100_),
    .A2(\rbzero.debug_overlay.vplaneX[-9] ),
    .B1(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__xnor2_1 _17710_ (.A(_01979_),
    .B(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__mux2_1 _17711_ (.A0(_01976_),
    .A1(_01982_),
    .S(_03339_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _17712_ (.A0(\rbzero.wall_tracer.rayAddendX[0] ),
    .A1(_01983_),
    .S(_03509_),
    .X(_01984_));
 sky130_fd_sc_hd__clkbuf_1 _17713_ (.A(_01984_),
    .X(_00631_));
 sky130_fd_sc_hd__buf_2 _17714_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_01985_));
 sky130_fd_sc_hd__nand2_1 _17715_ (.A(_01985_),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_01986_));
 sky130_fd_sc_hd__or2_1 _17716_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_01987_));
 sky130_fd_sc_hd__o21a_1 _17717_ (.A1(_01972_),
    .A2(\rbzero.wall_tracer.rayAddendX[0] ),
    .B1(_01971_),
    .X(_01988_));
 sky130_fd_sc_hd__a211o_1 _17718_ (.A1(_01986_),
    .A2(_01987_),
    .B1(_01988_),
    .C1(_01974_),
    .X(_01989_));
 sky130_fd_sc_hd__o211ai_2 _17719_ (.A1(_01974_),
    .A2(_01988_),
    .B1(_01987_),
    .C1(_01986_),
    .Y(_01990_));
 sky130_fd_sc_hd__a21oi_1 _17720_ (.A1(_04100_),
    .A2(\rbzero.debug_overlay.vplaneX[-9] ),
    .B1(_01979_),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_1 _17721_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_01992_));
 sky130_fd_sc_hd__and2_1 _17722_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_01993_));
 sky130_fd_sc_hd__nor2_1 _17723_ (.A(_01992_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__xnor2_1 _17724_ (.A(_01977_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__o21a_1 _17725_ (.A1(_01980_),
    .A2(_01991_),
    .B1(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__inv_2 _17726_ (.A(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__or3_1 _17727_ (.A(_01980_),
    .B(_01995_),
    .C(_01991_),
    .X(_01998_));
 sky130_fd_sc_hd__a32o_1 _17728_ (.A1(_01722_),
    .A2(_01997_),
    .A3(_01998_),
    .B1(_08448_),
    .B2(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_01999_));
 sky130_fd_sc_hd__a31o_1 _17729_ (.A1(_08458_),
    .A2(_01989_),
    .A3(_01990_),
    .B1(_01999_),
    .X(_00632_));
 sky130_fd_sc_hd__clkbuf_4 _17730_ (.A(_01985_),
    .X(_02000_));
 sky130_fd_sc_hd__clkbuf_4 _17731_ (.A(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__xnor2_1 _17732_ (.A(_02001_),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_02002_));
 sky130_fd_sc_hd__a21oi_1 _17733_ (.A1(_01986_),
    .A2(_01990_),
    .B1(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__a311oi_1 _17734_ (.A1(_01986_),
    .A2(_01990_),
    .A3(_02002_),
    .B1(_02003_),
    .C1(_03486_),
    .Y(_02004_));
 sky130_fd_sc_hd__xor2_1 _17735_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_02005_));
 sky130_fd_sc_hd__o31ai_1 _17736_ (.A1(_01977_),
    .A2(_01992_),
    .A3(_01993_),
    .B1(_01997_),
    .Y(_02006_));
 sky130_fd_sc_hd__xnor2_1 _17737_ (.A(_02005_),
    .B(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__xnor2_1 _17738_ (.A(_01992_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__a21o_1 _17739_ (.A1(_01714_),
    .A2(_02008_),
    .B1(_08448_),
    .X(_02009_));
 sky130_fd_sc_hd__o22a_1 _17740_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(_00013_),
    .B1(_02004_),
    .B2(_02009_),
    .X(_00633_));
 sky130_fd_sc_hd__o21ai_1 _17741_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[1] ),
    .B1(_01985_),
    .Y(_02010_));
 sky130_fd_sc_hd__o21bai_1 _17742_ (.A1(_01985_),
    .A2(\rbzero.wall_tracer.rayAddendX[2] ),
    .B1_N(_01990_),
    .Y(_02011_));
 sky130_fd_sc_hd__and2_1 _17743_ (.A(_01985_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02012_));
 sky130_fd_sc_hd__nor2_1 _17744_ (.A(_01985_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02013_));
 sky130_fd_sc_hd__a211o_1 _17745_ (.A1(_02010_),
    .A2(_02011_),
    .B1(_02012_),
    .C1(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__o211ai_1 _17746_ (.A1(_02012_),
    .A2(_02013_),
    .B1(_02010_),
    .C1(_02011_),
    .Y(_02015_));
 sky130_fd_sc_hd__or2_1 _17747_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_04100_),
    .X(_02016_));
 sky130_fd_sc_hd__nand2_1 _17748_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_04100_),
    .Y(_02017_));
 sky130_fd_sc_hd__and4bb_1 _17749_ (.A_N(\rbzero.debug_overlay.vplaneX[-2] ),
    .B_N(\rbzero.debug_overlay.vplaneX[-6] ),
    .C(_02016_),
    .D(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__a2bb2o_1 _17750_ (.A1_N(\rbzero.debug_overlay.vplaneX[-2] ),
    .A2_N(\rbzero.debug_overlay.vplaneX[-6] ),
    .B1(_02016_),
    .B2(_02017_),
    .X(_02019_));
 sky130_fd_sc_hd__and2b_1 _17751_ (.A_N(_02018_),
    .B(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__o21a_1 _17752_ (.A1(_01996_),
    .A2(_02005_),
    .B1(_01992_),
    .X(_02021_));
 sky130_fd_sc_hd__a21o_1 _17753_ (.A1(_02005_),
    .A2(_02006_),
    .B1(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__and2_1 _17754_ (.A(_02020_),
    .B(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__o21ai_1 _17755_ (.A1(_02020_),
    .A2(_02022_),
    .B1(_03340_),
    .Y(_02024_));
 sky130_fd_sc_hd__a2bb2o_1 _17756_ (.A1_N(_02023_),
    .A2_N(_02024_),
    .B1(\rbzero.wall_tracer.rayAddendX[3] ),
    .B2(_08447_),
    .X(_02025_));
 sky130_fd_sc_hd__a31o_1 _17757_ (.A1(_08458_),
    .A2(_02014_),
    .A3(_02015_),
    .B1(_02025_),
    .X(_00634_));
 sky130_fd_sc_hd__xor2_1 _17758_ (.A(_01972_),
    .B(_04102_),
    .X(_02026_));
 sky130_fd_sc_hd__o21a_1 _17759_ (.A1(_02018_),
    .A2(_02023_),
    .B1(_02026_),
    .X(_02027_));
 sky130_fd_sc_hd__nor3_1 _17760_ (.A(_02018_),
    .B(_02023_),
    .C(_02026_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _17761_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_04100_),
    .Y(_02029_));
 sky130_fd_sc_hd__o21ai_1 _17762_ (.A1(_02027_),
    .A2(_02028_),
    .B1(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__o31a_1 _17763_ (.A1(_02029_),
    .A2(_02027_),
    .A3(_02028_),
    .B1(_03339_),
    .X(_02031_));
 sky130_fd_sc_hd__xor2_1 _17764_ (.A(_01985_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_02032_));
 sky130_fd_sc_hd__or2b_1 _17765_ (.A(_02012_),
    .B_N(_02014_),
    .X(_02033_));
 sky130_fd_sc_hd__xor2_1 _17766_ (.A(_02032_),
    .B(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__o2bb2a_1 _17767_ (.A1_N(_02030_),
    .A2_N(_02031_),
    .B1(_03339_),
    .B2(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _17768_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02035_),
    .S(_03509_),
    .X(_02036_));
 sky130_fd_sc_hd__clkbuf_1 _17769_ (.A(_02036_),
    .X(_00635_));
 sky130_fd_sc_hd__or2b_1 _17770_ (.A(_02014_),
    .B_N(_02032_),
    .X(_02037_));
 sky130_fd_sc_hd__o21ai_1 _17771_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02001_),
    .Y(_02038_));
 sky130_fd_sc_hd__xnor2_1 _17772_ (.A(_02000_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02039_));
 sky130_fd_sc_hd__a21oi_1 _17773_ (.A1(_02037_),
    .A2(_02038_),
    .B1(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__a31o_1 _17774_ (.A1(_02039_),
    .A2(_02037_),
    .A3(_02038_),
    .B1(_08464_),
    .X(_02041_));
 sky130_fd_sc_hd__nor2_1 _17775_ (.A(_01985_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .Y(_02042_));
 sky130_fd_sc_hd__and2_1 _17776_ (.A(_01985_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_02043_));
 sky130_fd_sc_hd__o22a_1 _17777_ (.A1(_01972_),
    .A2(_04102_),
    .B1(_02042_),
    .B2(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__nor4_1 _17778_ (.A(_01972_),
    .B(_04102_),
    .C(_02042_),
    .D(_02043_),
    .Y(_02045_));
 sky130_fd_sc_hd__nor2_1 _17779_ (.A(_02044_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__o22a_1 _17780_ (.A1(_02023_),
    .A2(_02026_),
    .B1(_02027_),
    .B2(_02029_),
    .X(_02047_));
 sky130_fd_sc_hd__xnor2_1 _17781_ (.A(_02046_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__o2bb2a_1 _17782_ (.A1_N(\rbzero.wall_tracer.rayAddendX[5] ),
    .A2_N(_08460_),
    .B1(_02048_),
    .B2(_03497_),
    .X(_02049_));
 sky130_fd_sc_hd__o21ai_1 _17783_ (.A1(_02040_),
    .A2(_02041_),
    .B1(_02049_),
    .Y(_00636_));
 sky130_fd_sc_hd__xor2_1 _17784_ (.A(_02000_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_02050_));
 sky130_fd_sc_hd__a21o_1 _17785_ (.A1(_02001_),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .B1(_02040_),
    .X(_02051_));
 sky130_fd_sc_hd__nand2_1 _17786_ (.A(_02050_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__or2_1 _17787_ (.A(_02050_),
    .B(_02051_),
    .X(_02053_));
 sky130_fd_sc_hd__or2_1 _17788_ (.A(_01985_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_02054_));
 sky130_fd_sc_hd__nand2_1 _17789_ (.A(_02000_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .Y(_02055_));
 sky130_fd_sc_hd__a21o_1 _17790_ (.A1(_02054_),
    .A2(_02055_),
    .B1(_02042_),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _17791_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(_02042_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_1 _17792_ (.A(_02056_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__a21o_1 _17793_ (.A1(_02046_),
    .A2(_02047_),
    .B1(_02045_),
    .X(_02059_));
 sky130_fd_sc_hd__xnor2_1 _17794_ (.A(_02058_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__a22o_1 _17795_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(_08447_),
    .B1(_02060_),
    .B2(_01722_),
    .X(_02061_));
 sky130_fd_sc_hd__a31o_1 _17796_ (.A1(_08458_),
    .A2(_02052_),
    .A3(_02053_),
    .B1(_02061_),
    .X(_00637_));
 sky130_fd_sc_hd__nand2_1 _17797_ (.A(_02000_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_02062_));
 sky130_fd_sc_hd__or2_1 _17798_ (.A(_02000_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02063_));
 sky130_fd_sc_hd__nor3b_1 _17799_ (.A(_02039_),
    .B(_02037_),
    .C_N(_02050_),
    .Y(_02064_));
 sky130_fd_sc_hd__o41a_1 _17800_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .A3(\rbzero.wall_tracer.rayAddendX[4] ),
    .A4(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02000_),
    .X(_02065_));
 sky130_fd_sc_hd__a211o_1 _17801_ (.A1(_02062_),
    .A2(_02063_),
    .B1(_02064_),
    .C1(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__o211ai_2 _17802_ (.A1(_02064_),
    .A2(_02065_),
    .B1(_02062_),
    .C1(_02063_),
    .Y(_02067_));
 sky130_fd_sc_hd__inv_2 _17803_ (.A(_02057_),
    .Y(_02068_));
 sky130_fd_sc_hd__and3_1 _17804_ (.A(_02056_),
    .B(_02057_),
    .C(_02059_),
    .X(_02069_));
 sky130_fd_sc_hd__nor2_1 _17805_ (.A(_02000_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .Y(_02070_));
 sky130_fd_sc_hd__and2_1 _17806_ (.A(_02000_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_02071_));
 sky130_fd_sc_hd__o21ai_1 _17807_ (.A1(_02070_),
    .A2(_02071_),
    .B1(_02054_),
    .Y(_02072_));
 sky130_fd_sc_hd__or3_1 _17808_ (.A(_02054_),
    .B(_02070_),
    .C(_02071_),
    .X(_02073_));
 sky130_fd_sc_hd__o211ai_2 _17809_ (.A1(_02068_),
    .A2(_02069_),
    .B1(_02072_),
    .C1(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__a211o_1 _17810_ (.A1(_02072_),
    .A2(_02073_),
    .B1(_02068_),
    .C1(_02069_),
    .X(_02075_));
 sky130_fd_sc_hd__a32o_1 _17811_ (.A1(_03340_),
    .A2(_02074_),
    .A3(_02075_),
    .B1(_08448_),
    .B2(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02076_));
 sky130_fd_sc_hd__a31o_1 _17812_ (.A1(_08458_),
    .A2(_02066_),
    .A3(_02067_),
    .B1(_02076_),
    .X(_00638_));
 sky130_fd_sc_hd__xnor2_1 _17813_ (.A(_02000_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_02077_));
 sky130_fd_sc_hd__a21oi_1 _17814_ (.A1(_02062_),
    .A2(_02067_),
    .B1(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__a31o_1 _17815_ (.A1(_02062_),
    .A2(_02067_),
    .A3(_02077_),
    .B1(_03340_),
    .X(_02079_));
 sky130_fd_sc_hd__nor2_1 _17816_ (.A(_02078_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__inv_2 _17817_ (.A(_01972_),
    .Y(_02081_));
 sky130_fd_sc_hd__a21oi_1 _17818_ (.A1(_01972_),
    .A2(\rbzero.debug_overlay.vplaneX[-1] ),
    .B1(_02001_),
    .Y(_02082_));
 sky130_fd_sc_hd__a21oi_1 _17819_ (.A1(_02001_),
    .A2(_01972_),
    .B1(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__a21oi_1 _17820_ (.A1(_02081_),
    .A2(_02070_),
    .B1(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__a21o_1 _17821_ (.A1(_02073_),
    .A2(_02074_),
    .B1(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__nand3_1 _17822_ (.A(_02073_),
    .B(_02074_),
    .C(_02084_),
    .Y(_02086_));
 sky130_fd_sc_hd__a31o_1 _17823_ (.A1(_01722_),
    .A2(_02085_),
    .A3(_02086_),
    .B1(_08460_),
    .X(_02087_));
 sky130_fd_sc_hd__o22a_1 _17824_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(_00013_),
    .B1(_02080_),
    .B2(_02087_),
    .X(_00639_));
 sky130_fd_sc_hd__or2_1 _17825_ (.A(_02001_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_02088_));
 sky130_fd_sc_hd__nand2_1 _17826_ (.A(_02001_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_1 _17827_ (.A(_02088_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__o21ai_1 _17828_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[7] ),
    .B1(_02001_),
    .Y(_02091_));
 sky130_fd_sc_hd__o21ai_1 _17829_ (.A1(_02067_),
    .A2(_02077_),
    .B1(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__xnor2_1 _17830_ (.A(_02090_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__inv_2 _17831_ (.A(_02001_),
    .Y(_02094_));
 sky130_fd_sc_hd__a21oi_1 _17832_ (.A1(_02094_),
    .A2(_02081_),
    .B1(_02085_),
    .Y(_02095_));
 sky130_fd_sc_hd__a211o_1 _17833_ (.A1(_02082_),
    .A2(_02085_),
    .B1(_02095_),
    .C1(_03497_),
    .X(_02096_));
 sky130_fd_sc_hd__o221a_1 _17834_ (.A1(\rbzero.wall_tracer.rayAddendX[9] ),
    .A2(_03509_),
    .B1(_08464_),
    .B2(_02093_),
    .C1(_02096_),
    .X(_00640_));
 sky130_fd_sc_hd__a21bo_1 _17835_ (.A1(_02088_),
    .A2(_02092_),
    .B1_N(_02089_),
    .X(_02097_));
 sky130_fd_sc_hd__xnor2_1 _17836_ (.A(_02001_),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_02098_));
 sky130_fd_sc_hd__xnor2_1 _17837_ (.A(_02097_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__o211a_1 _17838_ (.A1(_01972_),
    .A2(_02085_),
    .B1(_03340_),
    .C1(_02094_),
    .X(_02100_));
 sky130_fd_sc_hd__o22a_1 _17839_ (.A1(_01714_),
    .A2(_02099_),
    .B1(_02100_),
    .B2(_08458_),
    .X(_02101_));
 sky130_fd_sc_hd__a21o_1 _17840_ (.A1(\rbzero.wall_tracer.rayAddendX[10] ),
    .A2(_08449_),
    .B1(_02101_),
    .X(_00641_));
 sky130_fd_sc_hd__nor2b_2 _17841_ (.A(\rbzero.spi_registers.sclk_buffer[2] ),
    .B_N(\rbzero.spi_registers.sclk_buffer[1] ),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_4 _17842_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_02981_),
    .Y(_02103_));
 sky130_fd_sc_hd__inv_2 _17843_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .Y(_02104_));
 sky130_fd_sc_hd__nand2_1 _17844_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .Y(_02105_));
 sky130_fd_sc_hd__or2_1 _17845_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(\rbzero.spi_registers.spi_counter[2] ),
    .X(_02106_));
 sky130_fd_sc_hd__clkbuf_2 _17846_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02107_));
 sky130_fd_sc_hd__o21a_1 _17847_ (.A1(_02107_),
    .A2(\rbzero.spi_registers.spi_cmd[1] ),
    .B1(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_02108_));
 sky130_fd_sc_hd__a211o_1 _17848_ (.A1(_02107_),
    .A2(\rbzero.spi_registers.spi_cmd[1] ),
    .B1(\rbzero.spi_registers.spi_cmd[3] ),
    .C1(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .Y(_02110_));
 sky130_fd_sc_hd__and3_1 _17850_ (.A(_02107_),
    .B(\rbzero.spi_registers.spi_cmd[1] ),
    .C(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__and2_1 _17851_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02112_));
 sky130_fd_sc_hd__or2_1 _17852_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02113_));
 sky130_fd_sc_hd__nor4_1 _17853_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_01660_),
    .C(_02111_),
    .D(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__a31o_1 _17854_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(_02111_),
    .A3(_02112_),
    .B1(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__nand2_1 _17855_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__o311a_1 _17856_ (.A1(_01659_),
    .A2(_02105_),
    .A3(_02106_),
    .B1(_02109_),
    .C1(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__a211oi_1 _17857_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_01659_),
    .B1(\rbzero.spi_registers.spi_counter[6] ),
    .C1(\rbzero.spi_registers.spi_counter[5] ),
    .Y(_02118_));
 sky130_fd_sc_hd__o21ai_1 _17858_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_01659_),
    .B1(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _17859_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(\rbzero.spi_registers.spi_counter[1] ),
    .Y(_02120_));
 sky130_fd_sc_hd__a31o_1 _17860_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(\rbzero.spi_registers.spi_counter[0] ),
    .A3(_02120_),
    .B1(_02109_),
    .X(_02121_));
 sky130_fd_sc_hd__or3b_2 _17861_ (.A(_02117_),
    .B(_02119_),
    .C_N(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__nand2b_2 _17862_ (.A_N(\rbzero.spi_registers.sclk_buffer[2] ),
    .B(\rbzero.spi_registers.sclk_buffer[1] ),
    .Y(_02123_));
 sky130_fd_sc_hd__a21o_1 _17863_ (.A1(_02104_),
    .A2(_02122_),
    .B1(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__o211a_1 _17864_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02102_),
    .B1(_02103_),
    .C1(_02124_),
    .X(_00642_));
 sky130_fd_sc_hd__a31o_1 _17865_ (.A1(_02113_),
    .A2(_02105_),
    .A3(_02122_),
    .B1(_02123_),
    .X(_02125_));
 sky130_fd_sc_hd__o211a_1 _17866_ (.A1(\rbzero.spi_registers.spi_counter[1] ),
    .A2(_02102_),
    .B1(_02103_),
    .C1(_02125_),
    .X(_00643_));
 sky130_fd_sc_hd__o21ai_1 _17867_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(_02112_),
    .B1(_02122_),
    .Y(_02126_));
 sky130_fd_sc_hd__a21oi_1 _17868_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(_02112_),
    .B1(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__or2_1 _17869_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(_02102_),
    .X(_02128_));
 sky130_fd_sc_hd__o211a_1 _17870_ (.A1(_02123_),
    .A2(_02127_),
    .B1(_02128_),
    .C1(_02103_),
    .X(_00644_));
 sky130_fd_sc_hd__and3_1 _17871_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(\rbzero.spi_registers.spi_counter[2] ),
    .C(_02112_),
    .X(_02129_));
 sky130_fd_sc_hd__inv_2 _17872_ (.A(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__a31o_1 _17873_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(\rbzero.spi_registers.spi_counter[1] ),
    .A3(\rbzero.spi_registers.spi_counter[0] ),
    .B1(\rbzero.spi_registers.spi_counter[3] ),
    .X(_02131_));
 sky130_fd_sc_hd__a31o_1 _17874_ (.A1(_02122_),
    .A2(_02130_),
    .A3(_02131_),
    .B1(_02123_),
    .X(_02132_));
 sky130_fd_sc_hd__o211a_1 _17875_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(_02102_),
    .B1(_02103_),
    .C1(_02132_),
    .X(_00645_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02129_),
    .Y(_02133_));
 sky130_fd_sc_hd__or2_1 _17877_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02129_),
    .X(_02134_));
 sky130_fd_sc_hd__a31o_1 _17878_ (.A1(_02122_),
    .A2(_02133_),
    .A3(_02134_),
    .B1(_02123_),
    .X(_02135_));
 sky130_fd_sc_hd__o211a_1 _17879_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_02102_),
    .B1(_02103_),
    .C1(_02135_),
    .X(_00646_));
 sky130_fd_sc_hd__nor2_1 _17880_ (.A(_02123_),
    .B(_02133_),
    .Y(_02136_));
 sky130_fd_sc_hd__and2_1 _17881_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__or2_1 _17882_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(_02136_),
    .X(_02138_));
 sky130_fd_sc_hd__and3b_1 _17883_ (.A_N(_02137_),
    .B(_02103_),
    .C(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__clkbuf_1 _17884_ (.A(_02139_),
    .X(_00647_));
 sky130_fd_sc_hd__o21ai_1 _17885_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02137_),
    .B1(_02103_),
    .Y(_02140_));
 sky130_fd_sc_hd__a21oi_1 _17886_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02137_),
    .B1(_02140_),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _17887_ (.A(\rbzero.pov.spi_done ),
    .B(_02907_),
    .Y(_02141_));
 sky130_fd_sc_hd__clkbuf_4 _17888_ (.A(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__clkbuf_4 _17889_ (.A(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _17890_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.ready_buffer[0] ),
    .S(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__clkbuf_1 _17891_ (.A(_02144_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _17892_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.ready_buffer[1] ),
    .S(_02143_),
    .X(_02145_));
 sky130_fd_sc_hd__clkbuf_1 _17893_ (.A(_02145_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _17894_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.ready_buffer[2] ),
    .S(_02143_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_1 _17895_ (.A(_02146_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _17896_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.ready_buffer[3] ),
    .S(_02143_),
    .X(_02147_));
 sky130_fd_sc_hd__clkbuf_1 _17897_ (.A(_02147_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _17898_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.ready_buffer[4] ),
    .S(_02143_),
    .X(_02148_));
 sky130_fd_sc_hd__clkbuf_1 _17899_ (.A(_02148_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _17900_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.ready_buffer[5] ),
    .S(_02143_),
    .X(_02149_));
 sky130_fd_sc_hd__clkbuf_1 _17901_ (.A(_02149_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _17902_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.ready_buffer[6] ),
    .S(_02143_),
    .X(_02150_));
 sky130_fd_sc_hd__clkbuf_1 _17903_ (.A(_02150_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _17904_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.ready_buffer[7] ),
    .S(_02143_),
    .X(_02151_));
 sky130_fd_sc_hd__clkbuf_1 _17905_ (.A(_02151_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _17906_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.ready_buffer[8] ),
    .S(_02143_),
    .X(_02152_));
 sky130_fd_sc_hd__clkbuf_1 _17907_ (.A(_02152_),
    .X(_00657_));
 sky130_fd_sc_hd__clkbuf_4 _17908_ (.A(_02142_),
    .X(_02153_));
 sky130_fd_sc_hd__mux2_1 _17909_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.ready_buffer[9] ),
    .S(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__clkbuf_1 _17910_ (.A(_02154_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _17911_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.ready_buffer[10] ),
    .S(_02153_),
    .X(_02155_));
 sky130_fd_sc_hd__clkbuf_1 _17912_ (.A(_02155_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _17913_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.ready_buffer[11] ),
    .S(_02153_),
    .X(_02156_));
 sky130_fd_sc_hd__clkbuf_1 _17914_ (.A(_02156_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _17915_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.ready_buffer[12] ),
    .S(_02153_),
    .X(_02157_));
 sky130_fd_sc_hd__clkbuf_1 _17916_ (.A(_02157_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _17917_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.ready_buffer[13] ),
    .S(_02153_),
    .X(_02158_));
 sky130_fd_sc_hd__clkbuf_1 _17918_ (.A(_02158_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _17919_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.ready_buffer[14] ),
    .S(_02153_),
    .X(_02159_));
 sky130_fd_sc_hd__clkbuf_1 _17920_ (.A(_02159_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _17921_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.ready_buffer[15] ),
    .S(_02153_),
    .X(_02160_));
 sky130_fd_sc_hd__clkbuf_1 _17922_ (.A(_02160_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _17923_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.ready_buffer[16] ),
    .S(_02153_),
    .X(_02161_));
 sky130_fd_sc_hd__clkbuf_1 _17924_ (.A(_02161_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _17925_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.ready_buffer[17] ),
    .S(_02153_),
    .X(_02162_));
 sky130_fd_sc_hd__clkbuf_1 _17926_ (.A(_02162_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _17927_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.ready_buffer[18] ),
    .S(_02153_),
    .X(_02163_));
 sky130_fd_sc_hd__clkbuf_1 _17928_ (.A(_02163_),
    .X(_00667_));
 sky130_fd_sc_hd__buf_4 _17929_ (.A(_02142_),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _17930_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.ready_buffer[19] ),
    .S(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__clkbuf_1 _17931_ (.A(_02165_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _17932_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.ready_buffer[20] ),
    .S(_02164_),
    .X(_02166_));
 sky130_fd_sc_hd__clkbuf_1 _17933_ (.A(_02166_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _17934_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.ready_buffer[21] ),
    .S(_02164_),
    .X(_02167_));
 sky130_fd_sc_hd__clkbuf_1 _17935_ (.A(_02167_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _17936_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.ready_buffer[22] ),
    .S(_02164_),
    .X(_02168_));
 sky130_fd_sc_hd__clkbuf_1 _17937_ (.A(_02168_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _17938_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.ready_buffer[23] ),
    .S(_02164_),
    .X(_02169_));
 sky130_fd_sc_hd__clkbuf_1 _17939_ (.A(_02169_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _17940_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.ready_buffer[24] ),
    .S(_02164_),
    .X(_02170_));
 sky130_fd_sc_hd__clkbuf_1 _17941_ (.A(_02170_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _17942_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.ready_buffer[25] ),
    .S(_02164_),
    .X(_02171_));
 sky130_fd_sc_hd__clkbuf_1 _17943_ (.A(_02171_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _17944_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.ready_buffer[26] ),
    .S(_02164_),
    .X(_02172_));
 sky130_fd_sc_hd__clkbuf_1 _17945_ (.A(_02172_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _17946_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.ready_buffer[27] ),
    .S(_02164_),
    .X(_02173_));
 sky130_fd_sc_hd__clkbuf_1 _17947_ (.A(_02173_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _17948_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.ready_buffer[28] ),
    .S(_02164_),
    .X(_02174_));
 sky130_fd_sc_hd__clkbuf_1 _17949_ (.A(_02174_),
    .X(_00677_));
 sky130_fd_sc_hd__clkbuf_4 _17950_ (.A(_02142_),
    .X(_02175_));
 sky130_fd_sc_hd__mux2_1 _17951_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.ready_buffer[29] ),
    .S(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__clkbuf_1 _17952_ (.A(_02176_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _17953_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.ready_buffer[30] ),
    .S(_02175_),
    .X(_02177_));
 sky130_fd_sc_hd__clkbuf_1 _17954_ (.A(_02177_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _17955_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.ready_buffer[31] ),
    .S(_02175_),
    .X(_02178_));
 sky130_fd_sc_hd__clkbuf_1 _17956_ (.A(_02178_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _17957_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.ready_buffer[32] ),
    .S(_02175_),
    .X(_02179_));
 sky130_fd_sc_hd__clkbuf_1 _17958_ (.A(_02179_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _17959_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.ready_buffer[33] ),
    .S(_02175_),
    .X(_02180_));
 sky130_fd_sc_hd__clkbuf_1 _17960_ (.A(_02180_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _17961_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.ready_buffer[34] ),
    .S(_02175_),
    .X(_02181_));
 sky130_fd_sc_hd__clkbuf_1 _17962_ (.A(_02181_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _17963_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.ready_buffer[35] ),
    .S(_02175_),
    .X(_02182_));
 sky130_fd_sc_hd__clkbuf_1 _17964_ (.A(_02182_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _17965_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.ready_buffer[36] ),
    .S(_02175_),
    .X(_02183_));
 sky130_fd_sc_hd__clkbuf_1 _17966_ (.A(_02183_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _17967_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.ready_buffer[37] ),
    .S(_02175_),
    .X(_02184_));
 sky130_fd_sc_hd__clkbuf_1 _17968_ (.A(_02184_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _17969_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.ready_buffer[38] ),
    .S(_02175_),
    .X(_02185_));
 sky130_fd_sc_hd__clkbuf_1 _17970_ (.A(_02185_),
    .X(_00687_));
 sky130_fd_sc_hd__clkbuf_4 _17971_ (.A(_02142_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _17972_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.ready_buffer[39] ),
    .S(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__clkbuf_1 _17973_ (.A(_02187_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _17974_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.ready_buffer[40] ),
    .S(_02186_),
    .X(_02188_));
 sky130_fd_sc_hd__clkbuf_1 _17975_ (.A(_02188_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _17976_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.ready_buffer[41] ),
    .S(_02186_),
    .X(_02189_));
 sky130_fd_sc_hd__clkbuf_1 _17977_ (.A(_02189_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _17978_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.ready_buffer[42] ),
    .S(_02186_),
    .X(_02190_));
 sky130_fd_sc_hd__clkbuf_1 _17979_ (.A(_02190_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _17980_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.ready_buffer[43] ),
    .S(_02186_),
    .X(_02191_));
 sky130_fd_sc_hd__clkbuf_1 _17981_ (.A(_02191_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _17982_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_02186_),
    .X(_02192_));
 sky130_fd_sc_hd__clkbuf_1 _17983_ (.A(_02192_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _17984_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.ready_buffer[45] ),
    .S(_02186_),
    .X(_02193_));
 sky130_fd_sc_hd__clkbuf_1 _17985_ (.A(_02193_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _17986_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.ready_buffer[46] ),
    .S(_02186_),
    .X(_02194_));
 sky130_fd_sc_hd__clkbuf_1 _17987_ (.A(_02194_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _17988_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.ready_buffer[47] ),
    .S(_02186_),
    .X(_02195_));
 sky130_fd_sc_hd__clkbuf_1 _17989_ (.A(_02195_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _17990_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.ready_buffer[48] ),
    .S(_02186_),
    .X(_02196_));
 sky130_fd_sc_hd__clkbuf_1 _17991_ (.A(_02196_),
    .X(_00697_));
 sky130_fd_sc_hd__clkbuf_4 _17992_ (.A(_02141_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _17993_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.ready_buffer[49] ),
    .S(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__clkbuf_1 _17994_ (.A(_02198_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _17995_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.ready_buffer[50] ),
    .S(_02197_),
    .X(_02199_));
 sky130_fd_sc_hd__clkbuf_1 _17996_ (.A(_02199_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _17997_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.ready_buffer[51] ),
    .S(_02197_),
    .X(_02200_));
 sky130_fd_sc_hd__clkbuf_1 _17998_ (.A(_02200_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _17999_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.ready_buffer[52] ),
    .S(_02197_),
    .X(_02201_));
 sky130_fd_sc_hd__clkbuf_1 _18000_ (.A(_02201_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _18001_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.ready_buffer[53] ),
    .S(_02197_),
    .X(_02202_));
 sky130_fd_sc_hd__clkbuf_1 _18002_ (.A(_02202_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _18003_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.ready_buffer[54] ),
    .S(_02197_),
    .X(_02203_));
 sky130_fd_sc_hd__clkbuf_1 _18004_ (.A(_02203_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _18005_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.ready_buffer[55] ),
    .S(_02197_),
    .X(_02204_));
 sky130_fd_sc_hd__clkbuf_1 _18006_ (.A(_02204_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _18007_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.ready_buffer[56] ),
    .S(_02197_),
    .X(_02205_));
 sky130_fd_sc_hd__clkbuf_1 _18008_ (.A(_02205_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _18009_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.ready_buffer[57] ),
    .S(_02197_),
    .X(_02206_));
 sky130_fd_sc_hd__clkbuf_1 _18010_ (.A(_02206_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _18011_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.ready_buffer[58] ),
    .S(_02197_),
    .X(_02207_));
 sky130_fd_sc_hd__clkbuf_1 _18012_ (.A(_02207_),
    .X(_00707_));
 sky130_fd_sc_hd__buf_4 _18013_ (.A(_02141_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _18014_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__clkbuf_1 _18015_ (.A(_02209_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _18016_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.ready_buffer[60] ),
    .S(_02208_),
    .X(_02210_));
 sky130_fd_sc_hd__clkbuf_1 _18017_ (.A(_02210_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _18018_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.ready_buffer[61] ),
    .S(_02208_),
    .X(_02211_));
 sky130_fd_sc_hd__clkbuf_1 _18019_ (.A(_02211_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _18020_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.ready_buffer[62] ),
    .S(_02208_),
    .X(_02212_));
 sky130_fd_sc_hd__clkbuf_1 _18021_ (.A(_02212_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _18022_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.ready_buffer[63] ),
    .S(_02208_),
    .X(_02213_));
 sky130_fd_sc_hd__clkbuf_1 _18023_ (.A(_02213_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _18024_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.ready_buffer[64] ),
    .S(_02208_),
    .X(_02214_));
 sky130_fd_sc_hd__clkbuf_1 _18025_ (.A(_02214_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _18026_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.ready_buffer[65] ),
    .S(_02208_),
    .X(_02215_));
 sky130_fd_sc_hd__clkbuf_1 _18027_ (.A(_02215_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _18028_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.ready_buffer[66] ),
    .S(_02208_),
    .X(_02216_));
 sky130_fd_sc_hd__clkbuf_1 _18029_ (.A(_02216_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _18030_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.ready_buffer[67] ),
    .S(_02208_),
    .X(_02217_));
 sky130_fd_sc_hd__clkbuf_1 _18031_ (.A(_02217_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _18032_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.ready_buffer[68] ),
    .S(_02208_),
    .X(_02218_));
 sky130_fd_sc_hd__clkbuf_1 _18033_ (.A(_02218_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _18034_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.ready_buffer[69] ),
    .S(_02142_),
    .X(_02219_));
 sky130_fd_sc_hd__clkbuf_1 _18035_ (.A(_02219_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _18036_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.ready_buffer[70] ),
    .S(_02142_),
    .X(_02220_));
 sky130_fd_sc_hd__clkbuf_1 _18037_ (.A(_02220_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _18038_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.ready_buffer[71] ),
    .S(_02142_),
    .X(_02221_));
 sky130_fd_sc_hd__clkbuf_1 _18039_ (.A(_02221_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _18040_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.ready_buffer[72] ),
    .S(_02142_),
    .X(_02222_));
 sky130_fd_sc_hd__clkbuf_1 _18041_ (.A(_02222_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _18042_ (.A0(\rbzero.pov.spi_buffer[73] ),
    .A1(\rbzero.pov.ready_buffer[73] ),
    .S(_02142_),
    .X(_02223_));
 sky130_fd_sc_hd__clkbuf_1 _18043_ (.A(_02223_),
    .X(_00722_));
 sky130_fd_sc_hd__or4_1 _18044_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(\rbzero.spi_registers.spi_counter[5] ),
    .C(\rbzero.spi_registers.spi_counter[4] ),
    .D(_02106_),
    .X(_02224_));
 sky130_fd_sc_hd__and3_1 _18045_ (.A(_02102_),
    .B(_02103_),
    .C(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__buf_2 _18046_ (.A(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__clkbuf_4 _18047_ (.A(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _18048_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__clkbuf_1 _18049_ (.A(_02228_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _18050_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02227_),
    .X(_02229_));
 sky130_fd_sc_hd__clkbuf_1 _18051_ (.A(_02229_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _18052_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02227_),
    .X(_02230_));
 sky130_fd_sc_hd__clkbuf_1 _18053_ (.A(_02230_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _18054_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02227_),
    .X(_02231_));
 sky130_fd_sc_hd__clkbuf_1 _18055_ (.A(_02231_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _18056_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02227_),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_1 _18057_ (.A(_02232_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _18058_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02227_),
    .X(_02233_));
 sky130_fd_sc_hd__clkbuf_1 _18059_ (.A(_02233_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _18060_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_02227_),
    .X(_02234_));
 sky130_fd_sc_hd__clkbuf_1 _18061_ (.A(_02234_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _18062_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02227_),
    .X(_02235_));
 sky130_fd_sc_hd__clkbuf_1 _18063_ (.A(_02235_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _18064_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02227_),
    .X(_02236_));
 sky130_fd_sc_hd__clkbuf_1 _18065_ (.A(_02236_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _18066_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02227_),
    .X(_02237_));
 sky130_fd_sc_hd__clkbuf_1 _18067_ (.A(_02237_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _18068_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02226_),
    .X(_02238_));
 sky130_fd_sc_hd__clkbuf_1 _18069_ (.A(_02238_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _18070_ (.A0(\rbzero.spi_registers.spi_buffer[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02226_),
    .X(_02239_));
 sky130_fd_sc_hd__clkbuf_1 _18071_ (.A(_02239_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _18072_ (.A0(\rbzero.spi_registers.spi_buffer[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_02226_),
    .X(_02240_));
 sky130_fd_sc_hd__clkbuf_1 _18073_ (.A(_02240_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _18074_ (.A0(\rbzero.spi_registers.spi_buffer[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_02226_),
    .X(_02241_));
 sky130_fd_sc_hd__clkbuf_1 _18075_ (.A(_02241_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _18076_ (.A0(\rbzero.spi_registers.spi_buffer[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_02226_),
    .X(_02242_));
 sky130_fd_sc_hd__clkbuf_1 _18077_ (.A(_02242_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _18078_ (.A0(\rbzero.spi_registers.spi_buffer[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_02226_),
    .X(_02243_));
 sky130_fd_sc_hd__clkbuf_1 _18079_ (.A(_02243_),
    .X(_00738_));
 sky130_fd_sc_hd__nand2_1 _18080_ (.A(_02102_),
    .B(_02103_),
    .Y(_02244_));
 sky130_fd_sc_hd__or2_2 _18081_ (.A(_02244_),
    .B(_02224_),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _18082_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(_02107_),
    .S(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__clkbuf_1 _18083_ (.A(_02246_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _18084_ (.A0(_02107_),
    .A1(\rbzero.spi_registers.spi_cmd[1] ),
    .S(_02245_),
    .X(_02247_));
 sky130_fd_sc_hd__clkbuf_1 _18085_ (.A(_02247_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _18086_ (.A0(\rbzero.spi_registers.spi_cmd[1] ),
    .A1(\rbzero.spi_registers.spi_cmd[2] ),
    .S(_02245_),
    .X(_02248_));
 sky130_fd_sc_hd__clkbuf_1 _18087_ (.A(_02248_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _18088_ (.A0(\rbzero.spi_registers.spi_cmd[2] ),
    .A1(\rbzero.spi_registers.spi_cmd[3] ),
    .S(_02245_),
    .X(_02249_));
 sky130_fd_sc_hd__clkbuf_1 _18089_ (.A(_02249_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _18090_ (.A0(net43),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_03337_),
    .X(_02250_));
 sky130_fd_sc_hd__clkbuf_1 _18091_ (.A(_02250_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _18092_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_04834_),
    .X(_02251_));
 sky130_fd_sc_hd__clkbuf_1 _18093_ (.A(_02251_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _18094_ (.A0(net42),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_03337_),
    .X(_02252_));
 sky130_fd_sc_hd__clkbuf_1 _18095_ (.A(_02252_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _18096_ (.A0(\rbzero.spi_registers.ss_buffer[1] ),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_04834_),
    .X(_02253_));
 sky130_fd_sc_hd__clkbuf_1 _18097_ (.A(_02253_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _18098_ (.A0(net44),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_03337_),
    .X(_02254_));
 sky130_fd_sc_hd__clkbuf_1 _18099_ (.A(_02254_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _18100_ (.A0(\rbzero.spi_registers.sclk_buffer[1] ),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_04834_),
    .X(_02255_));
 sky130_fd_sc_hd__clkbuf_1 _18101_ (.A(_02255_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _18102_ (.A0(\rbzero.spi_registers.sclk_buffer[2] ),
    .A1(\rbzero.spi_registers.sclk_buffer[1] ),
    .S(_04834_),
    .X(_02256_));
 sky130_fd_sc_hd__clkbuf_1 _18103_ (.A(_02256_),
    .X(_00749_));
 sky130_fd_sc_hd__inv_2 _18104_ (.A(_03906_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor3_2 _18105_ (.A(_03909_),
    .B(_02257_),
    .C(_03907_),
    .Y(_02258_));
 sky130_fd_sc_hd__and4_1 _18106_ (.A(_03517_),
    .B(\gpout0.vpos[2] ),
    .C(\gpout0.vpos[1] ),
    .D(\gpout0.vpos[0] ),
    .X(_02259_));
 sky130_fd_sc_hd__and3_1 _18107_ (.A(_03834_),
    .B(_03506_),
    .C(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__and3_4 _18108_ (.A(_03852_),
    .B(_02258_),
    .C(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__buf_4 _18109_ (.A(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__nand2_2 _18110_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__buf_2 _18111_ (.A(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_1 _18112_ (.A(_03881_),
    .B(_02263_),
    .Y(_02265_));
 sky130_fd_sc_hd__clkbuf_4 _18113_ (.A(_04828_),
    .X(_02266_));
 sky130_fd_sc_hd__o211a_1 _18114_ (.A1(\rbzero.spi_registers.new_other[6] ),
    .A2(_02264_),
    .B1(_02265_),
    .C1(_02266_),
    .X(_00750_));
 sky130_fd_sc_hd__nand2_1 _18115_ (.A(_03430_),
    .B(_02263_),
    .Y(_02267_));
 sky130_fd_sc_hd__o211a_1 _18116_ (.A1(\rbzero.spi_registers.new_other[7] ),
    .A2(_02264_),
    .B1(_02267_),
    .C1(_02266_),
    .X(_00751_));
 sky130_fd_sc_hd__and2_1 _18117_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02262_),
    .X(_02268_));
 sky130_fd_sc_hd__or2_1 _18118_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .B(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__o211a_1 _18119_ (.A1(\rbzero.spi_registers.new_other[8] ),
    .A2(_02264_),
    .B1(_02269_),
    .C1(_02266_),
    .X(_00752_));
 sky130_fd_sc_hd__nand2_1 _18120_ (.A(_03872_),
    .B(_02263_),
    .Y(_02270_));
 sky130_fd_sc_hd__o211a_1 _18121_ (.A1(\rbzero.spi_registers.new_other[9] ),
    .A2(_02264_),
    .B1(_02270_),
    .C1(_02266_),
    .X(_00753_));
 sky130_fd_sc_hd__nand2_1 _18122_ (.A(_03441_),
    .B(_02263_),
    .Y(_02271_));
 sky130_fd_sc_hd__o211a_1 _18123_ (.A1(\rbzero.spi_registers.new_other[10] ),
    .A2(_02264_),
    .B1(_02271_),
    .C1(_02266_),
    .X(_00754_));
 sky130_fd_sc_hd__nand2_1 _18124_ (.A(_03437_),
    .B(_02263_),
    .Y(_02272_));
 sky130_fd_sc_hd__o211a_1 _18125_ (.A1(\rbzero.spi_registers.new_other[0] ),
    .A2(_02264_),
    .B1(_02272_),
    .C1(_02266_),
    .X(_00755_));
 sky130_fd_sc_hd__or2_1 _18126_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(_02268_),
    .X(_02273_));
 sky130_fd_sc_hd__o211a_1 _18127_ (.A1(\rbzero.spi_registers.new_other[1] ),
    .A2(_02264_),
    .B1(_02273_),
    .C1(_02266_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _18128_ (.A(\rbzero.map_overlay.i_othery[2] ),
    .B(_02268_),
    .X(_02274_));
 sky130_fd_sc_hd__buf_2 _18129_ (.A(_04828_),
    .X(_02275_));
 sky130_fd_sc_hd__o211a_1 _18130_ (.A1(\rbzero.spi_registers.new_other[2] ),
    .A2(_02264_),
    .B1(_02274_),
    .C1(_02275_),
    .X(_00757_));
 sky130_fd_sc_hd__nand2_1 _18131_ (.A(_03873_),
    .B(_02263_),
    .Y(_02276_));
 sky130_fd_sc_hd__o211a_1 _18132_ (.A1(\rbzero.spi_registers.new_other[3] ),
    .A2(_02264_),
    .B1(_02276_),
    .C1(_02275_),
    .X(_00758_));
 sky130_fd_sc_hd__nand2_1 _18133_ (.A(_03871_),
    .B(_02263_),
    .Y(_02277_));
 sky130_fd_sc_hd__o211a_1 _18134_ (.A1(\rbzero.spi_registers.new_other[4] ),
    .A2(_02264_),
    .B1(_02277_),
    .C1(_02275_),
    .X(_00759_));
 sky130_fd_sc_hd__inv_2 _18135_ (.A(\rbzero.spi_registers.got_new_vinf ),
    .Y(_02278_));
 sky130_fd_sc_hd__and4b_1 _18136_ (.A_N(_03467_),
    .B(_03503_),
    .C(_03911_),
    .D(_03505_),
    .X(_02279_));
 sky130_fd_sc_hd__and2_1 _18137_ (.A(_02279_),
    .B(_02259_),
    .X(_02280_));
 sky130_fd_sc_hd__nand2_1 _18138_ (.A(_04503_),
    .B(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__or3b_1 _18139_ (.A(_02281_),
    .B(_03902_),
    .C_N(_02258_),
    .X(_02282_));
 sky130_fd_sc_hd__buf_2 _18140_ (.A(_02282_),
    .X(_02283_));
 sky130_fd_sc_hd__a21o_1 _18141_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_02262_),
    .B1(\rbzero.row_render.vinf ),
    .X(_02284_));
 sky130_fd_sc_hd__buf_4 _18142_ (.A(_04834_),
    .X(_02285_));
 sky130_fd_sc_hd__o311a_1 _18143_ (.A1(\rbzero.spi_registers.new_vinf ),
    .A2(_02278_),
    .A3(_02283_),
    .B1(_02284_),
    .C1(_02285_),
    .X(_00760_));
 sky130_fd_sc_hd__and2_1 _18144_ (.A(\gpout0.vpos[0] ),
    .B(_08450_),
    .X(_02286_));
 sky130_fd_sc_hd__and3_1 _18145_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__and4b_2 _18146_ (.A_N(_03901_),
    .B(_02287_),
    .C(_02258_),
    .D(_03852_),
    .X(_02288_));
 sky130_fd_sc_hd__nand2_2 _18147_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__buf_2 _18148_ (.A(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__and2_1 _18149_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_02261_),
    .X(_02291_));
 sky130_fd_sc_hd__clkbuf_2 _18150_ (.A(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__or2_1 _18151_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__o211a_1 _18152_ (.A1(\rbzero.spi_registers.new_mapd[10] ),
    .A2(_02290_),
    .B1(_02293_),
    .C1(_02275_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _18153_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .B(_02292_),
    .X(_02294_));
 sky130_fd_sc_hd__o211a_1 _18154_ (.A1(\rbzero.spi_registers.new_mapd[11] ),
    .A2(_02290_),
    .B1(_02294_),
    .C1(_02275_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _18155_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_02292_),
    .X(_02295_));
 sky130_fd_sc_hd__o211a_1 _18156_ (.A1(\rbzero.spi_registers.new_mapd[12] ),
    .A2(_02290_),
    .B1(_02295_),
    .C1(_02275_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _18157_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_02292_),
    .X(_02296_));
 sky130_fd_sc_hd__o211a_1 _18158_ (.A1(\rbzero.spi_registers.new_mapd[13] ),
    .A2(_02290_),
    .B1(_02296_),
    .C1(_02275_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _18159_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .B(_02292_),
    .X(_02297_));
 sky130_fd_sc_hd__o211a_1 _18160_ (.A1(\rbzero.spi_registers.new_mapd[14] ),
    .A2(_02290_),
    .B1(_02297_),
    .C1(_02275_),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _18161_ (.A(\rbzero.map_overlay.i_mapdx[5] ),
    .B(_02292_),
    .X(_02298_));
 sky130_fd_sc_hd__o211a_1 _18162_ (.A1(\rbzero.spi_registers.new_mapd[15] ),
    .A2(_02290_),
    .B1(_02298_),
    .C1(_02275_),
    .X(_00766_));
 sky130_fd_sc_hd__or2_1 _18163_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(_02292_),
    .X(_02299_));
 sky130_fd_sc_hd__o211a_1 _18164_ (.A1(\rbzero.spi_registers.new_mapd[4] ),
    .A2(_02290_),
    .B1(_02299_),
    .C1(_02275_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _18165_ (.A(\rbzero.map_overlay.i_mapdy[1] ),
    .B(_02292_),
    .X(_02300_));
 sky130_fd_sc_hd__clkbuf_4 _18166_ (.A(_04828_),
    .X(_02301_));
 sky130_fd_sc_hd__o211a_1 _18167_ (.A1(\rbzero.spi_registers.new_mapd[5] ),
    .A2(_02290_),
    .B1(_02300_),
    .C1(_02301_),
    .X(_00768_));
 sky130_fd_sc_hd__or2_1 _18168_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(_02292_),
    .X(_02302_));
 sky130_fd_sc_hd__o211a_1 _18169_ (.A1(\rbzero.spi_registers.new_mapd[6] ),
    .A2(_02290_),
    .B1(_02302_),
    .C1(_02301_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _18170_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(_02292_),
    .X(_02303_));
 sky130_fd_sc_hd__o211a_1 _18171_ (.A1(\rbzero.spi_registers.new_mapd[7] ),
    .A2(_02290_),
    .B1(_02303_),
    .C1(_02301_),
    .X(_00770_));
 sky130_fd_sc_hd__or2_1 _18172_ (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .B(_02291_),
    .X(_02304_));
 sky130_fd_sc_hd__o211a_1 _18173_ (.A1(\rbzero.spi_registers.new_mapd[8] ),
    .A2(_02289_),
    .B1(_02304_),
    .C1(_02301_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _18174_ (.A(\rbzero.map_overlay.i_mapdy[5] ),
    .B(_02291_),
    .X(_02305_));
 sky130_fd_sc_hd__o211a_1 _18175_ (.A1(\rbzero.spi_registers.new_mapd[9] ),
    .A2(_02289_),
    .B1(_02305_),
    .C1(_02301_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _18176_ (.A(\rbzero.mapdxw[0] ),
    .B(_02291_),
    .X(_02306_));
 sky130_fd_sc_hd__o211a_1 _18177_ (.A1(\rbzero.spi_registers.new_mapd[2] ),
    .A2(_02289_),
    .B1(_02306_),
    .C1(_02301_),
    .X(_00773_));
 sky130_fd_sc_hd__or2_1 _18178_ (.A(\rbzero.mapdxw[1] ),
    .B(_02291_),
    .X(_02307_));
 sky130_fd_sc_hd__o211a_1 _18179_ (.A1(\rbzero.spi_registers.new_mapd[3] ),
    .A2(_02289_),
    .B1(_02307_),
    .C1(_02301_),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _18180_ (.A(\rbzero.mapdyw[0] ),
    .B(_02291_),
    .X(_02308_));
 sky130_fd_sc_hd__o211a_1 _18181_ (.A1(\rbzero.spi_registers.new_mapd[0] ),
    .A2(_02289_),
    .B1(_02308_),
    .C1(_02301_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _18182_ (.A(\rbzero.mapdyw[1] ),
    .B(_02291_),
    .X(_02309_));
 sky130_fd_sc_hd__o211a_1 _18183_ (.A1(\rbzero.spi_registers.new_mapd[1] ),
    .A2(_02289_),
    .B1(_02309_),
    .C1(_02301_),
    .X(_00776_));
 sky130_fd_sc_hd__nand2_2 _18184_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02262_),
    .Y(_02310_));
 sky130_fd_sc_hd__and2_1 _18185_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02262_),
    .X(_02311_));
 sky130_fd_sc_hd__or2_1 _18186_ (.A(\rbzero.floor_leak[0] ),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__o211a_1 _18187_ (.A1(\rbzero.spi_registers.new_leak[0] ),
    .A2(_02310_),
    .B1(_02312_),
    .C1(_02301_),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _18188_ (.A(\rbzero.floor_leak[1] ),
    .B(_02311_),
    .X(_02313_));
 sky130_fd_sc_hd__buf_2 _18189_ (.A(_04828_),
    .X(_02314_));
 sky130_fd_sc_hd__o211a_1 _18190_ (.A1(\rbzero.spi_registers.new_leak[1] ),
    .A2(_02310_),
    .B1(_02313_),
    .C1(_02314_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _18191_ (.A(\rbzero.floor_leak[2] ),
    .B(_02311_),
    .X(_02315_));
 sky130_fd_sc_hd__o211a_1 _18192_ (.A1(\rbzero.spi_registers.new_leak[2] ),
    .A2(_02310_),
    .B1(_02315_),
    .C1(_02314_),
    .X(_00779_));
 sky130_fd_sc_hd__or2_1 _18193_ (.A(\rbzero.floor_leak[3] ),
    .B(_02311_),
    .X(_02316_));
 sky130_fd_sc_hd__o211a_1 _18194_ (.A1(\rbzero.spi_registers.new_leak[3] ),
    .A2(_02310_),
    .B1(_02316_),
    .C1(_02314_),
    .X(_00780_));
 sky130_fd_sc_hd__or2_1 _18195_ (.A(\rbzero.floor_leak[4] ),
    .B(_02311_),
    .X(_02317_));
 sky130_fd_sc_hd__o211a_1 _18196_ (.A1(\rbzero.spi_registers.new_leak[4] ),
    .A2(_02310_),
    .B1(_02317_),
    .C1(_02314_),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _18197_ (.A(\rbzero.floor_leak[5] ),
    .B(_02311_),
    .X(_02318_));
 sky130_fd_sc_hd__o211a_1 _18198_ (.A1(\rbzero.spi_registers.new_leak[5] ),
    .A2(_02310_),
    .B1(_02318_),
    .C1(_02314_),
    .X(_00782_));
 sky130_fd_sc_hd__buf_6 _18199_ (.A(_03337_),
    .X(_02319_));
 sky130_fd_sc_hd__and2_2 _18200_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_02261_),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _18201_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.spi_registers.new_sky[0] ),
    .S(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__or2_1 _18202_ (.A(_02319_),
    .B(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__clkbuf_1 _18203_ (.A(_02322_),
    .X(_00783_));
 sky130_fd_sc_hd__clkbuf_4 _18204_ (.A(_04827_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _18205_ (.A0(\rbzero.color_sky[1] ),
    .A1(\rbzero.spi_registers.new_sky[1] ),
    .S(_02320_),
    .X(_02324_));
 sky130_fd_sc_hd__and2_1 _18206_ (.A(_02323_),
    .B(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__clkbuf_1 _18207_ (.A(_02325_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _18208_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.spi_registers.new_sky[2] ),
    .S(_02320_),
    .X(_02326_));
 sky130_fd_sc_hd__or2_1 _18209_ (.A(_03338_),
    .B(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__clkbuf_1 _18210_ (.A(_02327_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _18211_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.spi_registers.new_sky[3] ),
    .S(_02320_),
    .X(_02328_));
 sky130_fd_sc_hd__and2_1 _18212_ (.A(_02323_),
    .B(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__clkbuf_1 _18213_ (.A(_02329_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _18214_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.spi_registers.new_sky[4] ),
    .S(_02320_),
    .X(_02330_));
 sky130_fd_sc_hd__or2_1 _18215_ (.A(_03338_),
    .B(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__clkbuf_1 _18216_ (.A(_02331_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _18217_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.spi_registers.new_sky[5] ),
    .S(_02320_),
    .X(_02332_));
 sky130_fd_sc_hd__and2_1 _18218_ (.A(_02323_),
    .B(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__clkbuf_1 _18219_ (.A(_02333_),
    .X(_00788_));
 sky130_fd_sc_hd__buf_4 _18220_ (.A(_04827_),
    .X(_02334_));
 sky130_fd_sc_hd__and2_2 _18221_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_02261_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _18222_ (.A0(\rbzero.color_floor[0] ),
    .A1(\rbzero.spi_registers.new_floor[0] ),
    .S(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__and2_1 _18223_ (.A(_02334_),
    .B(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__clkbuf_1 _18224_ (.A(_02337_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _18225_ (.A0(\rbzero.color_floor[1] ),
    .A1(\rbzero.spi_registers.new_floor[1] ),
    .S(_02335_),
    .X(_02338_));
 sky130_fd_sc_hd__or2_1 _18226_ (.A(_03338_),
    .B(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__clkbuf_1 _18227_ (.A(_02339_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _18228_ (.A0(\rbzero.color_floor[2] ),
    .A1(\rbzero.spi_registers.new_floor[2] ),
    .S(_02335_),
    .X(_02340_));
 sky130_fd_sc_hd__and2_1 _18229_ (.A(_02334_),
    .B(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__clkbuf_1 _18230_ (.A(_02341_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _18231_ (.A0(\rbzero.color_floor[3] ),
    .A1(\rbzero.spi_registers.new_floor[3] ),
    .S(_02335_),
    .X(_02342_));
 sky130_fd_sc_hd__or2_1 _18232_ (.A(_03338_),
    .B(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__clkbuf_1 _18233_ (.A(_02343_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _18234_ (.A0(\rbzero.color_floor[4] ),
    .A1(\rbzero.spi_registers.new_floor[4] ),
    .S(_02335_),
    .X(_02344_));
 sky130_fd_sc_hd__and2_1 _18235_ (.A(_02334_),
    .B(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__clkbuf_1 _18236_ (.A(_02345_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _18237_ (.A0(\rbzero.color_floor[5] ),
    .A1(\rbzero.spi_registers.new_floor[5] ),
    .S(_02335_),
    .X(_02346_));
 sky130_fd_sc_hd__or2_1 _18238_ (.A(_03338_),
    .B(_02346_),
    .X(_02347_));
 sky130_fd_sc_hd__clkbuf_1 _18239_ (.A(_02347_),
    .X(_00794_));
 sky130_fd_sc_hd__nand2_2 _18240_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02262_),
    .Y(_02348_));
 sky130_fd_sc_hd__and2_1 _18241_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02262_),
    .X(_02349_));
 sky130_fd_sc_hd__or2_1 _18242_ (.A(\rbzero.spi_registers.vshift[0] ),
    .B(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__o211a_1 _18243_ (.A1(\rbzero.spi_registers.new_vshift[0] ),
    .A2(_02348_),
    .B1(_02350_),
    .C1(_02314_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _18244_ (.A(\rbzero.spi_registers.vshift[1] ),
    .B(_02349_),
    .X(_02351_));
 sky130_fd_sc_hd__o211a_1 _18245_ (.A1(\rbzero.spi_registers.new_vshift[1] ),
    .A2(_02348_),
    .B1(_02351_),
    .C1(_02314_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _18246_ (.A(\rbzero.spi_registers.vshift[2] ),
    .B(_02349_),
    .X(_02352_));
 sky130_fd_sc_hd__o211a_1 _18247_ (.A1(\rbzero.spi_registers.new_vshift[2] ),
    .A2(_02348_),
    .B1(_02352_),
    .C1(_02314_),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _18248_ (.A(\rbzero.spi_registers.vshift[3] ),
    .B(_02349_),
    .X(_02353_));
 sky130_fd_sc_hd__o211a_1 _18249_ (.A1(\rbzero.spi_registers.new_vshift[3] ),
    .A2(_02348_),
    .B1(_02353_),
    .C1(_02314_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _18250_ (.A(\rbzero.spi_registers.vshift[4] ),
    .B(_02349_),
    .X(_02354_));
 sky130_fd_sc_hd__o211a_1 _18251_ (.A1(\rbzero.spi_registers.new_vshift[4] ),
    .A2(_02348_),
    .B1(_02354_),
    .C1(_02314_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _18252_ (.A(\rbzero.spi_registers.vshift[5] ),
    .B(_02349_),
    .X(_02355_));
 sky130_fd_sc_hd__buf_4 _18253_ (.A(_04828_),
    .X(_02356_));
 sky130_fd_sc_hd__o211a_1 _18254_ (.A1(\rbzero.spi_registers.new_vshift[5] ),
    .A2(_02348_),
    .B1(_02355_),
    .C1(_02356_),
    .X(_00800_));
 sky130_fd_sc_hd__nor2_1 _18255_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02244_),
    .Y(_02357_));
 sky130_fd_sc_hd__and4bb_1 _18256_ (.A_N(_02117_),
    .B_N(_02119_),
    .C(_02121_),
    .D(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__clkbuf_1 _18257_ (.A(_02358_),
    .X(_00801_));
 sky130_fd_sc_hd__nand2_1 _18258_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02110_),
    .Y(_02359_));
 sky130_fd_sc_hd__or4_1 _18259_ (.A(_02107_),
    .B(\rbzero.spi_registers.spi_cmd[1] ),
    .C(_02981_),
    .D(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__clkbuf_4 _18260_ (.A(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _18261_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_sky[0] ),
    .S(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__clkbuf_1 _18262_ (.A(_02362_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _18263_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_sky[1] ),
    .S(_02361_),
    .X(_02363_));
 sky130_fd_sc_hd__clkbuf_1 _18264_ (.A(_02363_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _18265_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_sky[2] ),
    .S(_02361_),
    .X(_02364_));
 sky130_fd_sc_hd__clkbuf_1 _18266_ (.A(_02364_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _18267_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_sky[3] ),
    .S(_02361_),
    .X(_02365_));
 sky130_fd_sc_hd__clkbuf_1 _18268_ (.A(_02365_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _18269_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_sky[4] ),
    .S(_02361_),
    .X(_02366_));
 sky130_fd_sc_hd__clkbuf_1 _18270_ (.A(_02366_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _18271_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_sky[5] ),
    .S(_02361_),
    .X(_02367_));
 sky130_fd_sc_hd__clkbuf_1 _18272_ (.A(_02367_),
    .X(_00807_));
 sky130_fd_sc_hd__inv_2 _18273_ (.A(_02361_),
    .Y(_02368_));
 sky130_fd_sc_hd__a31o_1 _18274_ (.A1(\rbzero.spi_registers.got_new_sky ),
    .A2(_02285_),
    .A3(_02283_),
    .B1(_02368_),
    .X(_00808_));
 sky130_fd_sc_hd__or4b_1 _18275_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(_02981_),
    .C(_02359_),
    .D_N(_02107_),
    .X(_02369_));
 sky130_fd_sc_hd__clkbuf_4 _18276_ (.A(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_1 _18277_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_floor[0] ),
    .S(_02370_),
    .X(_02371_));
 sky130_fd_sc_hd__clkbuf_1 _18278_ (.A(_02371_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _18279_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_floor[1] ),
    .S(_02370_),
    .X(_02372_));
 sky130_fd_sc_hd__clkbuf_1 _18280_ (.A(_02372_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _18281_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_floor[2] ),
    .S(_02370_),
    .X(_02373_));
 sky130_fd_sc_hd__clkbuf_1 _18282_ (.A(_02373_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _18283_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_floor[3] ),
    .S(_02370_),
    .X(_02374_));
 sky130_fd_sc_hd__clkbuf_1 _18284_ (.A(_02374_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _18285_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_floor[4] ),
    .S(_02370_),
    .X(_02375_));
 sky130_fd_sc_hd__clkbuf_1 _18286_ (.A(_02375_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _18287_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_floor[5] ),
    .S(_02370_),
    .X(_02376_));
 sky130_fd_sc_hd__clkbuf_1 _18288_ (.A(_02376_),
    .X(_00814_));
 sky130_fd_sc_hd__inv_2 _18289_ (.A(_02370_),
    .Y(_02377_));
 sky130_fd_sc_hd__a31o_1 _18290_ (.A1(\rbzero.spi_registers.got_new_floor ),
    .A2(_02323_),
    .A3(_02283_),
    .B1(_02377_),
    .X(_00815_));
 sky130_fd_sc_hd__or4_1 _18291_ (.A(_02107_),
    .B(_01658_),
    .C(_02981_),
    .D(_02359_),
    .X(_02378_));
 sky130_fd_sc_hd__clkbuf_4 _18292_ (.A(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__mux2_1 _18293_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_leak[0] ),
    .S(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__clkbuf_1 _18294_ (.A(_02380_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _18295_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_leak[1] ),
    .S(_02379_),
    .X(_02381_));
 sky130_fd_sc_hd__clkbuf_1 _18296_ (.A(_02381_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _18297_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_leak[2] ),
    .S(_02379_),
    .X(_02382_));
 sky130_fd_sc_hd__clkbuf_1 _18298_ (.A(_02382_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _18299_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_leak[3] ),
    .S(_02379_),
    .X(_02383_));
 sky130_fd_sc_hd__clkbuf_1 _18300_ (.A(_02383_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _18301_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_leak[4] ),
    .S(_02379_),
    .X(_02384_));
 sky130_fd_sc_hd__clkbuf_1 _18302_ (.A(_02384_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _18303_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_leak[5] ),
    .S(_02379_),
    .X(_02385_));
 sky130_fd_sc_hd__clkbuf_1 _18304_ (.A(_02385_),
    .X(_00821_));
 sky130_fd_sc_hd__inv_2 _18305_ (.A(_02379_),
    .Y(_02386_));
 sky130_fd_sc_hd__a31o_1 _18306_ (.A1(\rbzero.spi_registers.got_new_leak ),
    .A2(_02323_),
    .A3(_02283_),
    .B1(_02386_),
    .X(_00822_));
 sky130_fd_sc_hd__and3_1 _18307_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02907_),
    .C(_02111_),
    .X(_02387_));
 sky130_fd_sc_hd__clkbuf_4 _18308_ (.A(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _18309_ (.A0(\rbzero.spi_registers.new_other[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__clkbuf_1 _18310_ (.A(_02389_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _18311_ (.A0(\rbzero.spi_registers.new_other[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02388_),
    .X(_02390_));
 sky130_fd_sc_hd__clkbuf_1 _18312_ (.A(_02390_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _18313_ (.A0(\rbzero.spi_registers.new_other[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02388_),
    .X(_02391_));
 sky130_fd_sc_hd__clkbuf_1 _18314_ (.A(_02391_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _18315_ (.A0(\rbzero.spi_registers.new_other[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02388_),
    .X(_02392_));
 sky130_fd_sc_hd__clkbuf_1 _18316_ (.A(_02392_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _18317_ (.A0(\rbzero.spi_registers.new_other[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02388_),
    .X(_02393_));
 sky130_fd_sc_hd__clkbuf_1 _18318_ (.A(_02393_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _18319_ (.A0(\rbzero.spi_registers.new_other[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02388_),
    .X(_02394_));
 sky130_fd_sc_hd__clkbuf_1 _18320_ (.A(_02394_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _18321_ (.A0(\rbzero.spi_registers.new_other[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02388_),
    .X(_02395_));
 sky130_fd_sc_hd__clkbuf_1 _18322_ (.A(_02395_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _18323_ (.A0(\rbzero.spi_registers.new_other[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02388_),
    .X(_02396_));
 sky130_fd_sc_hd__clkbuf_1 _18324_ (.A(_02396_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _18325_ (.A0(\rbzero.spi_registers.new_other[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02388_),
    .X(_02397_));
 sky130_fd_sc_hd__clkbuf_1 _18326_ (.A(_02397_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _18327_ (.A0(\rbzero.spi_registers.new_other[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02387_),
    .X(_02398_));
 sky130_fd_sc_hd__clkbuf_1 _18328_ (.A(_02398_),
    .X(_00832_));
 sky130_fd_sc_hd__a31o_1 _18329_ (.A1(\rbzero.spi_registers.got_new_other ),
    .A2(_02323_),
    .A3(_02283_),
    .B1(_02388_),
    .X(_00833_));
 sky130_fd_sc_hd__and3b_1 _18330_ (.A_N(\rbzero.spi_registers.spi_cmd[3] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .C(\rbzero.spi_registers.spi_done ),
    .X(_02399_));
 sky130_fd_sc_hd__and4b_1 _18331_ (.A_N(_02107_),
    .B(_01658_),
    .C(_02907_),
    .D(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__clkbuf_4 _18332_ (.A(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _18333_ (.A0(\rbzero.spi_registers.new_vshift[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__clkbuf_1 _18334_ (.A(_02402_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _18335_ (.A0(\rbzero.spi_registers.new_vshift[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02401_),
    .X(_02403_));
 sky130_fd_sc_hd__clkbuf_1 _18336_ (.A(_02403_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _18337_ (.A0(\rbzero.spi_registers.new_vshift[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02401_),
    .X(_02404_));
 sky130_fd_sc_hd__clkbuf_1 _18338_ (.A(_02404_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _18339_ (.A0(\rbzero.spi_registers.new_vshift[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02401_),
    .X(_02405_));
 sky130_fd_sc_hd__clkbuf_1 _18340_ (.A(_02405_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _18341_ (.A0(\rbzero.spi_registers.new_vshift[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02401_),
    .X(_02406_));
 sky130_fd_sc_hd__clkbuf_1 _18342_ (.A(_02406_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _18343_ (.A0(\rbzero.spi_registers.new_vshift[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_02401_),
    .X(_02407_));
 sky130_fd_sc_hd__clkbuf_1 _18344_ (.A(_02407_),
    .X(_00839_));
 sky130_fd_sc_hd__a31o_1 _18345_ (.A1(\rbzero.spi_registers.got_new_vshift ),
    .A2(_02323_),
    .A3(_02283_),
    .B1(_02401_),
    .X(_00840_));
 sky130_fd_sc_hd__and4_1 _18346_ (.A(_02107_),
    .B(_01658_),
    .C(_02907_),
    .D(_02399_),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _18347_ (.A0(\rbzero.spi_registers.new_vinf ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__clkbuf_1 _18348_ (.A(_02409_),
    .X(_00841_));
 sky130_fd_sc_hd__a31o_1 _18349_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_02323_),
    .A3(_02283_),
    .B1(_02408_),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _18350_ (.A(net40),
    .B(net39),
    .X(_02410_));
 sky130_fd_sc_hd__clkbuf_4 _18351_ (.A(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__nand2_2 _18352_ (.A(_02261_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__clkbuf_4 _18353_ (.A(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__o211a_1 _18354_ (.A1(\rbzero.pov.spi_done ),
    .A2(\rbzero.pov.ready ),
    .B1(_02285_),
    .C1(_02413_),
    .X(_00843_));
 sky130_fd_sc_hd__nor2b_2 _18355_ (.A(\rbzero.pov.sclk_buffer[2] ),
    .B_N(\rbzero.pov.sclk_buffer[1] ),
    .Y(_02414_));
 sky130_fd_sc_hd__nor2_2 _18356_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(_02981_),
    .Y(_02415_));
 sky130_fd_sc_hd__o21ai_1 _18357_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_02414_),
    .B1(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__a21oi_1 _18358_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_02414_),
    .B1(_02416_),
    .Y(_00844_));
 sky130_fd_sc_hd__and3_1 _18359_ (.A(\rbzero.pov.spi_counter[1] ),
    .B(\rbzero.pov.spi_counter[0] ),
    .C(_02414_),
    .X(_02417_));
 sky130_fd_sc_hd__a21o_1 _18360_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_02414_),
    .B1(\rbzero.pov.spi_counter[1] ),
    .X(_02418_));
 sky130_fd_sc_hd__and4bb_1 _18361_ (.A_N(\rbzero.pov.spi_counter[5] ),
    .B_N(\rbzero.pov.spi_counter[4] ),
    .C(\rbzero.pov.spi_counter[3] ),
    .D(\rbzero.pov.spi_counter[6] ),
    .X(_02419_));
 sky130_fd_sc_hd__and4bb_1 _18362_ (.A_N(\rbzero.pov.spi_counter[2] ),
    .B_N(\rbzero.pov.spi_counter[1] ),
    .C(\rbzero.pov.spi_counter[0] ),
    .D(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__a21boi_1 _18363_ (.A1(_02414_),
    .A2(_02420_),
    .B1_N(_02415_),
    .Y(_02421_));
 sky130_fd_sc_hd__and3b_1 _18364_ (.A_N(_02417_),
    .B(_02418_),
    .C(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__clkbuf_1 _18365_ (.A(_02422_),
    .X(_00845_));
 sky130_fd_sc_hd__and2_1 _18366_ (.A(\rbzero.pov.spi_counter[2] ),
    .B(_02417_),
    .X(_02423_));
 sky130_fd_sc_hd__o21ai_1 _18367_ (.A1(\rbzero.pov.spi_counter[2] ),
    .A2(_02417_),
    .B1(_02415_),
    .Y(_02424_));
 sky130_fd_sc_hd__nor2_1 _18368_ (.A(_02423_),
    .B(_02424_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _18369_ (.A(\rbzero.pov.spi_counter[3] ),
    .B(_02423_),
    .Y(_02425_));
 sky130_fd_sc_hd__o211a_1 _18370_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_02423_),
    .B1(_02425_),
    .C1(_02421_),
    .X(_00847_));
 sky130_fd_sc_hd__and3_1 _18371_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[3] ),
    .C(_02423_),
    .X(_02426_));
 sky130_fd_sc_hd__a31o_1 _18372_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(\rbzero.pov.spi_counter[2] ),
    .A3(_02417_),
    .B1(\rbzero.pov.spi_counter[4] ),
    .X(_02427_));
 sky130_fd_sc_hd__and3b_1 _18373_ (.A_N(_02426_),
    .B(_02415_),
    .C(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__clkbuf_1 _18374_ (.A(_02428_),
    .X(_00848_));
 sky130_fd_sc_hd__a21boi_1 _18375_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_02426_),
    .B1_N(_02415_),
    .Y(_02429_));
 sky130_fd_sc_hd__o21a_1 _18376_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_02426_),
    .B1(_02429_),
    .X(_00849_));
 sky130_fd_sc_hd__a21o_1 _18377_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_02426_),
    .B1(\rbzero.pov.spi_counter[6] ),
    .X(_02430_));
 sky130_fd_sc_hd__nand3_1 _18378_ (.A(\rbzero.pov.spi_counter[6] ),
    .B(\rbzero.pov.spi_counter[5] ),
    .C(_02426_),
    .Y(_02431_));
 sky130_fd_sc_hd__and3_1 _18379_ (.A(_02421_),
    .B(_02430_),
    .C(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__clkbuf_1 _18380_ (.A(_02432_),
    .X(_00850_));
 sky130_fd_sc_hd__buf_1 _18381_ (.A(clknet_1_0__leaf__04486_),
    .X(_02433_));
 sky130_fd_sc_hd__buf_1 _18382_ (.A(clknet_1_1__leaf__02433_),
    .X(_02434_));
 sky130_fd_sc_hd__inv_2 _18384__28 (.A(clknet_1_1__leaf__02434_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _18385__29 (.A(clknet_1_0__leaf__02434_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _18386__30 (.A(clknet_1_0__leaf__02434_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _18387__31 (.A(clknet_1_0__leaf__02434_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _18388__32 (.A(clknet_1_0__leaf__02434_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _18389__33 (.A(clknet_1_0__leaf__02434_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _18390__34 (.A(clknet_1_1__leaf__02434_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _18391__35 (.A(clknet_1_1__leaf__02434_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _18392__36 (.A(clknet_1_1__leaf__02434_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _18394__37 (.A(clknet_1_0__leaf__02435_),
    .Y(net159));
 sky130_fd_sc_hd__buf_1 _18393_ (.A(clknet_1_1__leaf__02433_),
    .X(_02435_));
 sky130_fd_sc_hd__inv_2 _18395__38 (.A(clknet_1_0__leaf__02435_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _18396__39 (.A(clknet_1_0__leaf__02435_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _18397__40 (.A(clknet_1_0__leaf__02435_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _18398__41 (.A(clknet_1_1__leaf__02435_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _18399__42 (.A(clknet_1_1__leaf__02435_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _18400__43 (.A(clknet_1_1__leaf__02435_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _18401__44 (.A(clknet_1_1__leaf__02435_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _18402__45 (.A(clknet_1_1__leaf__02435_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _18403__46 (.A(clknet_1_0__leaf__02435_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _18405__47 (.A(clknet_1_0__leaf__02436_),
    .Y(net169));
 sky130_fd_sc_hd__buf_1 _18404_ (.A(clknet_1_1__leaf__02433_),
    .X(_02436_));
 sky130_fd_sc_hd__inv_2 _18406__48 (.A(clknet_1_0__leaf__02436_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _18407__49 (.A(clknet_1_0__leaf__02436_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _18408__50 (.A(clknet_1_0__leaf__02436_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _18409__51 (.A(clknet_1_0__leaf__02436_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _18410__52 (.A(clknet_1_1__leaf__02436_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _18411__53 (.A(clknet_1_1__leaf__02436_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _18412__54 (.A(clknet_1_1__leaf__02436_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _18413__55 (.A(clknet_1_1__leaf__02436_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _18414__56 (.A(clknet_1_1__leaf__02436_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _18416__57 (.A(clknet_1_1__leaf__02437_),
    .Y(net179));
 sky130_fd_sc_hd__buf_1 _18415_ (.A(clknet_1_1__leaf__02433_),
    .X(_02437_));
 sky130_fd_sc_hd__inv_2 _18417__58 (.A(clknet_1_1__leaf__02437_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _18418__59 (.A(clknet_1_1__leaf__02437_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _18419__60 (.A(clknet_1_1__leaf__02437_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _18420__61 (.A(clknet_1_1__leaf__02437_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _18421__62 (.A(clknet_1_1__leaf__02437_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _18422__63 (.A(clknet_1_0__leaf__02437_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _18423__64 (.A(clknet_1_0__leaf__02437_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _18424__65 (.A(clknet_1_0__leaf__02437_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _18425__66 (.A(clknet_1_0__leaf__02437_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _18427__67 (.A(clknet_1_1__leaf__02438_),
    .Y(net189));
 sky130_fd_sc_hd__buf_1 _18426_ (.A(clknet_1_0__leaf__02433_),
    .X(_02438_));
 sky130_fd_sc_hd__inv_2 _18428__68 (.A(clknet_1_1__leaf__02438_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _18429__69 (.A(clknet_1_1__leaf__02438_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _18430__70 (.A(clknet_1_0__leaf__02438_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _18431__71 (.A(clknet_1_0__leaf__02438_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _18432__72 (.A(clknet_1_0__leaf__02438_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _18433__73 (.A(clknet_1_0__leaf__02438_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _18434__74 (.A(clknet_1_0__leaf__02438_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _18435__75 (.A(clknet_1_1__leaf__02438_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _18436__76 (.A(clknet_1_1__leaf__02438_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _18438__77 (.A(clknet_1_1__leaf__02439_),
    .Y(net199));
 sky130_fd_sc_hd__buf_1 _18437_ (.A(clknet_1_0__leaf__02433_),
    .X(_02439_));
 sky130_fd_sc_hd__inv_2 _18439__78 (.A(clknet_1_1__leaf__02439_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _18440__79 (.A(clknet_1_0__leaf__02439_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _18441__80 (.A(clknet_1_0__leaf__02439_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _18442__81 (.A(clknet_1_0__leaf__02439_),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _18443__82 (.A(clknet_1_1__leaf__02439_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _18444__83 (.A(clknet_1_1__leaf__02439_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _18445__84 (.A(clknet_1_0__leaf__02439_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _18446__85 (.A(clknet_1_0__leaf__02439_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _18447__86 (.A(clknet_1_0__leaf__02439_),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _18450__87 (.A(clknet_1_0__leaf__02441_),
    .Y(net209));
 sky130_fd_sc_hd__buf_1 _18448_ (.A(clknet_1_0__leaf__04486_),
    .X(_02440_));
 sky130_fd_sc_hd__buf_1 _18449_ (.A(clknet_1_0__leaf__02440_),
    .X(_02441_));
 sky130_fd_sc_hd__inv_2 _18451__88 (.A(clknet_1_0__leaf__02441_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _18452__89 (.A(clknet_1_0__leaf__02441_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _18453__90 (.A(clknet_1_1__leaf__02441_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _18904__91 (.A(clknet_1_1__leaf__02441_),
    .Y(net213));
 sky130_fd_sc_hd__nand2_1 _18454_ (.A(_02415_),
    .B(_02414_),
    .Y(_02442_));
 sky130_fd_sc_hd__clkbuf_4 _18455_ (.A(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__clkbuf_4 _18456_ (.A(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _18457_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.spi_buffer[0] ),
    .S(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__clkbuf_1 _18458_ (.A(_02445_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _18459_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.spi_buffer[1] ),
    .S(_02444_),
    .X(_02446_));
 sky130_fd_sc_hd__clkbuf_1 _18460_ (.A(_02446_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _18461_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.spi_buffer[2] ),
    .S(_02444_),
    .X(_02447_));
 sky130_fd_sc_hd__clkbuf_1 _18462_ (.A(_02447_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _18463_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.spi_buffer[3] ),
    .S(_02444_),
    .X(_02448_));
 sky130_fd_sc_hd__clkbuf_1 _18464_ (.A(_02448_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _18465_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.spi_buffer[4] ),
    .S(_02444_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_1 _18466_ (.A(_02449_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _18467_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.spi_buffer[5] ),
    .S(_02444_),
    .X(_02450_));
 sky130_fd_sc_hd__clkbuf_1 _18468_ (.A(_02450_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _18469_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.spi_buffer[6] ),
    .S(_02444_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _18470_ (.A(_02451_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _18471_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.spi_buffer[7] ),
    .S(_02444_),
    .X(_02452_));
 sky130_fd_sc_hd__clkbuf_1 _18472_ (.A(_02452_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _18473_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.spi_buffer[8] ),
    .S(_02444_),
    .X(_02453_));
 sky130_fd_sc_hd__clkbuf_1 _18474_ (.A(_02453_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _18475_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.spi_buffer[9] ),
    .S(_02444_),
    .X(_02454_));
 sky130_fd_sc_hd__clkbuf_1 _18476_ (.A(_02454_),
    .X(_00924_));
 sky130_fd_sc_hd__clkbuf_4 _18477_ (.A(_02443_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _18478_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.spi_buffer[10] ),
    .S(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__clkbuf_1 _18479_ (.A(_02456_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _18480_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.spi_buffer[11] ),
    .S(_02455_),
    .X(_02457_));
 sky130_fd_sc_hd__clkbuf_1 _18481_ (.A(_02457_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _18482_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.spi_buffer[12] ),
    .S(_02455_),
    .X(_02458_));
 sky130_fd_sc_hd__clkbuf_1 _18483_ (.A(_02458_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _18484_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.spi_buffer[13] ),
    .S(_02455_),
    .X(_02459_));
 sky130_fd_sc_hd__clkbuf_1 _18485_ (.A(_02459_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _18486_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.spi_buffer[14] ),
    .S(_02455_),
    .X(_02460_));
 sky130_fd_sc_hd__clkbuf_1 _18487_ (.A(_02460_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _18488_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.spi_buffer[15] ),
    .S(_02455_),
    .X(_02461_));
 sky130_fd_sc_hd__clkbuf_1 _18489_ (.A(_02461_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _18490_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.spi_buffer[16] ),
    .S(_02455_),
    .X(_02462_));
 sky130_fd_sc_hd__clkbuf_1 _18491_ (.A(_02462_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _18492_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.spi_buffer[17] ),
    .S(_02455_),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_1 _18493_ (.A(_02463_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _18494_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.spi_buffer[18] ),
    .S(_02455_),
    .X(_02464_));
 sky130_fd_sc_hd__clkbuf_1 _18495_ (.A(_02464_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _18496_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.spi_buffer[19] ),
    .S(_02455_),
    .X(_02465_));
 sky130_fd_sc_hd__clkbuf_1 _18497_ (.A(_02465_),
    .X(_00934_));
 sky130_fd_sc_hd__clkbuf_4 _18498_ (.A(_02443_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _18499_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.spi_buffer[20] ),
    .S(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__clkbuf_1 _18500_ (.A(_02467_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _18501_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.spi_buffer[21] ),
    .S(_02466_),
    .X(_02468_));
 sky130_fd_sc_hd__clkbuf_1 _18502_ (.A(_02468_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _18503_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.spi_buffer[22] ),
    .S(_02466_),
    .X(_02469_));
 sky130_fd_sc_hd__clkbuf_1 _18504_ (.A(_02469_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _18505_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.spi_buffer[23] ),
    .S(_02466_),
    .X(_02470_));
 sky130_fd_sc_hd__clkbuf_1 _18506_ (.A(_02470_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _18507_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.spi_buffer[24] ),
    .S(_02466_),
    .X(_02471_));
 sky130_fd_sc_hd__clkbuf_1 _18508_ (.A(_02471_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _18509_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.spi_buffer[25] ),
    .S(_02466_),
    .X(_02472_));
 sky130_fd_sc_hd__clkbuf_1 _18510_ (.A(_02472_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _18511_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.spi_buffer[26] ),
    .S(_02466_),
    .X(_02473_));
 sky130_fd_sc_hd__clkbuf_1 _18512_ (.A(_02473_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _18513_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.spi_buffer[27] ),
    .S(_02466_),
    .X(_02474_));
 sky130_fd_sc_hd__clkbuf_1 _18514_ (.A(_02474_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _18515_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.spi_buffer[28] ),
    .S(_02466_),
    .X(_02475_));
 sky130_fd_sc_hd__clkbuf_1 _18516_ (.A(_02475_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _18517_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.spi_buffer[29] ),
    .S(_02466_),
    .X(_02476_));
 sky130_fd_sc_hd__clkbuf_1 _18518_ (.A(_02476_),
    .X(_00944_));
 sky130_fd_sc_hd__clkbuf_4 _18519_ (.A(_02443_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _18520_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.spi_buffer[30] ),
    .S(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__clkbuf_1 _18521_ (.A(_02478_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _18522_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.spi_buffer[31] ),
    .S(_02477_),
    .X(_02479_));
 sky130_fd_sc_hd__clkbuf_1 _18523_ (.A(_02479_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _18524_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.spi_buffer[32] ),
    .S(_02477_),
    .X(_02480_));
 sky130_fd_sc_hd__clkbuf_1 _18525_ (.A(_02480_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _18526_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.spi_buffer[33] ),
    .S(_02477_),
    .X(_02481_));
 sky130_fd_sc_hd__clkbuf_1 _18527_ (.A(_02481_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _18528_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.spi_buffer[34] ),
    .S(_02477_),
    .X(_02482_));
 sky130_fd_sc_hd__clkbuf_1 _18529_ (.A(_02482_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _18530_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.spi_buffer[35] ),
    .S(_02477_),
    .X(_02483_));
 sky130_fd_sc_hd__clkbuf_1 _18531_ (.A(_02483_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _18532_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.spi_buffer[36] ),
    .S(_02477_),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_1 _18533_ (.A(_02484_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _18534_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.spi_buffer[37] ),
    .S(_02477_),
    .X(_02485_));
 sky130_fd_sc_hd__clkbuf_1 _18535_ (.A(_02485_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _18536_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.spi_buffer[38] ),
    .S(_02477_),
    .X(_02486_));
 sky130_fd_sc_hd__clkbuf_1 _18537_ (.A(_02486_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _18538_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.spi_buffer[39] ),
    .S(_02477_),
    .X(_02487_));
 sky130_fd_sc_hd__clkbuf_1 _18539_ (.A(_02487_),
    .X(_00954_));
 sky130_fd_sc_hd__clkbuf_4 _18540_ (.A(_02443_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _18541_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.spi_buffer[40] ),
    .S(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__clkbuf_1 _18542_ (.A(_02489_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _18543_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.spi_buffer[41] ),
    .S(_02488_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _18544_ (.A(_02490_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _18545_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.spi_buffer[42] ),
    .S(_02488_),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_1 _18546_ (.A(_02491_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _18547_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.spi_buffer[43] ),
    .S(_02488_),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_1 _18548_ (.A(_02492_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _18549_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.spi_buffer[44] ),
    .S(_02488_),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _18550_ (.A(_02493_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _18551_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.spi_buffer[45] ),
    .S(_02488_),
    .X(_02494_));
 sky130_fd_sc_hd__clkbuf_1 _18552_ (.A(_02494_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _18553_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.spi_buffer[46] ),
    .S(_02488_),
    .X(_02495_));
 sky130_fd_sc_hd__clkbuf_1 _18554_ (.A(_02495_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _18555_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.spi_buffer[47] ),
    .S(_02488_),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_1 _18556_ (.A(_02496_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _18557_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.spi_buffer[48] ),
    .S(_02488_),
    .X(_02497_));
 sky130_fd_sc_hd__clkbuf_1 _18558_ (.A(_02497_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _18559_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.spi_buffer[49] ),
    .S(_02488_),
    .X(_02498_));
 sky130_fd_sc_hd__clkbuf_1 _18560_ (.A(_02498_),
    .X(_00964_));
 sky130_fd_sc_hd__clkbuf_4 _18561_ (.A(_02443_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _18562_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.spi_buffer[50] ),
    .S(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__clkbuf_1 _18563_ (.A(_02500_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _18564_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.spi_buffer[51] ),
    .S(_02499_),
    .X(_02501_));
 sky130_fd_sc_hd__clkbuf_1 _18565_ (.A(_02501_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _18566_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.spi_buffer[52] ),
    .S(_02499_),
    .X(_02502_));
 sky130_fd_sc_hd__clkbuf_1 _18567_ (.A(_02502_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _18568_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.spi_buffer[53] ),
    .S(_02499_),
    .X(_02503_));
 sky130_fd_sc_hd__clkbuf_1 _18569_ (.A(_02503_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _18570_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.spi_buffer[54] ),
    .S(_02499_),
    .X(_02504_));
 sky130_fd_sc_hd__clkbuf_1 _18571_ (.A(_02504_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _18572_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.spi_buffer[55] ),
    .S(_02499_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _18573_ (.A(_02505_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _18574_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.spi_buffer[56] ),
    .S(_02499_),
    .X(_02506_));
 sky130_fd_sc_hd__clkbuf_1 _18575_ (.A(_02506_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _18576_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.spi_buffer[57] ),
    .S(_02499_),
    .X(_02507_));
 sky130_fd_sc_hd__clkbuf_1 _18577_ (.A(_02507_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _18578_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.spi_buffer[58] ),
    .S(_02499_),
    .X(_02508_));
 sky130_fd_sc_hd__clkbuf_1 _18579_ (.A(_02508_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _18580_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.spi_buffer[59] ),
    .S(_02499_),
    .X(_02509_));
 sky130_fd_sc_hd__clkbuf_1 _18581_ (.A(_02509_),
    .X(_00974_));
 sky130_fd_sc_hd__buf_4 _18582_ (.A(_02442_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _18583_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.spi_buffer[60] ),
    .S(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__clkbuf_1 _18584_ (.A(_02511_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _18585_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.spi_buffer[61] ),
    .S(_02510_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _18586_ (.A(_02512_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _18587_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.spi_buffer[62] ),
    .S(_02510_),
    .X(_02513_));
 sky130_fd_sc_hd__clkbuf_1 _18588_ (.A(_02513_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _18589_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.spi_buffer[63] ),
    .S(_02510_),
    .X(_02514_));
 sky130_fd_sc_hd__clkbuf_1 _18590_ (.A(_02514_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _18591_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.spi_buffer[64] ),
    .S(_02510_),
    .X(_02515_));
 sky130_fd_sc_hd__clkbuf_1 _18592_ (.A(_02515_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _18593_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.spi_buffer[65] ),
    .S(_02510_),
    .X(_02516_));
 sky130_fd_sc_hd__clkbuf_1 _18594_ (.A(_02516_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _18595_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.spi_buffer[66] ),
    .S(_02510_),
    .X(_02517_));
 sky130_fd_sc_hd__clkbuf_1 _18596_ (.A(_02517_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _18597_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.spi_buffer[67] ),
    .S(_02510_),
    .X(_02518_));
 sky130_fd_sc_hd__clkbuf_1 _18598_ (.A(_02518_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _18599_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.spi_buffer[68] ),
    .S(_02510_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_1 _18600_ (.A(_02519_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _18601_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.spi_buffer[69] ),
    .S(_02510_),
    .X(_02520_));
 sky130_fd_sc_hd__clkbuf_1 _18602_ (.A(_02520_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _18603_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.spi_buffer[70] ),
    .S(_02443_),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _18604_ (.A(_02521_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _18605_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.spi_buffer[71] ),
    .S(_02443_),
    .X(_02522_));
 sky130_fd_sc_hd__clkbuf_1 _18606_ (.A(_02522_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _18607_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.spi_buffer[72] ),
    .S(_02443_),
    .X(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _18608_ (.A(_02523_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _18609_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.spi_buffer[73] ),
    .S(_02443_),
    .X(_02524_));
 sky130_fd_sc_hd__clkbuf_1 _18610_ (.A(_02524_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _18611_ (.A0(_04532_),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_03337_),
    .X(_02525_));
 sky130_fd_sc_hd__clkbuf_1 _18612_ (.A(_02525_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _18613_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_04827_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_1 _18614_ (.A(_02526_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _18615_ (.A0(net51),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_03337_),
    .X(_02527_));
 sky130_fd_sc_hd__clkbuf_1 _18616_ (.A(_02527_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _18617_ (.A0(\rbzero.pov.ss_buffer[1] ),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_04827_),
    .X(_02528_));
 sky130_fd_sc_hd__clkbuf_1 _18618_ (.A(_02528_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _18619_ (.A0(net53),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_03337_),
    .X(_02529_));
 sky130_fd_sc_hd__clkbuf_1 _18620_ (.A(_02529_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _18621_ (.A0(\rbzero.pov.sclk_buffer[1] ),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_04827_),
    .X(_02530_));
 sky130_fd_sc_hd__clkbuf_1 _18622_ (.A(_02530_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _18623_ (.A0(\rbzero.pov.sclk_buffer[2] ),
    .A1(\rbzero.pov.sclk_buffer[1] ),
    .S(_04827_),
    .X(_02531_));
 sky130_fd_sc_hd__clkbuf_1 _18624_ (.A(_02531_),
    .X(_00995_));
 sky130_fd_sc_hd__and2_1 _18625_ (.A(\rbzero.pov.ready ),
    .B(_02412_),
    .X(_02532_));
 sky130_fd_sc_hd__o21ai_4 _18626_ (.A1(net39),
    .A2(_02532_),
    .B1(_02262_),
    .Y(_02533_));
 sky130_fd_sc_hd__clkbuf_4 _18627_ (.A(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__clkbuf_4 _18628_ (.A(_02412_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _18629_ (.A0(_07145_),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__nand2_1 _18630_ (.A(_07145_),
    .B(_02533_),
    .Y(_02537_));
 sky130_fd_sc_hd__o211a_1 _18631_ (.A1(_02534_),
    .A2(_02536_),
    .B1(_02537_),
    .C1(_02356_),
    .X(_00996_));
 sky130_fd_sc_hd__and2_1 _18632_ (.A(_02261_),
    .B(_02411_),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_4 _18633_ (.A(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__clkbuf_4 _18634_ (.A(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _18635_ (.A0(\rbzero.pov.ready_buffer[60] ),
    .A1(_06912_),
    .S(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__o21a_2 _18636_ (.A1(net39),
    .A2(_02532_),
    .B1(_02261_),
    .X(_02542_));
 sky130_fd_sc_hd__clkbuf_4 _18637_ (.A(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__or2_1 _18638_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__o211a_1 _18639_ (.A1(_02534_),
    .A2(_02541_),
    .B1(_02544_),
    .C1(_02356_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _18640_ (.A0(\rbzero.pov.ready_buffer[61] ),
    .A1(_06890_),
    .S(_02540_),
    .X(_02545_));
 sky130_fd_sc_hd__or2_1 _18641_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(_02542_),
    .X(_02546_));
 sky130_fd_sc_hd__o211a_1 _18642_ (.A1(_02534_),
    .A2(_02545_),
    .B1(_02546_),
    .C1(_02356_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _18643_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(_06929_),
    .S(_02540_),
    .X(_02547_));
 sky130_fd_sc_hd__or2_1 _18644_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_02542_),
    .X(_02548_));
 sky130_fd_sc_hd__o211a_1 _18645_ (.A1(_02534_),
    .A2(_02547_),
    .B1(_02548_),
    .C1(_02356_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _18646_ (.A0(\rbzero.pov.ready_buffer[63] ),
    .A1(_06946_),
    .S(_02540_),
    .X(_02549_));
 sky130_fd_sc_hd__or2_1 _18647_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_02542_),
    .X(_02550_));
 sky130_fd_sc_hd__o211a_1 _18648_ (.A1(_02534_),
    .A2(_02549_),
    .B1(_02550_),
    .C1(_02356_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _18649_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(_06963_),
    .S(_02539_),
    .X(_02551_));
 sky130_fd_sc_hd__or2_1 _18650_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(_02542_),
    .X(_02552_));
 sky130_fd_sc_hd__o211a_1 _18651_ (.A1(_02534_),
    .A2(_02551_),
    .B1(_02552_),
    .C1(_02356_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _18652_ (.A0(\rbzero.pov.ready_buffer[65] ),
    .A1(_06989_),
    .S(_02539_),
    .X(_02553_));
 sky130_fd_sc_hd__nand2_1 _18653_ (.A(_06990_),
    .B(_02533_),
    .Y(_02554_));
 sky130_fd_sc_hd__o211a_1 _18654_ (.A1(_02534_),
    .A2(_02553_),
    .B1(_02554_),
    .C1(_02356_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _18655_ (.A0(\rbzero.pov.ready_buffer[66] ),
    .A1(_07021_),
    .S(_02539_),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _18656_ (.A(_07022_),
    .B(_02533_),
    .Y(_02556_));
 sky130_fd_sc_hd__o211a_1 _18657_ (.A1(_02534_),
    .A2(_02555_),
    .B1(_02556_),
    .C1(_02356_),
    .X(_01003_));
 sky130_fd_sc_hd__inv_2 _18658_ (.A(_07034_),
    .Y(_02557_));
 sky130_fd_sc_hd__o221a_1 _18659_ (.A1(\rbzero.pov.ready_buffer[67] ),
    .A2(_02411_),
    .B1(_02413_),
    .B2(_02557_),
    .C1(_02543_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_4 _18660_ (.A(_03338_),
    .X(_02559_));
 sky130_fd_sc_hd__a211o_1 _18661_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_02534_),
    .B1(_02558_),
    .C1(_02559_),
    .X(_01004_));
 sky130_fd_sc_hd__nand2_1 _18662_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_07032_),
    .Y(_02560_));
 sky130_fd_sc_hd__or2_1 _18663_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_07032_),
    .X(_02561_));
 sky130_fd_sc_hd__nand2_1 _18664_ (.A(_02560_),
    .B(_02561_),
    .Y(_02562_));
 sky130_fd_sc_hd__o221a_1 _18665_ (.A1(\rbzero.pov.ready_buffer[68] ),
    .A2(_02411_),
    .B1(_02413_),
    .B2(_02562_),
    .C1(_02543_),
    .X(_02563_));
 sky130_fd_sc_hd__a211o_1 _18666_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_02534_),
    .B1(_02563_),
    .C1(_02559_),
    .X(_01005_));
 sky130_fd_sc_hd__xnor2_1 _18667_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_02561_),
    .Y(_02564_));
 sky130_fd_sc_hd__o221a_1 _18668_ (.A1(\rbzero.pov.ready_buffer[69] ),
    .A2(_02411_),
    .B1(_02535_),
    .B2(_02564_),
    .C1(_02543_),
    .X(_02565_));
 sky130_fd_sc_hd__a211o_1 _18669_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_02533_),
    .B1(_02565_),
    .C1(_02559_),
    .X(_01006_));
 sky130_fd_sc_hd__or3_1 _18670_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .B(\rbzero.debug_overlay.playerX[1] ),
    .C(_02561_),
    .X(_02566_));
 sky130_fd_sc_hd__o21ai_1 _18671_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_02561_),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .Y(_02567_));
 sky130_fd_sc_hd__a21oi_1 _18672_ (.A1(_02566_),
    .A2(_02567_),
    .B1(_02535_),
    .Y(_02568_));
 sky130_fd_sc_hd__a211o_1 _18673_ (.A1(\rbzero.pov.ready_buffer[70] ),
    .A2(_02413_),
    .B1(_02533_),
    .C1(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__o211a_1 _18674_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_02543_),
    .B1(_02569_),
    .C1(_02356_),
    .X(_01007_));
 sky130_fd_sc_hd__or2_1 _18675_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_02566_),
    .X(_02570_));
 sky130_fd_sc_hd__inv_2 _18676_ (.A(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__a21o_1 _18677_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_02566_),
    .B1(_02412_),
    .X(_02572_));
 sky130_fd_sc_hd__o221a_1 _18678_ (.A1(\rbzero.pov.ready_buffer[71] ),
    .A2(_02540_),
    .B1(_02571_),
    .B2(_02572_),
    .C1(_02543_),
    .X(_02573_));
 sky130_fd_sc_hd__a211o_1 _18679_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_02533_),
    .B1(_02573_),
    .C1(_02559_),
    .X(_01008_));
 sky130_fd_sc_hd__nand2_1 _18680_ (.A(_02411_),
    .B(_02570_),
    .Y(_02574_));
 sky130_fd_sc_hd__a21oi_1 _18681_ (.A1(_02543_),
    .A2(_02574_),
    .B1(_03350_),
    .Y(_02575_));
 sky130_fd_sc_hd__o21ai_1 _18682_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_02570_),
    .B1(_02411_),
    .Y(_02576_));
 sky130_fd_sc_hd__o211a_1 _18683_ (.A1(\rbzero.pov.ready_buffer[72] ),
    .A2(_02540_),
    .B1(_02543_),
    .C1(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__o21a_1 _18684_ (.A1(_02575_),
    .A2(_02577_),
    .B1(_02266_),
    .X(_01009_));
 sky130_fd_sc_hd__a21boi_1 _18685_ (.A1(_02543_),
    .A2(_02576_),
    .B1_N(\rbzero.debug_overlay.playerX[5] ),
    .Y(_02578_));
 sky130_fd_sc_hd__o31ai_1 _18686_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(\rbzero.debug_overlay.playerX[4] ),
    .A3(_02570_),
    .B1(_02540_),
    .Y(_02579_));
 sky130_fd_sc_hd__o211a_1 _18687_ (.A1(\rbzero.pov.ready_buffer[73] ),
    .A2(_02540_),
    .B1(_02543_),
    .C1(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__o21a_1 _18688_ (.A1(_02578_),
    .A2(_02580_),
    .B1(_02266_),
    .X(_01010_));
 sky130_fd_sc_hd__o21ai_1 _18689_ (.A1(net40),
    .A2(_02532_),
    .B1(_02262_),
    .Y(_02581_));
 sky130_fd_sc_hd__buf_2 _18690_ (.A(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__inv_2 _18691_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_02583_));
 sky130_fd_sc_hd__mux2_1 _18692_ (.A0(_02583_),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_02535_),
    .X(_02584_));
 sky130_fd_sc_hd__nand2_1 _18693_ (.A(_02583_),
    .B(_02582_),
    .Y(_02585_));
 sky130_fd_sc_hd__clkbuf_4 _18694_ (.A(_04828_),
    .X(_02586_));
 sky130_fd_sc_hd__o211a_1 _18695_ (.A1(_02582_),
    .A2(_02584_),
    .B1(_02585_),
    .C1(_02586_),
    .X(_01011_));
 sky130_fd_sc_hd__o21a_2 _18696_ (.A1(net40),
    .A2(_02532_),
    .B1(_02262_),
    .X(_02587_));
 sky130_fd_sc_hd__buf_2 _18697_ (.A(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__inv_2 _18698_ (.A(\rbzero.pov.ready_buffer[45] ),
    .Y(_02589_));
 sky130_fd_sc_hd__mux2_1 _18699_ (.A0(_02589_),
    .A1(_06909_),
    .S(_02539_),
    .X(_02590_));
 sky130_fd_sc_hd__nor2_1 _18700_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(_02588_),
    .Y(_02591_));
 sky130_fd_sc_hd__a211oi_1 _18701_ (.A1(_02588_),
    .A2(_02590_),
    .B1(_02591_),
    .C1(_02319_),
    .Y(_01012_));
 sky130_fd_sc_hd__nor2_1 _18702_ (.A(_06879_),
    .B(_02535_),
    .Y(_02592_));
 sky130_fd_sc_hd__a211o_1 _18703_ (.A1(\rbzero.pov.ready_buffer[46] ),
    .A2(_02413_),
    .B1(_02582_),
    .C1(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__o211a_1 _18704_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_02588_),
    .B1(_02593_),
    .C1(_02586_),
    .X(_01013_));
 sky130_fd_sc_hd__nor2_1 _18705_ (.A(_06924_),
    .B(_02535_),
    .Y(_02594_));
 sky130_fd_sc_hd__a211o_1 _18706_ (.A1(\rbzero.pov.ready_buffer[47] ),
    .A2(_02413_),
    .B1(_02582_),
    .C1(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__o211a_1 _18707_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_02588_),
    .B1(_02595_),
    .C1(_02586_),
    .X(_01014_));
 sky130_fd_sc_hd__inv_2 _18708_ (.A(\rbzero.pov.ready_buffer[48] ),
    .Y(_02596_));
 sky130_fd_sc_hd__mux2_1 _18709_ (.A0(_02596_),
    .A1(_06943_),
    .S(_02539_),
    .X(_02597_));
 sky130_fd_sc_hd__mux2_1 _18710_ (.A0(_06942_),
    .A1(_02597_),
    .S(_02587_),
    .X(_02598_));
 sky130_fd_sc_hd__nor2_1 _18711_ (.A(net61),
    .B(_02598_),
    .Y(_01015_));
 sky130_fd_sc_hd__nor2_1 _18712_ (.A(_06958_),
    .B(_02535_),
    .Y(_02599_));
 sky130_fd_sc_hd__a211o_1 _18713_ (.A1(\rbzero.pov.ready_buffer[49] ),
    .A2(_02413_),
    .B1(_02582_),
    .C1(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__o211a_1 _18714_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_02588_),
    .B1(_02600_),
    .C1(_02586_),
    .X(_01016_));
 sky130_fd_sc_hd__nor2_1 _18715_ (.A(_06982_),
    .B(_02535_),
    .Y(_02601_));
 sky130_fd_sc_hd__a211o_1 _18716_ (.A1(\rbzero.pov.ready_buffer[50] ),
    .A2(_02413_),
    .B1(_02582_),
    .C1(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__o211a_1 _18717_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_02588_),
    .B1(_02602_),
    .C1(_02586_),
    .X(_01017_));
 sky130_fd_sc_hd__inv_2 _18718_ (.A(\rbzero.pov.ready_buffer[51] ),
    .Y(_02603_));
 sky130_fd_sc_hd__mux2_1 _18719_ (.A0(_02603_),
    .A1(_07017_),
    .S(_02539_),
    .X(_02604_));
 sky130_fd_sc_hd__mux2_1 _18720_ (.A0(_07016_),
    .A1(_02604_),
    .S(_02587_),
    .X(_02605_));
 sky130_fd_sc_hd__nor2_1 _18721_ (.A(net61),
    .B(_02605_),
    .Y(_01018_));
 sky130_fd_sc_hd__o221a_1 _18722_ (.A1(\rbzero.pov.ready_buffer[52] ),
    .A2(_02411_),
    .B1(_02535_),
    .B2(_07028_),
    .C1(_02587_),
    .X(_02606_));
 sky130_fd_sc_hd__a211o_1 _18723_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_02582_),
    .B1(_02606_),
    .C1(_02559_),
    .X(_01019_));
 sky130_fd_sc_hd__nor2_1 _18724_ (.A(net40),
    .B(net39),
    .Y(_02607_));
 sky130_fd_sc_hd__xnor2_1 _18725_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_07026_),
    .Y(_02608_));
 sky130_fd_sc_hd__a221o_1 _18726_ (.A1(\rbzero.pov.ready_buffer[53] ),
    .A2(_02607_),
    .B1(_02540_),
    .B2(_02608_),
    .C1(_02581_),
    .X(_02609_));
 sky130_fd_sc_hd__o211a_1 _18727_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_02588_),
    .B1(_02609_),
    .C1(_02586_),
    .X(_01020_));
 sky130_fd_sc_hd__or3_1 _18728_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .C(_07026_),
    .X(_02610_));
 sky130_fd_sc_hd__o21ai_1 _18729_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_07026_),
    .B1(\rbzero.debug_overlay.playerY[1] ),
    .Y(_02611_));
 sky130_fd_sc_hd__nand2_1 _18730_ (.A(_02610_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__o221a_1 _18731_ (.A1(\rbzero.pov.ready_buffer[54] ),
    .A2(_02411_),
    .B1(_02535_),
    .B2(_02612_),
    .C1(_02587_),
    .X(_02613_));
 sky130_fd_sc_hd__a211o_1 _18732_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_02582_),
    .B1(_02613_),
    .C1(_02559_),
    .X(_01021_));
 sky130_fd_sc_hd__or2_1 _18733_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(_02610_),
    .X(_02614_));
 sky130_fd_sc_hd__nand2_1 _18734_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(_02610_),
    .Y(_02615_));
 sky130_fd_sc_hd__a21oi_1 _18735_ (.A1(_02614_),
    .A2(_02615_),
    .B1(_02412_),
    .Y(_02616_));
 sky130_fd_sc_hd__a211o_1 _18736_ (.A1(\rbzero.pov.ready_buffer[55] ),
    .A2(_02413_),
    .B1(_02582_),
    .C1(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__o211a_1 _18737_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_02588_),
    .B1(_02617_),
    .C1(_02586_),
    .X(_01022_));
 sky130_fd_sc_hd__nor2_1 _18738_ (.A(_03347_),
    .B(_02587_),
    .Y(_02618_));
 sky130_fd_sc_hd__or2_1 _18739_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .B(_02614_),
    .X(_02619_));
 sky130_fd_sc_hd__inv_2 _18740_ (.A(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__a21o_1 _18741_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_02614_),
    .B1(_02412_),
    .X(_02621_));
 sky130_fd_sc_hd__o221a_1 _18742_ (.A1(\rbzero.pov.ready_buffer[56] ),
    .A2(_02539_),
    .B1(_02620_),
    .B2(_02621_),
    .C1(_02587_),
    .X(_02622_));
 sky130_fd_sc_hd__or3_1 _18743_ (.A(_03337_),
    .B(_02618_),
    .C(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_1 _18744_ (.A(_02623_),
    .X(_01023_));
 sky130_fd_sc_hd__nor2_1 _18745_ (.A(_02607_),
    .B(_02620_),
    .Y(_02624_));
 sky130_fd_sc_hd__o21a_1 _18746_ (.A1(_02582_),
    .A2(_02624_),
    .B1(\rbzero.debug_overlay.playerY[4] ),
    .X(_02625_));
 sky130_fd_sc_hd__o21ai_1 _18747_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_02619_),
    .B1(_02411_),
    .Y(_02626_));
 sky130_fd_sc_hd__o211a_1 _18748_ (.A1(\rbzero.pov.ready_buffer[57] ),
    .A2(_02540_),
    .B1(_02588_),
    .C1(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__o21a_1 _18749_ (.A1(_02625_),
    .A2(_02627_),
    .B1(_02266_),
    .X(_01024_));
 sky130_fd_sc_hd__a21o_1 _18750_ (.A1(_02588_),
    .A2(_02626_),
    .B1(_03360_),
    .X(_02628_));
 sky130_fd_sc_hd__inv_2 _18751_ (.A(\rbzero.pov.ready_buffer[58] ),
    .Y(_02629_));
 sky130_fd_sc_hd__o31a_1 _18752_ (.A1(\rbzero.debug_overlay.playerY[5] ),
    .A2(\rbzero.debug_overlay.playerY[4] ),
    .A3(_02619_),
    .B1(_02539_),
    .X(_02630_));
 sky130_fd_sc_hd__a211o_1 _18753_ (.A1(_02629_),
    .A2(_02413_),
    .B1(_02581_),
    .C1(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__a21oi_1 _18754_ (.A1(_02628_),
    .A2(_02631_),
    .B1(_02559_),
    .Y(_01025_));
 sky130_fd_sc_hd__and2_1 _18755_ (.A(\rbzero.pov.ready ),
    .B(_02607_),
    .X(_02632_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(_02288_),
    .B(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__buf_2 _18757_ (.A(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__buf_2 _18758_ (.A(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__buf_2 _18759_ (.A(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__and2_1 _18760_ (.A(_02288_),
    .B(_02632_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_2 _18761_ (.A(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__or2_1 _18762_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__o211a_1 _18763_ (.A1(\rbzero.pov.ready_buffer[33] ),
    .A2(_02636_),
    .B1(_02639_),
    .C1(_02586_),
    .X(_01026_));
 sky130_fd_sc_hd__or2_1 _18764_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(_02638_),
    .X(_02640_));
 sky130_fd_sc_hd__o211a_1 _18765_ (.A1(\rbzero.pov.ready_buffer[34] ),
    .A2(_02636_),
    .B1(_02640_),
    .C1(_02586_),
    .X(_01027_));
 sky130_fd_sc_hd__or2_1 _18766_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(_02638_),
    .X(_02641_));
 sky130_fd_sc_hd__o211a_1 _18767_ (.A1(\rbzero.pov.ready_buffer[35] ),
    .A2(_02636_),
    .B1(_02641_),
    .C1(_02586_),
    .X(_01028_));
 sky130_fd_sc_hd__or2_1 _18768_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(_02638_),
    .X(_02642_));
 sky130_fd_sc_hd__buf_2 _18769_ (.A(_04828_),
    .X(_02643_));
 sky130_fd_sc_hd__o211a_1 _18770_ (.A1(\rbzero.pov.ready_buffer[36] ),
    .A2(_02636_),
    .B1(_02642_),
    .C1(_02643_),
    .X(_01029_));
 sky130_fd_sc_hd__clkbuf_4 _18771_ (.A(_02638_),
    .X(_02644_));
 sky130_fd_sc_hd__buf_2 _18772_ (.A(_02633_),
    .X(_02645_));
 sky130_fd_sc_hd__and2_1 _18773_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__a211o_1 _18774_ (.A1(\rbzero.pov.ready_buffer[37] ),
    .A2(_02644_),
    .B1(_02646_),
    .C1(_02559_),
    .X(_01030_));
 sky130_fd_sc_hd__and2_1 _18775_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(_02645_),
    .X(_02647_));
 sky130_fd_sc_hd__a211o_1 _18776_ (.A1(\rbzero.pov.ready_buffer[38] ),
    .A2(_02644_),
    .B1(_02647_),
    .C1(_02559_),
    .X(_01031_));
 sky130_fd_sc_hd__and2_1 _18777_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(_02645_),
    .X(_02648_));
 sky130_fd_sc_hd__a211o_1 _18778_ (.A1(\rbzero.pov.ready_buffer[39] ),
    .A2(_02644_),
    .B1(_02648_),
    .C1(_02559_),
    .X(_01032_));
 sky130_fd_sc_hd__or2_1 _18779_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(_02638_),
    .X(_02649_));
 sky130_fd_sc_hd__o211a_1 _18780_ (.A1(\rbzero.pov.ready_buffer[40] ),
    .A2(_02636_),
    .B1(_02649_),
    .C1(_02643_),
    .X(_01033_));
 sky130_fd_sc_hd__and2_1 _18781_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(_02645_),
    .X(_02650_));
 sky130_fd_sc_hd__clkbuf_4 _18782_ (.A(_03338_),
    .X(_02651_));
 sky130_fd_sc_hd__a211o_1 _18783_ (.A1(\rbzero.pov.ready_buffer[41] ),
    .A2(_02644_),
    .B1(_02650_),
    .C1(_02651_),
    .X(_01034_));
 sky130_fd_sc_hd__or2_1 _18784_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(_02638_),
    .X(_02652_));
 sky130_fd_sc_hd__o211a_1 _18785_ (.A1(\rbzero.pov.ready_buffer[42] ),
    .A2(_02636_),
    .B1(_02652_),
    .C1(_02643_),
    .X(_01035_));
 sky130_fd_sc_hd__or2_1 _18786_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(_02638_),
    .X(_02653_));
 sky130_fd_sc_hd__o211a_1 _18787_ (.A1(\rbzero.pov.ready_buffer[43] ),
    .A2(_02636_),
    .B1(_02653_),
    .C1(_02643_),
    .X(_01036_));
 sky130_fd_sc_hd__and2_1 _18788_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(_02645_),
    .X(_02654_));
 sky130_fd_sc_hd__a211o_1 _18789_ (.A1(\rbzero.pov.ready_buffer[22] ),
    .A2(_02644_),
    .B1(_02654_),
    .C1(_02651_),
    .X(_01037_));
 sky130_fd_sc_hd__or2_1 _18790_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_02638_),
    .X(_02655_));
 sky130_fd_sc_hd__o211a_1 _18791_ (.A1(\rbzero.pov.ready_buffer[23] ),
    .A2(_02636_),
    .B1(_02655_),
    .C1(_02643_),
    .X(_01038_));
 sky130_fd_sc_hd__and2_1 _18792_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(_02645_),
    .X(_02656_));
 sky130_fd_sc_hd__a211o_1 _18793_ (.A1(\rbzero.pov.ready_buffer[24] ),
    .A2(_02644_),
    .B1(_02656_),
    .C1(_02651_),
    .X(_01039_));
 sky130_fd_sc_hd__and2_1 _18794_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(_02645_),
    .X(_02657_));
 sky130_fd_sc_hd__a211o_1 _18795_ (.A1(\rbzero.pov.ready_buffer[25] ),
    .A2(_02644_),
    .B1(_02657_),
    .C1(_02651_),
    .X(_01040_));
 sky130_fd_sc_hd__and2_1 _18796_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(_02645_),
    .X(_02658_));
 sky130_fd_sc_hd__a211o_1 _18797_ (.A1(\rbzero.pov.ready_buffer[26] ),
    .A2(_02644_),
    .B1(_02658_),
    .C1(_02651_),
    .X(_01041_));
 sky130_fd_sc_hd__or2_1 _18798_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(_02638_),
    .X(_02659_));
 sky130_fd_sc_hd__o211a_1 _18799_ (.A1(\rbzero.pov.ready_buffer[27] ),
    .A2(_02636_),
    .B1(_02659_),
    .C1(_02643_),
    .X(_01042_));
 sky130_fd_sc_hd__clkbuf_2 _18800_ (.A(_02637_),
    .X(_02660_));
 sky130_fd_sc_hd__or2_1 _18801_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__o211a_1 _18802_ (.A1(\rbzero.pov.ready_buffer[28] ),
    .A2(_02636_),
    .B1(_02661_),
    .C1(_02643_),
    .X(_01043_));
 sky130_fd_sc_hd__and2_1 _18803_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(_02645_),
    .X(_02662_));
 sky130_fd_sc_hd__a211o_1 _18804_ (.A1(\rbzero.pov.ready_buffer[29] ),
    .A2(_02644_),
    .B1(_02662_),
    .C1(_02651_),
    .X(_01044_));
 sky130_fd_sc_hd__buf_2 _18805_ (.A(_02645_),
    .X(_02663_));
 sky130_fd_sc_hd__or2_1 _18806_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(_02660_),
    .X(_02664_));
 sky130_fd_sc_hd__o211a_1 _18807_ (.A1(\rbzero.pov.ready_buffer[30] ),
    .A2(_02663_),
    .B1(_02664_),
    .C1(_02643_),
    .X(_01045_));
 sky130_fd_sc_hd__and2_1 _18808_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(_02634_),
    .X(_02665_));
 sky130_fd_sc_hd__a211o_1 _18809_ (.A1(\rbzero.pov.ready_buffer[31] ),
    .A2(_02644_),
    .B1(_02665_),
    .C1(_02651_),
    .X(_01046_));
 sky130_fd_sc_hd__clkbuf_4 _18810_ (.A(_02637_),
    .X(_02666_));
 sky130_fd_sc_hd__and2_1 _18811_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(_02634_),
    .X(_02667_));
 sky130_fd_sc_hd__a211o_1 _18812_ (.A1(\rbzero.pov.ready_buffer[32] ),
    .A2(_02666_),
    .B1(_02667_),
    .C1(_02651_),
    .X(_01047_));
 sky130_fd_sc_hd__nor2_1 _18813_ (.A(_01967_),
    .B(_02666_),
    .Y(_02668_));
 sky130_fd_sc_hd__a211o_1 _18814_ (.A1(\rbzero.pov.ready_buffer[11] ),
    .A2(_02666_),
    .B1(_02668_),
    .C1(_02651_),
    .X(_01048_));
 sky130_fd_sc_hd__or2_1 _18815_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(_02660_),
    .X(_02669_));
 sky130_fd_sc_hd__o211a_1 _18816_ (.A1(\rbzero.pov.ready_buffer[12] ),
    .A2(_02663_),
    .B1(_02669_),
    .C1(_02643_),
    .X(_01049_));
 sky130_fd_sc_hd__or2_1 _18817_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02660_),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_1 _18818_ (.A1(\rbzero.pov.ready_buffer[13] ),
    .A2(_02663_),
    .B1(_02670_),
    .C1(_02643_),
    .X(_01050_));
 sky130_fd_sc_hd__or2_1 _18819_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_02660_),
    .X(_02671_));
 sky130_fd_sc_hd__buf_2 _18820_ (.A(_04828_),
    .X(_02672_));
 sky130_fd_sc_hd__o211a_1 _18821_ (.A1(\rbzero.pov.ready_buffer[14] ),
    .A2(_02663_),
    .B1(_02671_),
    .C1(_02672_),
    .X(_01051_));
 sky130_fd_sc_hd__and2_1 _18822_ (.A(_04100_),
    .B(_02634_),
    .X(_02673_));
 sky130_fd_sc_hd__a211o_1 _18823_ (.A1(\rbzero.pov.ready_buffer[15] ),
    .A2(_02666_),
    .B1(_02673_),
    .C1(_02651_),
    .X(_01052_));
 sky130_fd_sc_hd__and2_1 _18824_ (.A(_04102_),
    .B(_02634_),
    .X(_02674_));
 sky130_fd_sc_hd__buf_4 _18825_ (.A(_03338_),
    .X(_02675_));
 sky130_fd_sc_hd__a211o_1 _18826_ (.A1(\rbzero.pov.ready_buffer[16] ),
    .A2(_02666_),
    .B1(_02674_),
    .C1(_02675_),
    .X(_01053_));
 sky130_fd_sc_hd__or2_1 _18827_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(_02660_),
    .X(_02676_));
 sky130_fd_sc_hd__o211a_1 _18828_ (.A1(\rbzero.pov.ready_buffer[17] ),
    .A2(_02663_),
    .B1(_02676_),
    .C1(_02672_),
    .X(_01054_));
 sky130_fd_sc_hd__and2_1 _18829_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(_02634_),
    .X(_02677_));
 sky130_fd_sc_hd__a211o_1 _18830_ (.A1(\rbzero.pov.ready_buffer[18] ),
    .A2(_02666_),
    .B1(_02677_),
    .C1(_02675_),
    .X(_01055_));
 sky130_fd_sc_hd__or2_1 _18831_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_02660_),
    .X(_02678_));
 sky130_fd_sc_hd__o211a_1 _18832_ (.A1(\rbzero.pov.ready_buffer[19] ),
    .A2(_02663_),
    .B1(_02678_),
    .C1(_02672_),
    .X(_01056_));
 sky130_fd_sc_hd__nand2_1 _18833_ (.A(_02081_),
    .B(_02635_),
    .Y(_02679_));
 sky130_fd_sc_hd__o211a_1 _18834_ (.A1(\rbzero.pov.ready_buffer[20] ),
    .A2(_02663_),
    .B1(_02679_),
    .C1(_02672_),
    .X(_01057_));
 sky130_fd_sc_hd__nand2_1 _18835_ (.A(_02094_),
    .B(_02635_),
    .Y(_02680_));
 sky130_fd_sc_hd__o211a_1 _18836_ (.A1(\rbzero.pov.ready_buffer[21] ),
    .A2(_02663_),
    .B1(_02680_),
    .C1(_02672_),
    .X(_01058_));
 sky130_fd_sc_hd__nand2_1 _18837_ (.A(_01752_),
    .B(_02635_),
    .Y(_02681_));
 sky130_fd_sc_hd__o211a_1 _18838_ (.A1(\rbzero.pov.ready_buffer[0] ),
    .A2(_02663_),
    .B1(_02681_),
    .C1(_02672_),
    .X(_01059_));
 sky130_fd_sc_hd__or2_1 _18839_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_02660_),
    .X(_02682_));
 sky130_fd_sc_hd__o211a_1 _18840_ (.A1(\rbzero.pov.ready_buffer[1] ),
    .A2(_02663_),
    .B1(_02682_),
    .C1(_02672_),
    .X(_01060_));
 sky130_fd_sc_hd__or2_1 _18841_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02660_),
    .X(_02683_));
 sky130_fd_sc_hd__o211a_1 _18842_ (.A1(\rbzero.pov.ready_buffer[2] ),
    .A2(_02635_),
    .B1(_02683_),
    .C1(_02672_),
    .X(_01061_));
 sky130_fd_sc_hd__and2_1 _18843_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_02634_),
    .X(_02684_));
 sky130_fd_sc_hd__a211o_1 _18844_ (.A1(\rbzero.pov.ready_buffer[3] ),
    .A2(_02666_),
    .B1(_02684_),
    .C1(_02675_),
    .X(_01062_));
 sky130_fd_sc_hd__and2_1 _18845_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(_02634_),
    .X(_02685_));
 sky130_fd_sc_hd__a211o_1 _18846_ (.A1(\rbzero.pov.ready_buffer[4] ),
    .A2(_02666_),
    .B1(_02685_),
    .C1(_02675_),
    .X(_01063_));
 sky130_fd_sc_hd__and2_1 _18847_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(_02634_),
    .X(_02686_));
 sky130_fd_sc_hd__a211o_1 _18848_ (.A1(\rbzero.pov.ready_buffer[5] ),
    .A2(_02666_),
    .B1(_02686_),
    .C1(_02675_),
    .X(_01064_));
 sky130_fd_sc_hd__or2_1 _18849_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(_02660_),
    .X(_02687_));
 sky130_fd_sc_hd__o211a_1 _18850_ (.A1(\rbzero.pov.ready_buffer[6] ),
    .A2(_02635_),
    .B1(_02687_),
    .C1(_02672_),
    .X(_01065_));
 sky130_fd_sc_hd__and2_1 _18851_ (.A(_04109_),
    .B(_02634_),
    .X(_02688_));
 sky130_fd_sc_hd__a211o_1 _18852_ (.A1(\rbzero.pov.ready_buffer[7] ),
    .A2(_02666_),
    .B1(_02688_),
    .C1(_02675_),
    .X(_01066_));
 sky130_fd_sc_hd__or2_1 _18853_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_02637_),
    .X(_02689_));
 sky130_fd_sc_hd__o211a_1 _18854_ (.A1(\rbzero.pov.ready_buffer[8] ),
    .A2(_02635_),
    .B1(_02689_),
    .C1(_02672_),
    .X(_01067_));
 sky130_fd_sc_hd__nand2_1 _18855_ (.A(_01871_),
    .B(_02635_),
    .Y(_02690_));
 sky130_fd_sc_hd__o211a_1 _18856_ (.A1(\rbzero.pov.ready_buffer[9] ),
    .A2(_02635_),
    .B1(_02690_),
    .C1(_02285_),
    .X(_01068_));
 sky130_fd_sc_hd__or2_1 _18857_ (.A(_01786_),
    .B(_02637_),
    .X(_02691_));
 sky130_fd_sc_hd__o211a_1 _18858_ (.A1(\rbzero.pov.ready_buffer[10] ),
    .A2(_02635_),
    .B1(_02691_),
    .C1(_02285_),
    .X(_01069_));
 sky130_fd_sc_hd__a31o_1 _18859_ (.A1(_02415_),
    .A2(_02414_),
    .A3(_02420_),
    .B1(\rbzero.pov.spi_done ),
    .X(_02692_));
 sky130_fd_sc_hd__and2_1 _18860_ (.A(_02143_),
    .B(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__clkbuf_1 _18861_ (.A(_02693_),
    .X(_01070_));
 sky130_fd_sc_hd__nor2_1 _18862_ (.A(_03852_),
    .B(_04503_),
    .Y(_02694_));
 sky130_fd_sc_hd__nand2_1 _18863_ (.A(_02258_),
    .B(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__or4bb_1 _18864_ (.A(_04500_),
    .B(_04499_),
    .C_N(_04508_),
    .D_N(_04507_),
    .X(_02696_));
 sky130_fd_sc_hd__and4bb_1 _18865_ (.A_N(_04507_),
    .B_N(_04499_),
    .C(_04500_),
    .D(_04508_),
    .X(_02697_));
 sky130_fd_sc_hd__a31o_1 _18866_ (.A1(_02258_),
    .A2(_02694_),
    .A3(_02697_),
    .B1(\rbzero.vga_sync.vsync ),
    .X(_02698_));
 sky130_fd_sc_hd__o211a_1 _18867_ (.A1(_02695_),
    .A2(_02696_),
    .B1(_02698_),
    .C1(_02285_),
    .X(_01071_));
 sky130_fd_sc_hd__or4_1 _18868_ (.A(_03865_),
    .B(_03459_),
    .C(_02903_),
    .D(_03529_),
    .X(_02699_));
 sky130_fd_sc_hd__and4b_1 _18869_ (.A_N(_02699_),
    .B(_03474_),
    .C(_03462_),
    .D(_03505_),
    .X(_02700_));
 sky130_fd_sc_hd__o41a_1 _18870_ (.A1(_04020_),
    .A2(_03464_),
    .A3(_04046_),
    .A4(_02699_),
    .B1(_02334_),
    .X(_02701_));
 sky130_fd_sc_hd__o21a_1 _18871_ (.A1(\rbzero.hsync ),
    .A2(_02700_),
    .B1(_02701_),
    .X(_01072_));
 sky130_fd_sc_hd__or4b_1 _18872_ (.A(_03906_),
    .B(_03531_),
    .C(_02696_),
    .D_N(_03909_),
    .X(_02702_));
 sky130_fd_sc_hd__a21o_1 _18873_ (.A1(_03506_),
    .A2(_02702_),
    .B1(_04499_),
    .X(_02703_));
 sky130_fd_sc_hd__and3b_1 _18874_ (.A_N(_02286_),
    .B(_02703_),
    .C(_04834_),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_1 _18875_ (.A(_02704_),
    .X(_01073_));
 sky130_fd_sc_hd__nand2_1 _18876_ (.A(_04500_),
    .B(_02286_),
    .Y(_02705_));
 sky130_fd_sc_hd__o211a_1 _18877_ (.A1(_04500_),
    .A2(_02286_),
    .B1(_02705_),
    .C1(_02285_),
    .X(_01074_));
 sky130_fd_sc_hd__a31o_1 _18878_ (.A1(_04500_),
    .A2(_04499_),
    .A3(_02279_),
    .B1(_04507_),
    .X(_02706_));
 sky130_fd_sc_hd__a21o_1 _18879_ (.A1(_04827_),
    .A2(_02702_),
    .B1(_08439_),
    .X(_02707_));
 sky130_fd_sc_hd__and3b_1 _18880_ (.A_N(_02287_),
    .B(_02706_),
    .C(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__clkbuf_1 _18881_ (.A(_02708_),
    .X(_01075_));
 sky130_fd_sc_hd__buf_4 _18882_ (.A(_08439_),
    .X(_02709_));
 sky130_fd_sc_hd__a31o_1 _18883_ (.A1(_04507_),
    .A2(_04500_),
    .A3(_04499_),
    .B1(_04508_),
    .X(_02710_));
 sky130_fd_sc_hd__and4b_1 _18884_ (.A_N(_02259_),
    .B(_02702_),
    .C(_02710_),
    .D(_02279_),
    .X(_02711_));
 sky130_fd_sc_hd__a22o_1 _18885_ (.A1(_04508_),
    .A2(_02709_),
    .B1(_02711_),
    .B2(_02285_),
    .X(_01076_));
 sky130_fd_sc_hd__o211a_1 _18886_ (.A1(_04503_),
    .A2(_02280_),
    .B1(_02281_),
    .C1(_02285_),
    .X(_01077_));
 sky130_fd_sc_hd__and3_1 _18887_ (.A(_03902_),
    .B(_04503_),
    .C(_02280_),
    .X(_02712_));
 sky130_fd_sc_hd__inv_2 _18888_ (.A(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__o211a_1 _18889_ (.A1(_03902_),
    .A2(_02260_),
    .B1(_02713_),
    .C1(_02285_),
    .X(_01078_));
 sky130_fd_sc_hd__and3_1 _18890_ (.A(_03520_),
    .B(_03902_),
    .C(_02260_),
    .X(_02714_));
 sky130_fd_sc_hd__or2_1 _18891_ (.A(_03520_),
    .B(_02712_),
    .X(_02715_));
 sky130_fd_sc_hd__and3b_1 _18892_ (.A_N(_02714_),
    .B(_04834_),
    .C(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__clkbuf_1 _18893_ (.A(_02716_),
    .X(_01079_));
 sky130_fd_sc_hd__o21a_1 _18894_ (.A1(_03515_),
    .A2(_02714_),
    .B1(_02323_),
    .X(_02717_));
 sky130_fd_sc_hd__o21a_1 _18895_ (.A1(_03907_),
    .A2(_02713_),
    .B1(_02717_),
    .X(_01080_));
 sky130_fd_sc_hd__a21o_1 _18896_ (.A1(_03515_),
    .A2(_02714_),
    .B1(_03906_),
    .X(_02718_));
 sky130_fd_sc_hd__or3_1 _18897_ (.A(_02257_),
    .B(_03907_),
    .C(_02713_),
    .X(_02719_));
 sky130_fd_sc_hd__and3_1 _18898_ (.A(_02334_),
    .B(_02718_),
    .C(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_1 _18899_ (.A(_02720_),
    .X(_01081_));
 sky130_fd_sc_hd__xnor2_1 _18900_ (.A(_03909_),
    .B(_02719_),
    .Y(_02721_));
 sky130_fd_sc_hd__and2_1 _18901_ (.A(_02707_),
    .B(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__clkbuf_1 _18902_ (.A(_02722_),
    .X(_01082_));
 sky130_fd_sc_hd__a31o_1 _18903_ (.A1(\rbzero.spi_registers.got_new_mapd ),
    .A2(_02323_),
    .A3(_02283_),
    .B1(_01663_),
    .X(_01083_));
 sky130_fd_sc_hd__inv_2 _18905__92 (.A(clknet_1_1__leaf__02441_),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _18906__93 (.A(clknet_1_1__leaf__02441_),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _18907__94 (.A(clknet_1_0__leaf__02441_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _18908__95 (.A(clknet_1_0__leaf__02441_),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _18909__96 (.A(clknet_1_0__leaf__02441_),
    .Y(net218));
 sky130_fd_sc_hd__inv_2 _18911__97 (.A(clknet_1_1__leaf__02723_),
    .Y(net219));
 sky130_fd_sc_hd__buf_1 _18910_ (.A(clknet_1_0__leaf__02440_),
    .X(_02723_));
 sky130_fd_sc_hd__inv_2 _18912__98 (.A(clknet_1_1__leaf__02723_),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _18913__99 (.A(clknet_1_1__leaf__02723_),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _18914__100 (.A(clknet_1_1__leaf__02723_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _18915__101 (.A(clknet_1_0__leaf__02723_),
    .Y(net223));
 sky130_fd_sc_hd__inv_2 _18916__102 (.A(clknet_1_0__leaf__02723_),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _18917__103 (.A(clknet_1_0__leaf__02723_),
    .Y(net225));
 sky130_fd_sc_hd__inv_2 _18918__104 (.A(clknet_1_0__leaf__02723_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _18919__105 (.A(clknet_1_0__leaf__02723_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _18920__106 (.A(clknet_1_0__leaf__02723_),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _18922__107 (.A(clknet_1_0__leaf__02724_),
    .Y(net229));
 sky130_fd_sc_hd__buf_1 _18921_ (.A(clknet_1_0__leaf__02440_),
    .X(_02724_));
 sky130_fd_sc_hd__inv_2 _18923__108 (.A(clknet_1_0__leaf__02724_),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _18924__109 (.A(clknet_1_0__leaf__02724_),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _18925__110 (.A(clknet_1_0__leaf__02724_),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _18926__111 (.A(clknet_1_0__leaf__02724_),
    .Y(net233));
 sky130_fd_sc_hd__inv_2 _18927__112 (.A(clknet_1_1__leaf__02724_),
    .Y(net234));
 sky130_fd_sc_hd__inv_2 _18928__113 (.A(clknet_1_1__leaf__02724_),
    .Y(net235));
 sky130_fd_sc_hd__inv_2 _18929__114 (.A(clknet_1_1__leaf__02724_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _18930__115 (.A(clknet_1_1__leaf__02724_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _18931__116 (.A(clknet_1_1__leaf__02724_),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _18933__117 (.A(clknet_1_0__leaf__02725_),
    .Y(net239));
 sky130_fd_sc_hd__buf_1 _18932_ (.A(clknet_1_0__leaf__02440_),
    .X(_02725_));
 sky130_fd_sc_hd__inv_2 _18934__118 (.A(clknet_1_1__leaf__02725_),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _18935__119 (.A(clknet_1_1__leaf__02725_),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _18936__120 (.A(clknet_1_1__leaf__02725_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _18937__121 (.A(clknet_1_1__leaf__02725_),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _18938__122 (.A(clknet_1_0__leaf__02725_),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _18939__123 (.A(clknet_1_0__leaf__02725_),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _18940__124 (.A(clknet_1_0__leaf__02725_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _18941__125 (.A(clknet_1_0__leaf__02725_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _18942__126 (.A(clknet_1_0__leaf__02725_),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _18944__127 (.A(clknet_1_0__leaf__02726_),
    .Y(net249));
 sky130_fd_sc_hd__buf_1 _18943_ (.A(clknet_1_1__leaf__02440_),
    .X(_02726_));
 sky130_fd_sc_hd__inv_2 _18945__128 (.A(clknet_1_0__leaf__02726_),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _18946__129 (.A(clknet_1_0__leaf__02726_),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _18947__130 (.A(clknet_1_1__leaf__02726_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _18948__131 (.A(clknet_1_1__leaf__02726_),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _18949__132 (.A(clknet_1_1__leaf__02726_),
    .Y(net254));
 sky130_fd_sc_hd__inv_2 _18950__133 (.A(clknet_1_1__leaf__02726_),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _18951__134 (.A(clknet_1_1__leaf__02726_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _18952__135 (.A(clknet_1_1__leaf__02726_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _18953__136 (.A(clknet_1_0__leaf__02726_),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _18955__137 (.A(clknet_1_0__leaf__02727_),
    .Y(net259));
 sky130_fd_sc_hd__buf_1 _18954_ (.A(clknet_1_1__leaf__02440_),
    .X(_02727_));
 sky130_fd_sc_hd__inv_2 _18956__138 (.A(clknet_1_0__leaf__02727_),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _18957__139 (.A(clknet_1_0__leaf__02727_),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _18958__140 (.A(clknet_1_0__leaf__02727_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _18959__141 (.A(clknet_1_1__leaf__02727_),
    .Y(net263));
 sky130_fd_sc_hd__inv_2 _18960__142 (.A(clknet_1_1__leaf__02727_),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _18961__143 (.A(clknet_1_1__leaf__02727_),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _18962__144 (.A(clknet_1_1__leaf__02727_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _18963__145 (.A(clknet_1_1__leaf__02727_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _18964__146 (.A(clknet_1_0__leaf__02727_),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _18966__147 (.A(clknet_1_0__leaf__02728_),
    .Y(net269));
 sky130_fd_sc_hd__buf_1 _18965_ (.A(clknet_1_1__leaf__02440_),
    .X(_02728_));
 sky130_fd_sc_hd__inv_2 _18967__148 (.A(clknet_1_1__leaf__02728_),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _18968__149 (.A(clknet_1_1__leaf__02728_),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _18969__150 (.A(clknet_1_1__leaf__02728_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _18970__151 (.A(clknet_1_1__leaf__02728_),
    .Y(net273));
 sky130_fd_sc_hd__inv_2 _18971__152 (.A(clknet_1_0__leaf__02728_),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _18972__153 (.A(clknet_1_0__leaf__02728_),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _18973__154 (.A(clknet_1_0__leaf__02728_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _18974__155 (.A(clknet_1_1__leaf__02728_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _18975__156 (.A(clknet_1_1__leaf__02728_),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _18977__157 (.A(clknet_1_1__leaf__02729_),
    .Y(net279));
 sky130_fd_sc_hd__buf_1 _18976_ (.A(clknet_1_1__leaf__02440_),
    .X(_02729_));
 sky130_fd_sc_hd__inv_2 _18978__158 (.A(clknet_1_1__leaf__02729_),
    .Y(net280));
 sky130_fd_sc_hd__inv_2 _18979__159 (.A(clknet_1_1__leaf__02729_),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _18980__160 (.A(clknet_1_1__leaf__02729_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _18981__161 (.A(clknet_1_1__leaf__02729_),
    .Y(net283));
 sky130_fd_sc_hd__inv_2 _18982__162 (.A(clknet_1_0__leaf__02729_),
    .Y(net284));
 sky130_fd_sc_hd__inv_2 _18983__163 (.A(clknet_1_0__leaf__02729_),
    .Y(net285));
 sky130_fd_sc_hd__inv_2 _18984__164 (.A(clknet_1_0__leaf__02729_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _18985__165 (.A(clknet_1_0__leaf__02729_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _18986__166 (.A(clknet_1_0__leaf__02729_),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _18988__167 (.A(clknet_1_0__leaf__02730_),
    .Y(net289));
 sky130_fd_sc_hd__buf_1 _18987_ (.A(clknet_1_1__leaf__02440_),
    .X(_02730_));
 sky130_fd_sc_hd__inv_2 _18989__168 (.A(clknet_1_1__leaf__02730_),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _18990__169 (.A(clknet_1_1__leaf__02730_),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _18991__170 (.A(clknet_1_1__leaf__02730_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _18992__171 (.A(clknet_1_0__leaf__02730_),
    .Y(net293));
 sky130_fd_sc_hd__inv_2 _18993__172 (.A(clknet_1_0__leaf__02730_),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _18994__173 (.A(clknet_1_0__leaf__02730_),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _18995__174 (.A(clknet_1_0__leaf__02730_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _18996__175 (.A(clknet_1_1__leaf__02730_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _18997__176 (.A(clknet_1_1__leaf__02730_),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _18999__177 (.A(clknet_1_1__leaf__02731_),
    .Y(net299));
 sky130_fd_sc_hd__buf_1 _18998_ (.A(clknet_1_1__leaf__02440_),
    .X(_02731_));
 sky130_fd_sc_hd__inv_2 _19000__178 (.A(clknet_1_1__leaf__02731_),
    .Y(net300));
 sky130_fd_sc_hd__inv_2 _19001__179 (.A(clknet_1_1__leaf__02731_),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _19002__180 (.A(clknet_1_1__leaf__02731_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _19003__181 (.A(clknet_1_1__leaf__02731_),
    .Y(net303));
 sky130_fd_sc_hd__inv_2 _19004__182 (.A(clknet_1_0__leaf__02731_),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _19005__183 (.A(clknet_1_0__leaf__02731_),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _19006__184 (.A(clknet_1_0__leaf__02731_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _19007__185 (.A(clknet_1_0__leaf__02731_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _19008__186 (.A(clknet_1_0__leaf__02731_),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _19011__187 (.A(clknet_1_1__leaf__02733_),
    .Y(net309));
 sky130_fd_sc_hd__buf_1 _19009_ (.A(clknet_1_1__leaf__04486_),
    .X(_02732_));
 sky130_fd_sc_hd__buf_1 _19010_ (.A(clknet_1_1__leaf__02732_),
    .X(_02733_));
 sky130_fd_sc_hd__inv_2 _19012__188 (.A(clknet_1_1__leaf__02733_),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 _19013__189 (.A(clknet_1_1__leaf__02733_),
    .Y(net311));
 sky130_fd_sc_hd__inv_2 _19014__190 (.A(clknet_1_1__leaf__02733_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _19015__191 (.A(clknet_1_1__leaf__02733_),
    .Y(net313));
 sky130_fd_sc_hd__inv_2 _19016__192 (.A(clknet_1_1__leaf__02733_),
    .Y(net314));
 sky130_fd_sc_hd__inv_2 _19017__193 (.A(clknet_1_0__leaf__02733_),
    .Y(net315));
 sky130_fd_sc_hd__inv_2 _19018__194 (.A(clknet_1_0__leaf__02733_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _19019__195 (.A(clknet_1_0__leaf__02733_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _19020__196 (.A(clknet_1_0__leaf__02733_),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _19022__197 (.A(clknet_1_1__leaf__02734_),
    .Y(net319));
 sky130_fd_sc_hd__buf_1 _19021_ (.A(clknet_1_1__leaf__02732_),
    .X(_02734_));
 sky130_fd_sc_hd__inv_2 _19023__198 (.A(clknet_1_1__leaf__02734_),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _19024__199 (.A(clknet_1_1__leaf__02734_),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _19025__200 (.A(clknet_1_1__leaf__02734_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _19026__201 (.A(clknet_1_1__leaf__02734_),
    .Y(net323));
 sky130_fd_sc_hd__inv_2 _19027__202 (.A(clknet_1_1__leaf__02734_),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _19028__203 (.A(clknet_1_0__leaf__02734_),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _19029__204 (.A(clknet_1_0__leaf__02734_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _19030__205 (.A(clknet_1_0__leaf__02734_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _19031__206 (.A(clknet_1_0__leaf__02734_),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _19033__207 (.A(clknet_1_1__leaf__02735_),
    .Y(net329));
 sky130_fd_sc_hd__buf_1 _19032_ (.A(clknet_1_1__leaf__02732_),
    .X(_02735_));
 sky130_fd_sc_hd__inv_2 _19034__208 (.A(clknet_1_1__leaf__02735_),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _19035__209 (.A(clknet_1_1__leaf__02735_),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _19036__210 (.A(clknet_1_1__leaf__02735_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _19037__211 (.A(clknet_1_1__leaf__02735_),
    .Y(net333));
 sky130_fd_sc_hd__inv_2 _19038__212 (.A(clknet_1_1__leaf__02735_),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _19039__213 (.A(clknet_1_0__leaf__02735_),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _19040__214 (.A(clknet_1_0__leaf__02735_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _19041__215 (.A(clknet_1_0__leaf__02735_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _19042__216 (.A(clknet_1_0__leaf__02735_),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _19044__217 (.A(clknet_1_0__leaf__02736_),
    .Y(net339));
 sky130_fd_sc_hd__buf_1 _19043_ (.A(clknet_1_0__leaf__02732_),
    .X(_02736_));
 sky130_fd_sc_hd__inv_2 _19045__218 (.A(clknet_1_0__leaf__02736_),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _19046__219 (.A(clknet_1_1__leaf__02736_),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _19047__220 (.A(clknet_1_1__leaf__02736_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _19048__221 (.A(clknet_1_1__leaf__02736_),
    .Y(net343));
 sky130_fd_sc_hd__inv_2 _19049__222 (.A(clknet_1_1__leaf__02736_),
    .Y(net344));
 sky130_fd_sc_hd__inv_2 _19050__223 (.A(clknet_1_1__leaf__02736_),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _19051__224 (.A(clknet_1_1__leaf__02736_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _19052__225 (.A(clknet_1_0__leaf__02736_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _19053__226 (.A(clknet_1_0__leaf__02736_),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _19055__227 (.A(clknet_1_1__leaf__02737_),
    .Y(net349));
 sky130_fd_sc_hd__buf_1 _19054_ (.A(clknet_1_0__leaf__02732_),
    .X(_02737_));
 sky130_fd_sc_hd__inv_2 _19056__228 (.A(clknet_1_1__leaf__02737_),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _19057__229 (.A(clknet_1_1__leaf__02737_),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _19058__230 (.A(clknet_1_1__leaf__02737_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _19059__231 (.A(clknet_1_0__leaf__02737_),
    .Y(net353));
 sky130_fd_sc_hd__inv_2 _19060__232 (.A(clknet_1_0__leaf__02737_),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _19061__233 (.A(clknet_1_1__leaf__02737_),
    .Y(net355));
 sky130_fd_sc_hd__inv_2 _19062__234 (.A(clknet_1_0__leaf__02737_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _19063__235 (.A(clknet_1_0__leaf__02737_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _19064__236 (.A(clknet_1_0__leaf__02737_),
    .Y(net358));
 sky130_fd_sc_hd__inv_2 _19066__237 (.A(clknet_1_1__leaf__02738_),
    .Y(net359));
 sky130_fd_sc_hd__buf_1 _19065_ (.A(clknet_1_0__leaf__02732_),
    .X(_02738_));
 sky130_fd_sc_hd__inv_2 _19067__238 (.A(clknet_1_1__leaf__02738_),
    .Y(net360));
 sky130_fd_sc_hd__inv_2 _19068__239 (.A(clknet_1_0__leaf__02738_),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 _19069__240 (.A(clknet_1_0__leaf__02738_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _19070__241 (.A(clknet_1_0__leaf__02738_),
    .Y(net363));
 sky130_fd_sc_hd__inv_2 _19071__242 (.A(clknet_1_0__leaf__02738_),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _19072__243 (.A(clknet_1_0__leaf__02738_),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _19073__244 (.A(clknet_1_1__leaf__02738_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _19074__245 (.A(clknet_1_1__leaf__02738_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _19075__246 (.A(clknet_1_1__leaf__02738_),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _19077__247 (.A(clknet_1_1__leaf__02739_),
    .Y(net369));
 sky130_fd_sc_hd__buf_1 _19076_ (.A(clknet_1_0__leaf__02732_),
    .X(_02739_));
 sky130_fd_sc_hd__inv_2 _19078__248 (.A(clknet_1_1__leaf__02739_),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _19079__249 (.A(clknet_1_1__leaf__02739_),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _19080__250 (.A(clknet_1_0__leaf__02739_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _19081__251 (.A(clknet_1_0__leaf__02739_),
    .Y(net373));
 sky130_fd_sc_hd__inv_2 _19082__252 (.A(clknet_1_0__leaf__02739_),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _19083__253 (.A(clknet_1_0__leaf__02739_),
    .Y(net375));
 sky130_fd_sc_hd__inv_2 _19084__254 (.A(clknet_1_0__leaf__02739_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _19085__255 (.A(clknet_1_1__leaf__02739_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _19086__256 (.A(clknet_1_1__leaf__02739_),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _19088__257 (.A(clknet_1_1__leaf__02740_),
    .Y(net379));
 sky130_fd_sc_hd__buf_1 _19087_ (.A(clknet_1_1__leaf__02732_),
    .X(_02740_));
 sky130_fd_sc_hd__inv_2 _19089__258 (.A(clknet_1_1__leaf__02740_),
    .Y(net380));
 sky130_fd_sc_hd__inv_2 _19090__259 (.A(clknet_1_0__leaf__02740_),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _19091__260 (.A(clknet_1_0__leaf__02740_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _19092__261 (.A(clknet_1_0__leaf__02740_),
    .Y(net383));
 sky130_fd_sc_hd__inv_2 _19093__262 (.A(clknet_1_0__leaf__02740_),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _19094__263 (.A(clknet_1_0__leaf__02740_),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _19095__264 (.A(clknet_1_1__leaf__02740_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _19096__265 (.A(clknet_1_1__leaf__02740_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _19097__266 (.A(clknet_1_1__leaf__02740_),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _19099__267 (.A(clknet_1_1__leaf__02741_),
    .Y(net389));
 sky130_fd_sc_hd__buf_1 _19098_ (.A(clknet_1_0__leaf__02732_),
    .X(_02741_));
 sky130_fd_sc_hd__inv_2 _19100__268 (.A(clknet_1_0__leaf__02741_),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _19101__269 (.A(clknet_1_0__leaf__02741_),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _19102__270 (.A(clknet_1_0__leaf__02741_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _19103__271 (.A(clknet_1_0__leaf__02741_),
    .Y(net393));
 sky130_fd_sc_hd__inv_2 _19104__272 (.A(clknet_1_0__leaf__02741_),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _19105__273 (.A(clknet_1_0__leaf__02741_),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _19106__274 (.A(clknet_1_1__leaf__02741_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _19107__275 (.A(clknet_1_1__leaf__02741_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _19108__276 (.A(clknet_1_1__leaf__02741_),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _19110__277 (.A(clknet_1_0__leaf__02742_),
    .Y(net399));
 sky130_fd_sc_hd__buf_1 _19109_ (.A(clknet_1_0__leaf__02732_),
    .X(_02742_));
 sky130_fd_sc_hd__inv_2 _19111__278 (.A(clknet_1_0__leaf__02742_),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _19112__279 (.A(clknet_1_0__leaf__02742_),
    .Y(net401));
 sky130_fd_sc_hd__inv_2 _19113__280 (.A(clknet_1_0__leaf__02742_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _19114__281 (.A(clknet_1_0__leaf__02742_),
    .Y(net403));
 sky130_fd_sc_hd__inv_2 _19115__282 (.A(clknet_1_0__leaf__02742_),
    .Y(net404));
 sky130_fd_sc_hd__inv_2 _19116__283 (.A(clknet_1_1__leaf__02742_),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _19117__284 (.A(clknet_1_1__leaf__02742_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _19118__285 (.A(clknet_1_1__leaf__02742_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _19119__286 (.A(clknet_1_1__leaf__02742_),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _19122__287 (.A(clknet_1_0__leaf__02744_),
    .Y(net409));
 sky130_fd_sc_hd__buf_1 _19120_ (.A(clknet_1_1__leaf__04486_),
    .X(_02743_));
 sky130_fd_sc_hd__buf_1 _19121_ (.A(clknet_1_1__leaf__02743_),
    .X(_02744_));
 sky130_fd_sc_hd__inv_2 _19123__288 (.A(clknet_1_0__leaf__02744_),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _19124__289 (.A(clknet_1_0__leaf__02744_),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _19125__290 (.A(clknet_1_0__leaf__02744_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _19126__291 (.A(clknet_1_0__leaf__02744_),
    .Y(net413));
 sky130_fd_sc_hd__inv_2 _19127__292 (.A(clknet_1_0__leaf__02744_),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _19128__293 (.A(clknet_1_1__leaf__02744_),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _19129__294 (.A(clknet_1_1__leaf__02744_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _19130__295 (.A(clknet_1_1__leaf__02744_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _19131__296 (.A(clknet_1_1__leaf__02744_),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _19133__297 (.A(clknet_1_0__leaf__02745_),
    .Y(net419));
 sky130_fd_sc_hd__buf_1 _19132_ (.A(clknet_1_1__leaf__02743_),
    .X(_02745_));
 sky130_fd_sc_hd__inv_2 _19134__298 (.A(clknet_1_0__leaf__02745_),
    .Y(net420));
 sky130_fd_sc_hd__inv_2 _19135__299 (.A(clknet_1_0__leaf__02745_),
    .Y(net421));
 sky130_fd_sc_hd__inv_2 _19136__300 (.A(clknet_1_0__leaf__02745_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _19137__301 (.A(clknet_1_0__leaf__02745_),
    .Y(net423));
 sky130_fd_sc_hd__inv_2 _19138__302 (.A(clknet_1_1__leaf__02745_),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _19139__303 (.A(clknet_1_1__leaf__02745_),
    .Y(net425));
 sky130_fd_sc_hd__inv_2 _19140__304 (.A(clknet_1_1__leaf__02745_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _19141__305 (.A(clknet_1_1__leaf__02745_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _19142__306 (.A(clknet_1_1__leaf__02745_),
    .Y(net428));
 sky130_fd_sc_hd__inv_2 _19144__307 (.A(clknet_1_1__leaf__02746_),
    .Y(net429));
 sky130_fd_sc_hd__buf_1 _19143_ (.A(clknet_1_1__leaf__02743_),
    .X(_02746_));
 sky130_fd_sc_hd__inv_2 _19145__308 (.A(clknet_1_1__leaf__02746_),
    .Y(net430));
 sky130_fd_sc_hd__inv_2 _19146__309 (.A(clknet_1_1__leaf__02746_),
    .Y(net431));
 sky130_fd_sc_hd__inv_2 _19147__310 (.A(clknet_1_1__leaf__02746_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _19148__311 (.A(clknet_1_1__leaf__02746_),
    .Y(net433));
 sky130_fd_sc_hd__inv_2 _19149__312 (.A(clknet_1_1__leaf__02746_),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _19150__313 (.A(clknet_1_0__leaf__02746_),
    .Y(net435));
 sky130_fd_sc_hd__inv_2 _19151__314 (.A(clknet_1_0__leaf__02746_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _19152__315 (.A(clknet_1_0__leaf__02746_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _19153__316 (.A(clknet_1_0__leaf__02746_),
    .Y(net438));
 sky130_fd_sc_hd__inv_2 _19155__317 (.A(clknet_1_1__leaf__02747_),
    .Y(net439));
 sky130_fd_sc_hd__buf_1 _19154_ (.A(clknet_1_1__leaf__02743_),
    .X(_02747_));
 sky130_fd_sc_hd__inv_2 _19156__318 (.A(clknet_1_1__leaf__02747_),
    .Y(net440));
 sky130_fd_sc_hd__inv_2 _19157__319 (.A(clknet_1_0__leaf__02747_),
    .Y(net441));
 sky130_fd_sc_hd__inv_2 _19158__320 (.A(clknet_1_0__leaf__02747_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _19159__321 (.A(clknet_1_0__leaf__02747_),
    .Y(net443));
 sky130_fd_sc_hd__inv_2 _19160__322 (.A(clknet_1_0__leaf__02747_),
    .Y(net444));
 sky130_fd_sc_hd__inv_2 _19161__323 (.A(clknet_1_0__leaf__02747_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _19162__324 (.A(clknet_1_1__leaf__02747_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _19163__325 (.A(clknet_1_1__leaf__02747_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _19164__326 (.A(clknet_1_1__leaf__02747_),
    .Y(net448));
 sky130_fd_sc_hd__inv_2 _19166__327 (.A(clknet_1_0__leaf__02748_),
    .Y(net449));
 sky130_fd_sc_hd__buf_1 _19165_ (.A(clknet_1_1__leaf__02743_),
    .X(_02748_));
 sky130_fd_sc_hd__inv_2 _19167__328 (.A(clknet_1_0__leaf__02748_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _19168__329 (.A(clknet_1_1__leaf__02748_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _19169__330 (.A(clknet_1_1__leaf__02748_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _19170__331 (.A(clknet_1_0__leaf__02748_),
    .Y(net453));
 sky130_fd_sc_hd__inv_2 _19171__332 (.A(clknet_1_0__leaf__02748_),
    .Y(net454));
 sky130_fd_sc_hd__inv_2 _19172__333 (.A(clknet_1_0__leaf__02748_),
    .Y(net455));
 sky130_fd_sc_hd__inv_2 _19173__334 (.A(clknet_1_1__leaf__02748_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _19174__335 (.A(clknet_1_1__leaf__02748_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _19175__336 (.A(clknet_1_1__leaf__02748_),
    .Y(net458));
 sky130_fd_sc_hd__inv_2 _19177__337 (.A(clknet_1_1__leaf__02749_),
    .Y(net459));
 sky130_fd_sc_hd__buf_1 _19176_ (.A(clknet_1_1__leaf__02743_),
    .X(_02749_));
 sky130_fd_sc_hd__inv_2 _19178__338 (.A(clknet_1_1__leaf__02749_),
    .Y(net460));
 sky130_fd_sc_hd__inv_2 _19179__339 (.A(clknet_1_1__leaf__02749_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _19180__340 (.A(clknet_1_1__leaf__02749_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _19181__341 (.A(clknet_1_1__leaf__02749_),
    .Y(net463));
 sky130_fd_sc_hd__inv_2 _19182__342 (.A(clknet_1_0__leaf__02749_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _19183__343 (.A(clknet_1_0__leaf__02749_),
    .Y(net465));
 sky130_fd_sc_hd__inv_2 _19184__344 (.A(clknet_1_0__leaf__02749_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _19185__345 (.A(clknet_1_0__leaf__02749_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _19186__346 (.A(clknet_1_0__leaf__02749_),
    .Y(net468));
 sky130_fd_sc_hd__inv_2 _19188__347 (.A(clknet_1_1__leaf__02750_),
    .Y(net469));
 sky130_fd_sc_hd__buf_1 _19187_ (.A(clknet_1_0__leaf__02743_),
    .X(_02750_));
 sky130_fd_sc_hd__inv_2 _19189__348 (.A(clknet_1_1__leaf__02750_),
    .Y(net470));
 sky130_fd_sc_hd__inv_2 _19190__349 (.A(clknet_1_1__leaf__02750_),
    .Y(net471));
 sky130_fd_sc_hd__inv_2 _19191__350 (.A(clknet_1_1__leaf__02750_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _19192__351 (.A(clknet_1_1__leaf__02750_),
    .Y(net473));
 sky130_fd_sc_hd__inv_2 _19193__352 (.A(clknet_1_1__leaf__02750_),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _19194__353 (.A(clknet_1_0__leaf__02750_),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _19195__354 (.A(clknet_1_0__leaf__02750_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _19196__355 (.A(clknet_1_0__leaf__02750_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _19197__356 (.A(clknet_1_0__leaf__02750_),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _19199__357 (.A(clknet_1_0__leaf__02751_),
    .Y(net479));
 sky130_fd_sc_hd__buf_1 _19198_ (.A(clknet_1_0__leaf__02743_),
    .X(_02751_));
 sky130_fd_sc_hd__inv_2 _19200__358 (.A(clknet_1_0__leaf__02751_),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _19201__359 (.A(clknet_1_0__leaf__02751_),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _19202__360 (.A(clknet_1_0__leaf__02751_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _19203__361 (.A(clknet_1_0__leaf__02751_),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _19204__362 (.A(clknet_1_1__leaf__02751_),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _19205__363 (.A(clknet_1_1__leaf__02751_),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _19206__364 (.A(clknet_1_1__leaf__02751_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _19207__365 (.A(clknet_1_1__leaf__02751_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _19208__366 (.A(clknet_1_1__leaf__02751_),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _19210__367 (.A(clknet_1_0__leaf__02752_),
    .Y(net489));
 sky130_fd_sc_hd__buf_1 _19209_ (.A(clknet_1_0__leaf__02743_),
    .X(_02752_));
 sky130_fd_sc_hd__inv_2 _19211__368 (.A(clknet_1_0__leaf__02752_),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _19212__369 (.A(clknet_1_0__leaf__02752_),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _19213__370 (.A(clknet_1_0__leaf__02752_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _19214__371 (.A(clknet_1_1__leaf__02752_),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _19215__372 (.A(clknet_1_1__leaf__02752_),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _19216__373 (.A(clknet_1_1__leaf__02752_),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _19217__374 (.A(clknet_1_1__leaf__02752_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _19218__375 (.A(clknet_1_1__leaf__02752_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _19219__376 (.A(clknet_1_1__leaf__02752_),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _19221__377 (.A(clknet_1_0__leaf__02753_),
    .Y(net499));
 sky130_fd_sc_hd__buf_1 _19220_ (.A(clknet_1_0__leaf__02743_),
    .X(_02753_));
 sky130_fd_sc_hd__inv_2 _19222__378 (.A(clknet_1_0__leaf__02753_),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _19223__379 (.A(clknet_1_0__leaf__02753_),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _19224__380 (.A(clknet_1_1__leaf__02753_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _19225__381 (.A(clknet_1_1__leaf__02753_),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _19226__382 (.A(clknet_1_1__leaf__02753_),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _19227__383 (.A(clknet_1_1__leaf__02753_),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _19228__384 (.A(clknet_1_0__leaf__02753_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _19229__385 (.A(clknet_1_0__leaf__02753_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _19230__386 (.A(clknet_1_0__leaf__02753_),
    .Y(net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__buf_1 _19231_ (.A(clknet_1_1__leaf__04486_),
    .X(_02754_));
 sky130_fd_sc_hd__inv_2 _19233__8 (.A(clknet_1_1__leaf__02754_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _19234__9 (.A(clknet_1_1__leaf__02754_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _19235__10 (.A(clknet_1_1__leaf__02754_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _19236__11 (.A(clknet_1_1__leaf__02754_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _19237__12 (.A(clknet_1_0__leaf__02754_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _19238__13 (.A(clknet_1_0__leaf__02754_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _19239__14 (.A(clknet_1_0__leaf__02754_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _19240__15 (.A(clknet_1_0__leaf__02754_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _19241__16 (.A(clknet_1_0__leaf__02754_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _19243__17 (.A(clknet_1_0__leaf__02755_),
    .Y(net139));
 sky130_fd_sc_hd__buf_1 _19242_ (.A(clknet_1_0__leaf__04486_),
    .X(_02755_));
 sky130_fd_sc_hd__inv_2 _19244__18 (.A(clknet_1_0__leaf__02755_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _19245__19 (.A(clknet_1_0__leaf__02755_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _19246__20 (.A(clknet_1_0__leaf__02755_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _19247__21 (.A(clknet_1_0__leaf__02755_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _19248__22 (.A(clknet_1_0__leaf__02755_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _19249__23 (.A(clknet_1_1__leaf__02755_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _19250__24 (.A(clknet_1_1__leaf__02755_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _19251__25 (.A(clknet_1_1__leaf__02755_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _19252__26 (.A(clknet_1_1__leaf__02755_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _18383__27 (.A(clknet_1_0__leaf__02434_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _19254__4 (.A(clknet_1_0__leaf__02433_),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _19255__5 (.A(clknet_1_0__leaf__02433_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _19256__6 (.A(clknet_1_0__leaf__02433_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _19232__7 (.A(clknet_1_1__leaf__02754_),
    .Y(net129));
 sky130_fd_sc_hd__nor2_1 _19257_ (.A(\gpout5.clk_div[0] ),
    .B(net61),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _19258_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .Y(_02756_));
 sky130_fd_sc_hd__or2_1 _19259_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .X(_02757_));
 sky130_fd_sc_hd__and3_1 _19260_ (.A(_02334_),
    .B(_02756_),
    .C(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__clkbuf_1 _19261_ (.A(_02758_),
    .X(_01405_));
 sky130_fd_sc_hd__clkbuf_4 _19262_ (.A(_08439_),
    .X(_02759_));
 sky130_fd_sc_hd__nand2_1 _19263_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .Y(_02760_));
 sky130_fd_sc_hd__or2_1 _19264_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .X(_02761_));
 sky130_fd_sc_hd__buf_4 _19265_ (.A(_03338_),
    .X(_02762_));
 sky130_fd_sc_hd__a32o_1 _19266_ (.A1(_02759_),
    .A2(_02760_),
    .A3(_02761_),
    .B1(_02762_),
    .B2(\rbzero.texV[-11] ),
    .X(_01406_));
 sky130_fd_sc_hd__or2_1 _19267_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .X(_02763_));
 sky130_fd_sc_hd__nand2_1 _19268_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_02764_));
 sky130_fd_sc_hd__nand3b_1 _19269_ (.A_N(_02760_),
    .B(_02763_),
    .C(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__a21bo_1 _19270_ (.A1(_02763_),
    .A2(_02764_),
    .B1_N(_02760_),
    .X(_02766_));
 sky130_fd_sc_hd__a32o_1 _19271_ (.A1(_02759_),
    .A2(_02765_),
    .A3(_02766_),
    .B1(_02762_),
    .B2(\rbzero.texV[-10] ),
    .X(_01407_));
 sky130_fd_sc_hd__and2_1 _19272_ (.A(_02764_),
    .B(_02765_),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_1 _19273_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_02768_));
 sky130_fd_sc_hd__nand2_1 _19274_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_02769_));
 sky130_fd_sc_hd__and2b_1 _19275_ (.A_N(_02768_),
    .B(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__xnor2_1 _19276_ (.A(_02767_),
    .B(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__a22o_1 _19277_ (.A1(\rbzero.texV[-9] ),
    .A2(_02675_),
    .B1(_02709_),
    .B2(_02771_),
    .X(_01408_));
 sky130_fd_sc_hd__or2_1 _19278_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .X(_02772_));
 sky130_fd_sc_hd__nand2_1 _19279_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_1 _19280_ (.A(_02772_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__o21ai_1 _19281_ (.A1(_02767_),
    .A2(_02768_),
    .B1(_02769_),
    .Y(_02775_));
 sky130_fd_sc_hd__xnor2_1 _19282_ (.A(_02774_),
    .B(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__a22o_1 _19283_ (.A1(\rbzero.texV[-8] ),
    .A2(_02675_),
    .B1(_02709_),
    .B2(_02776_),
    .X(_01409_));
 sky130_fd_sc_hd__nor2_1 _19284_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .Y(_02777_));
 sky130_fd_sc_hd__and2_1 _19285_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .X(_02778_));
 sky130_fd_sc_hd__a21boi_1 _19286_ (.A1(_02772_),
    .A2(_02775_),
    .B1_N(_02773_),
    .Y(_02779_));
 sky130_fd_sc_hd__o21ai_1 _19287_ (.A1(_02777_),
    .A2(_02778_),
    .B1(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__or3_1 _19288_ (.A(_02777_),
    .B(_02778_),
    .C(_02779_),
    .X(_02781_));
 sky130_fd_sc_hd__a32o_1 _19289_ (.A1(_02759_),
    .A2(_02780_),
    .A3(_02781_),
    .B1(_02762_),
    .B2(\rbzero.texV[-7] ),
    .X(_01410_));
 sky130_fd_sc_hd__xnor2_1 _19290_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_02782_));
 sky130_fd_sc_hd__o21bai_1 _19291_ (.A1(_02777_),
    .A2(_02779_),
    .B1_N(_02778_),
    .Y(_02783_));
 sky130_fd_sc_hd__xnor2_1 _19292_ (.A(_02782_),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__a22o_1 _19293_ (.A1(\rbzero.texV[-6] ),
    .A2(_02675_),
    .B1(_02709_),
    .B2(_02784_),
    .X(_01411_));
 sky130_fd_sc_hd__nor2_1 _19294_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_02785_));
 sky130_fd_sc_hd__and2_1 _19295_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .X(_02786_));
 sky130_fd_sc_hd__a21o_1 _19296_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_02783_),
    .X(_02787_));
 sky130_fd_sc_hd__o21ai_1 _19297_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__or3_1 _19298_ (.A(_02785_),
    .B(_02786_),
    .C(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__o21ai_1 _19299_ (.A1(_02785_),
    .A2(_02786_),
    .B1(_02788_),
    .Y(_02790_));
 sky130_fd_sc_hd__a32o_1 _19300_ (.A1(_02759_),
    .A2(_02789_),
    .A3(_02790_),
    .B1(_02762_),
    .B2(\rbzero.texV[-5] ),
    .X(_01412_));
 sky130_fd_sc_hd__xnor2_1 _19301_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_02791_));
 sky130_fd_sc_hd__o21bai_1 _19302_ (.A1(_02785_),
    .A2(_02788_),
    .B1_N(_02786_),
    .Y(_02792_));
 sky130_fd_sc_hd__xnor2_1 _19303_ (.A(_02791_),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__a22o_1 _19304_ (.A1(\rbzero.texV[-4] ),
    .A2(_02675_),
    .B1(_02709_),
    .B2(_02793_),
    .X(_01413_));
 sky130_fd_sc_hd__nor2_1 _19305_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_02794_));
 sky130_fd_sc_hd__and2_1 _19306_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .X(_02795_));
 sky130_fd_sc_hd__a21o_1 _19307_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_02792_),
    .X(_02796_));
 sky130_fd_sc_hd__o21ai_1 _19308_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_02796_),
    .Y(_02797_));
 sky130_fd_sc_hd__or3_1 _19309_ (.A(_02794_),
    .B(_02795_),
    .C(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__o21ai_1 _19310_ (.A1(_02794_),
    .A2(_02795_),
    .B1(_02797_),
    .Y(_02799_));
 sky130_fd_sc_hd__a32o_1 _19311_ (.A1(_02759_),
    .A2(_02798_),
    .A3(_02799_),
    .B1(_02762_),
    .B2(\rbzero.texV[-3] ),
    .X(_01414_));
 sky130_fd_sc_hd__or2_1 _19312_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .X(_02800_));
 sky130_fd_sc_hd__nand2_1 _19313_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .Y(_02801_));
 sky130_fd_sc_hd__o21bai_1 _19314_ (.A1(_02794_),
    .A2(_02797_),
    .B1_N(_02795_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand3_1 _19315_ (.A(_02800_),
    .B(_02801_),
    .C(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__a21o_1 _19316_ (.A1(_02800_),
    .A2(_02801_),
    .B1(_02802_),
    .X(_02804_));
 sky130_fd_sc_hd__a32o_1 _19317_ (.A1(_02759_),
    .A2(_02803_),
    .A3(_02804_),
    .B1(_02319_),
    .B2(\rbzero.texV[-2] ),
    .X(_01415_));
 sky130_fd_sc_hd__nor2_1 _19318_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .Y(_02805_));
 sky130_fd_sc_hd__and2_1 _19319_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .X(_02806_));
 sky130_fd_sc_hd__or2_1 _19320_ (.A(_02805_),
    .B(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__a21boi_1 _19321_ (.A1(_02800_),
    .A2(_02802_),
    .B1_N(_02801_),
    .Y(_02808_));
 sky130_fd_sc_hd__xor2_1 _19322_ (.A(_02807_),
    .B(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__a22o_1 _19323_ (.A1(\rbzero.texV[-1] ),
    .A2(_02762_),
    .B1(_02709_),
    .B2(_02809_),
    .X(_01416_));
 sky130_fd_sc_hd__nor2_1 _19324_ (.A(_02807_),
    .B(_02808_),
    .Y(_02810_));
 sky130_fd_sc_hd__or2_1 _19325_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .X(_02811_));
 sky130_fd_sc_hd__nand2_1 _19326_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .Y(_02812_));
 sky130_fd_sc_hd__o211a_1 _19327_ (.A1(_02806_),
    .A2(_02810_),
    .B1(_02811_),
    .C1(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__inv_2 _19328_ (.A(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__a211o_1 _19329_ (.A1(_02811_),
    .A2(_02812_),
    .B1(_02806_),
    .C1(_02810_),
    .X(_02815_));
 sky130_fd_sc_hd__a32o_1 _19330_ (.A1(_02759_),
    .A2(_02814_),
    .A3(_02815_),
    .B1(_02319_),
    .B2(\rbzero.texV[0] ),
    .X(_01417_));
 sky130_fd_sc_hd__or2_1 _19331_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .X(_02816_));
 sky130_fd_sc_hd__nand2_1 _19332_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .Y(_02817_));
 sky130_fd_sc_hd__nand2_1 _19333_ (.A(_02812_),
    .B(_02814_),
    .Y(_02818_));
 sky130_fd_sc_hd__and3_1 _19334_ (.A(_02816_),
    .B(_02817_),
    .C(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__inv_2 _19335_ (.A(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__a21o_1 _19336_ (.A1(_02816_),
    .A2(_02817_),
    .B1(_02818_),
    .X(_02821_));
 sky130_fd_sc_hd__a32o_1 _19337_ (.A1(_02759_),
    .A2(_02820_),
    .A3(_02821_),
    .B1(_02319_),
    .B2(\rbzero.texV[1] ),
    .X(_01418_));
 sky130_fd_sc_hd__or2_1 _19338_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .X(_02822_));
 sky130_fd_sc_hd__nand2_1 _19339_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _19340_ (.A(_02817_),
    .B(_02820_),
    .Y(_02824_));
 sky130_fd_sc_hd__and3_1 _19341_ (.A(_02822_),
    .B(_02823_),
    .C(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__inv_2 _19342_ (.A(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__a21o_1 _19343_ (.A1(_02822_),
    .A2(_02823_),
    .B1(_02824_),
    .X(_02827_));
 sky130_fd_sc_hd__a32o_1 _19344_ (.A1(_02759_),
    .A2(_02826_),
    .A3(_02827_),
    .B1(_02319_),
    .B2(\rbzero.texV[2] ),
    .X(_01419_));
 sky130_fd_sc_hd__or2_1 _19345_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .X(_02828_));
 sky130_fd_sc_hd__nand2_1 _19346_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _19347_ (.A(_02823_),
    .B(_02826_),
    .Y(_02830_));
 sky130_fd_sc_hd__and3_1 _19348_ (.A(_02828_),
    .B(_02829_),
    .C(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__inv_2 _19349_ (.A(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21o_1 _19350_ (.A1(_02828_),
    .A2(_02829_),
    .B1(_02830_),
    .X(_02833_));
 sky130_fd_sc_hd__a32o_1 _19351_ (.A1(_02759_),
    .A2(_02832_),
    .A3(_02833_),
    .B1(_02319_),
    .B2(\rbzero.texV[3] ),
    .X(_01420_));
 sky130_fd_sc_hd__or2_1 _19352_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .X(_02834_));
 sky130_fd_sc_hd__nand2_1 _19353_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_1 _19354_ (.A(_02829_),
    .B(_02832_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand3_1 _19355_ (.A(_02834_),
    .B(_02835_),
    .C(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__a21o_1 _19356_ (.A1(_02834_),
    .A2(_02835_),
    .B1(_02836_),
    .X(_02838_));
 sky130_fd_sc_hd__a32o_1 _19357_ (.A1(_08439_),
    .A2(_02837_),
    .A3(_02838_),
    .B1(_02319_),
    .B2(\rbzero.texV[4] ),
    .X(_01421_));
 sky130_fd_sc_hd__a21boi_1 _19358_ (.A1(_02834_),
    .A2(_02836_),
    .B1_N(_02835_),
    .Y(_02839_));
 sky130_fd_sc_hd__nor2_1 _19359_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_02840_));
 sky130_fd_sc_hd__nand2_1 _19360_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_02841_));
 sky130_fd_sc_hd__and2b_1 _19361_ (.A_N(_02840_),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__xnor2_1 _19362_ (.A(_02839_),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__a22o_1 _19363_ (.A1(\rbzero.texV[5] ),
    .A2(_02762_),
    .B1(_02709_),
    .B2(_02843_),
    .X(_01422_));
 sky130_fd_sc_hd__or2_1 _19364_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .X(_02844_));
 sky130_fd_sc_hd__nand2_1 _19365_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _19366_ (.A(_02844_),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__o21ai_1 _19367_ (.A1(_02839_),
    .A2(_02840_),
    .B1(_02841_),
    .Y(_02847_));
 sky130_fd_sc_hd__xnor2_1 _19368_ (.A(_02846_),
    .B(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hd__a22o_1 _19369_ (.A1(\rbzero.texV[6] ),
    .A2(_02762_),
    .B1(_02709_),
    .B2(_02848_),
    .X(_01423_));
 sky130_fd_sc_hd__nor2_1 _19370_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_02849_));
 sky130_fd_sc_hd__nand2_1 _19371_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_02850_));
 sky130_fd_sc_hd__and2b_1 _19372_ (.A_N(_02849_),
    .B(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__a21boi_1 _19373_ (.A1(_02844_),
    .A2(_02847_),
    .B1_N(_02845_),
    .Y(_02852_));
 sky130_fd_sc_hd__xnor2_1 _19374_ (.A(_02851_),
    .B(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__a22o_1 _19375_ (.A1(\rbzero.texV[7] ),
    .A2(_02762_),
    .B1(_02709_),
    .B2(_02853_),
    .X(_01424_));
 sky130_fd_sc_hd__or2_1 _19376_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _19377_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_02855_));
 sky130_fd_sc_hd__o21ai_1 _19378_ (.A1(_02849_),
    .A2(_02852_),
    .B1(_02850_),
    .Y(_02856_));
 sky130_fd_sc_hd__a21o_1 _19379_ (.A1(_02854_),
    .A2(_02855_),
    .B1(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__nand3_1 _19380_ (.A(_02854_),
    .B(_02855_),
    .C(_02856_),
    .Y(_02858_));
 sky130_fd_sc_hd__a32o_1 _19381_ (.A1(_08439_),
    .A2(_02857_),
    .A3(_02858_),
    .B1(_02319_),
    .B2(\rbzero.texV[8] ),
    .X(_01425_));
 sky130_fd_sc_hd__or2_1 _19382_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .X(_02859_));
 sky130_fd_sc_hd__nand2_1 _19383_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_02860_));
 sky130_fd_sc_hd__a21o_1 _19384_ (.A1(\rbzero.traced_texa[8] ),
    .A2(\rbzero.texV[8] ),
    .B1(_02856_),
    .X(_02861_));
 sky130_fd_sc_hd__a22o_1 _19385_ (.A1(_02859_),
    .A2(_02860_),
    .B1(_02861_),
    .B2(_02854_),
    .X(_02862_));
 sky130_fd_sc_hd__nand4_1 _19386_ (.A(_02854_),
    .B(_02859_),
    .C(_02860_),
    .D(_02861_),
    .Y(_02863_));
 sky130_fd_sc_hd__a32o_1 _19387_ (.A1(_08439_),
    .A2(_02862_),
    .A3(_02863_),
    .B1(_02319_),
    .B2(\rbzero.texV[9] ),
    .X(_01426_));
 sky130_fd_sc_hd__xnor2_1 _19388_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_02864_));
 sky130_fd_sc_hd__and3_1 _19389_ (.A(_02860_),
    .B(_02863_),
    .C(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__a21oi_1 _19390_ (.A1(_02860_),
    .A2(_02863_),
    .B1(_02864_),
    .Y(_02866_));
 sky130_fd_sc_hd__nor2_1 _19391_ (.A(_02865_),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__a22o_1 _19392_ (.A1(\rbzero.texV[10] ),
    .A2(_02762_),
    .B1(_02709_),
    .B2(_02867_),
    .X(_01427_));
 sky130_fd_sc_hd__a22o_1 _19393_ (.A1(\rbzero.traced_texVinit[0] ),
    .A2(_08463_),
    .B1(_07815_),
    .B2(_08455_),
    .X(_01428_));
 sky130_fd_sc_hd__a22o_1 _19394_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(_08463_),
    .B1(_07813_),
    .B2(_08455_),
    .X(_01429_));
 sky130_fd_sc_hd__a22o_1 _19395_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(_08463_),
    .B1(_07808_),
    .B2(_01745_),
    .X(_01430_));
 sky130_fd_sc_hd__a22o_1 _19396_ (.A1(\rbzero.traced_texVinit[3] ),
    .A2(_08463_),
    .B1(_07929_),
    .B2(_01745_),
    .X(_01431_));
 sky130_fd_sc_hd__buf_4 _19397_ (.A(_08460_),
    .X(_02868_));
 sky130_fd_sc_hd__a22o_1 _19398_ (.A1(\rbzero.traced_texVinit[4] ),
    .A2(_02868_),
    .B1(_08052_),
    .B2(_01745_),
    .X(_01432_));
 sky130_fd_sc_hd__a22o_1 _19399_ (.A1(\rbzero.traced_texVinit[5] ),
    .A2(_02868_),
    .B1(_08174_),
    .B2(_01745_),
    .X(_01433_));
 sky130_fd_sc_hd__a22o_1 _19400_ (.A1(\rbzero.traced_texVinit[6] ),
    .A2(_02868_),
    .B1(_08303_),
    .B2(_01745_),
    .X(_01434_));
 sky130_fd_sc_hd__a22o_1 _19401_ (.A1(\rbzero.traced_texVinit[7] ),
    .A2(_02868_),
    .B1(_08431_),
    .B2(_01745_),
    .X(_01435_));
 sky130_fd_sc_hd__a22o_1 _19402_ (.A1(\rbzero.traced_texVinit[8] ),
    .A2(_02868_),
    .B1(_08454_),
    .B2(_08716_),
    .X(_01436_));
 sky130_fd_sc_hd__a22o_1 _19403_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(_02868_),
    .B1(_08454_),
    .B2(_08834_),
    .X(_01437_));
 sky130_fd_sc_hd__a22o_1 _19404_ (.A1(\rbzero.traced_texVinit[10] ),
    .A2(_02868_),
    .B1(_08454_),
    .B2(_08958_),
    .X(_01438_));
 sky130_fd_sc_hd__nor2_1 _19405_ (.A(\gpout0.clk_div[0] ),
    .B(net61),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_1 _19406_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .Y(_02869_));
 sky130_fd_sc_hd__or2_1 _19407_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .X(_02870_));
 sky130_fd_sc_hd__and3_1 _19408_ (.A(_02334_),
    .B(_02869_),
    .C(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__clkbuf_1 _19409_ (.A(_02871_),
    .X(_01440_));
 sky130_fd_sc_hd__or2_1 _19410_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_02872_));
 sky130_fd_sc_hd__and3_1 _19411_ (.A(_08452_),
    .B(_01705_),
    .C(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__a21o_1 _19412_ (.A1(\rbzero.wall_tracer.rayAddendY[-9] ),
    .A2(_08449_),
    .B1(_02873_),
    .X(_01441_));
 sky130_fd_sc_hd__nor2_1 _19413_ (.A(_01707_),
    .B(_01706_),
    .Y(_02874_));
 sky130_fd_sc_hd__xnor2_1 _19414_ (.A(_01705_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__a22o_1 _19415_ (.A1(\rbzero.wall_tracer.rayAddendY[-8] ),
    .A2(_02868_),
    .B1(_08454_),
    .B2(_02875_),
    .X(_01442_));
 sky130_fd_sc_hd__and2b_1 _19416_ (.A_N(_01704_),
    .B(_01709_),
    .X(_02876_));
 sky130_fd_sc_hd__xnor2_1 _19417_ (.A(_01708_),
    .B(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__a22o_1 _19418_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_02868_),
    .B1(_08454_),
    .B2(_02877_),
    .X(_01443_));
 sky130_fd_sc_hd__a21oi_1 _19419_ (.A1(_01703_),
    .A2(_01711_),
    .B1(_01710_),
    .Y(_02878_));
 sky130_fd_sc_hd__a31o_1 _19420_ (.A1(_01703_),
    .A2(_01711_),
    .A3(_01710_),
    .B1(_08464_),
    .X(_02879_));
 sky130_fd_sc_hd__a2bb2o_1 _19421_ (.A1_N(_02878_),
    .A2_N(_02879_),
    .B1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B2(_08449_),
    .X(_01444_));
 sky130_fd_sc_hd__or2_1 _19422_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_02880_));
 sky130_fd_sc_hd__and3_1 _19423_ (.A(_08452_),
    .B(_01921_),
    .C(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__a21o_1 _19424_ (.A1(\rbzero.wall_tracer.rayAddendX[-9] ),
    .A2(_08449_),
    .B1(_02881_),
    .X(_01445_));
 sky130_fd_sc_hd__xor2_1 _19425_ (.A(_01921_),
    .B(_01924_),
    .X(_02882_));
 sky130_fd_sc_hd__a22o_1 _19426_ (.A1(\rbzero.wall_tracer.rayAddendX[-8] ),
    .A2(_02868_),
    .B1(_08454_),
    .B2(_02882_),
    .X(_01446_));
 sky130_fd_sc_hd__and2b_1 _19427_ (.A_N(_01920_),
    .B(_01926_),
    .X(_02883_));
 sky130_fd_sc_hd__xnor2_1 _19428_ (.A(_01925_),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__a22o_1 _19429_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_08448_),
    .B1(_08454_),
    .B2(_02884_),
    .X(_01447_));
 sky130_fd_sc_hd__a21oi_1 _19430_ (.A1(_01919_),
    .A2(_01928_),
    .B1(_01927_),
    .Y(_02885_));
 sky130_fd_sc_hd__a31o_1 _19431_ (.A1(_01919_),
    .A2(_01928_),
    .A3(_01927_),
    .B1(_08464_),
    .X(_02886_));
 sky130_fd_sc_hd__a2bb2o_1 _19432_ (.A1_N(_02885_),
    .A2_N(_02886_),
    .B1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B2(_08449_),
    .X(_01448_));
 sky130_fd_sc_hd__nor2_1 _19433_ (.A(\gpout1.clk_div[0] ),
    .B(net61),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_1 _19434_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .Y(_02887_));
 sky130_fd_sc_hd__or2_1 _19435_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .X(_02888_));
 sky130_fd_sc_hd__and3_1 _19436_ (.A(_02334_),
    .B(_02887_),
    .C(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__clkbuf_1 _19437_ (.A(_02889_),
    .X(_01450_));
 sky130_fd_sc_hd__nor2_1 _19438_ (.A(\gpout2.clk_div[0] ),
    .B(net61),
    .Y(_01451_));
 sky130_fd_sc_hd__nand2_1 _19439_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .Y(_02890_));
 sky130_fd_sc_hd__or2_1 _19440_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .X(_02891_));
 sky130_fd_sc_hd__and3_1 _19441_ (.A(_02334_),
    .B(_02890_),
    .C(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__clkbuf_1 _19442_ (.A(_02892_),
    .X(_01452_));
 sky130_fd_sc_hd__nor2_1 _19443_ (.A(\gpout3.clk_div[0] ),
    .B(net61),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_1 _19444_ (.A(\gpout3.clk_div[1] ),
    .B(\gpout3.clk_div[0] ),
    .Y(_02893_));
 sky130_fd_sc_hd__or2_1 _19445_ (.A(\gpout3.clk_div[1] ),
    .B(\gpout3.clk_div[0] ),
    .X(_02894_));
 sky130_fd_sc_hd__and3_1 _19446_ (.A(_02334_),
    .B(_02893_),
    .C(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _19447_ (.A(_02895_),
    .X(_01454_));
 sky130_fd_sc_hd__nor2_1 _19448_ (.A(\gpout4.clk_div[0] ),
    .B(net61),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _19449_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .Y(_02896_));
 sky130_fd_sc_hd__or2_1 _19450_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .X(_02897_));
 sky130_fd_sc_hd__and3_1 _19451_ (.A(_04828_),
    .B(_02896_),
    .C(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_1 _19452_ (.A(_02898_),
    .X(_01456_));
 sky130_fd_sc_hd__dfxtp_1 _19453_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00011_),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19454_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00012_),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19455_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00401_),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19456_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00402_),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19457_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00403_),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19458_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00404_),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19459_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00405_),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19460_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _19461_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _19462_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _19463_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _19464_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _19465_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _19466_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _19467_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00413_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _19468_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00414_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _19469_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00415_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _19470_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00416_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _19471_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00417_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19472_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00418_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19473_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00419_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19474_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00420_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19475_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00421_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19476_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00422_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19477_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00423_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19478_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00424_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19479_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00425_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_2 _19480_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00426_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_2 _19481_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00427_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19482_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00428_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_4 _19483_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00429_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _19484_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00430_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _19485_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00431_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _19486_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00432_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _19487_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00433_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _19488_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00434_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _19489_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _19490_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _19491_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _19492_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _19493_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_4 _19494_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19495_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19496_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19497_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_4 _19498_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_4 _19499_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_4 _19500_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_4 _19501_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_4 _19502_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_4 _19503_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19504_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _19505_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _19506_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _19507_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _19508_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _19509_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _19510_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _19511_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00457_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _19512_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00458_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _19513_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00459_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _19514_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00460_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _19515_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00461_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19516_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00462_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19517_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00463_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19518_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00464_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19519_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00465_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19520_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00466_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19521_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00467_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19522_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00468_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_2 _19523_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00469_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_2 _19524_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00470_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19525_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00471_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19526_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00013_),
    .Q(\rbzero.wall_tracer.state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _19527_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00015_),
    .Q(\rbzero.wall_tracer.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19528_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00000_),
    .Q(\rbzero.wall_tracer.state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _19529_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00001_),
    .Q(\rbzero.wall_tracer.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19530_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00002_),
    .Q(\rbzero.wall_tracer.state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19531_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00003_),
    .Q(\rbzero.wall_tracer.state[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19532_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00004_),
    .Q(\rbzero.wall_tracer.state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19533_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00005_),
    .Q(\rbzero.wall_tracer.state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19534_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00016_),
    .Q(\rbzero.wall_tracer.state[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19535_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00006_),
    .Q(\rbzero.wall_tracer.state[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19536_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00007_),
    .Q(\rbzero.wall_tracer.state[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19537_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00008_),
    .Q(\rbzero.wall_tracer.state[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19538_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00009_),
    .Q(\rbzero.wall_tracer.state[12] ));
 sky130_fd_sc_hd__dfxtp_2 _19539_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00010_),
    .Q(\rbzero.wall_tracer.state[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19540_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00014_),
    .Q(\rbzero.wall_tracer.state[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19541_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00472_),
    .Q(\rbzero.wall_tracer.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19542_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00473_),
    .Q(\rbzero.wall_tracer.wall[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19543_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00474_),
    .Q(\rbzero.wall_tracer.side ));
 sky130_fd_sc_hd__dfxtp_1 _19544_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00475_),
    .Q(\rbzero.wall_tracer.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19545_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00476_),
    .Q(\rbzero.wall_tracer.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19546_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00477_),
    .Q(\rbzero.wall_tracer.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19547_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00478_),
    .Q(\rbzero.wall_tracer.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19548_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00479_),
    .Q(\rbzero.wall_tracer.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19549_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00480_),
    .Q(\rbzero.wall_tracer.texu[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19550_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00481_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19551_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00482_),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19552_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00483_),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19553_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00484_),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19554_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00485_),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19555_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00486_),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19556_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00487_),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19557_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00488_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19558_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00489_),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_2 _19559_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00490_),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_4 _19560_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00491_),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _19561_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00492_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19562_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00493_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19563_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00494_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19564_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00495_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19565_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00496_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19566_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00497_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19567_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00498_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_2 _19568_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00499_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19569_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00500_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19570_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00501_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19571_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00502_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_2 _19572_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00503_),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19573_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00504_),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19574_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00505_),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_2 _19575_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00506_),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19576_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00507_),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19577_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00508_),
    .Q(\rbzero.row_render.texu[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19578_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00509_),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _19579_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00510_),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _19580_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00511_),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _19581_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00512_),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _19582_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00513_),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _19583_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00514_),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _19584_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00515_),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _19585_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00516_),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _19586_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00517_),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _19587_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00518_),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _19588_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00519_),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _19589_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00520_),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19590_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00521_),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19591_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00522_),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19592_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00523_),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19593_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00524_),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19594_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00525_),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19595_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00526_),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19596_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00527_),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19597_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00528_),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19598_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00529_),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19599_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00530_),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_2 _19600_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00531_),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19601_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00532_),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19602_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00533_),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19603_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00534_),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19604_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00535_),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19605_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00536_),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19606_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00537_),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19607_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00538_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _19608_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00539_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _19609_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00540_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _19610_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _19611_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _19612_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _19613_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _19614_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _19615_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _19616_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _19617_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _19618_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19619_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19620_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19621_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19622_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19623_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19624_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19625_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19626_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19627_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19628_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19629_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _19630_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _19631_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _19632_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _19633_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _19634_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _19635_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _19636_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _19637_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _19638_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _19639_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _19640_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19641_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00572_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19642_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00573_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19643_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00574_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19644_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00575_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19645_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00576_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19646_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00577_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19647_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00578_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19648_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00579_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19649_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00580_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19650_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00581_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19651_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00582_),
    .Q(\rbzero.spi_registers.new_mapd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19652_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00583_),
    .Q(\rbzero.spi_registers.new_mapd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19653_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00584_),
    .Q(\rbzero.spi_registers.new_mapd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19654_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00585_),
    .Q(\rbzero.spi_registers.new_mapd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19655_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00586_),
    .Q(\rbzero.spi_registers.new_mapd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19656_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00587_),
    .Q(\rbzero.spi_registers.new_mapd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19657_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00588_),
    .Q(\rbzero.spi_registers.new_mapd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19658_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00589_),
    .Q(\rbzero.spi_registers.new_mapd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19659_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00590_),
    .Q(\rbzero.spi_registers.new_mapd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19660_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00591_),
    .Q(\rbzero.spi_registers.new_mapd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19661_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00592_),
    .Q(\rbzero.spi_registers.new_mapd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19662_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00593_),
    .Q(\rbzero.spi_registers.new_mapd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19663_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00594_),
    .Q(\rbzero.spi_registers.new_mapd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19664_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00595_),
    .Q(\rbzero.spi_registers.new_mapd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19665_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00596_),
    .Q(\rbzero.spi_registers.new_mapd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19666_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00597_),
    .Q(\rbzero.spi_registers.new_mapd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19667_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00598_),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_1 _19668_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00599_),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_1 _19669_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00600_),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_1 _19670_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00601_),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_4 _19671_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00602_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19672_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00603_),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19673_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00604_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _19674_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00605_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _19675_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00606_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _19676_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00607_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _19677_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00608_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _19678_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00609_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19679_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00610_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19680_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00611_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _19681_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00612_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19682_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00613_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19683_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00614_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19684_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00615_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19685_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00616_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19686_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00617_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19687_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00618_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19688_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00619_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19689_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00620_),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_1 _19690_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00621_),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_1 _19691_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00622_),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_2 _19692_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00623_),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_4 _19693_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00624_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_2 _19694_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00625_),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19695_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00626_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _19696_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00627_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _19697_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00628_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _19698_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00629_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _19699_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00630_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _19700_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00631_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19701_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00632_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19702_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00633_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19703_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00634_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19704_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00635_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _19705_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00636_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19706_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00637_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19707_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00638_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19708_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00639_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19709_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00640_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19710_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00641_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19711_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00642_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19712_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00643_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19713_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00644_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19714_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00645_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19715_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00646_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19716_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00647_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19717_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00648_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19718_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00649_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19719_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00650_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19720_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00651_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19721_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00652_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19722_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00653_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19723_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00654_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19724_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00655_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19725_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00656_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19726_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00657_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19727_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00658_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19728_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00659_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19729_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00660_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19730_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00661_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19731_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00662_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19732_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00663_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19733_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00664_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19734_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00665_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19735_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00666_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19736_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00667_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19737_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00668_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19738_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00669_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19739_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00670_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19740_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00671_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19741_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00672_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19742_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00673_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19743_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00674_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19744_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00675_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19745_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00676_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19746_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00677_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19747_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00678_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19748_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00679_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19749_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00680_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19750_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00681_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _19751_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00682_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _19752_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00683_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _19753_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00684_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _19754_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00685_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _19755_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00686_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _19756_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00687_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _19757_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00688_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _19758_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00689_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _19759_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00690_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _19760_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00691_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _19761_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00692_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _19762_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00693_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _19763_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00694_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _19764_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00695_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _19765_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00696_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _19766_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00697_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _19767_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00698_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _19768_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00699_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _19769_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00700_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _19770_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00701_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _19771_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00702_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _19772_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00703_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _19773_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00704_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _19774_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00705_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _19775_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00706_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _19776_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00707_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _19777_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00708_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _19778_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00709_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _19779_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00710_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _19780_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00711_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _19781_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00712_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _19782_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00713_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _19783_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00714_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _19784_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00715_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _19785_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00716_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _19786_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00717_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _19787_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00718_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _19788_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00719_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _19789_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00720_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _19790_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00721_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _19791_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00722_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_2 _19792_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00723_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19793_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00724_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19794_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00725_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _19795_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00726_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19796_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00727_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_2 _19797_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00728_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19798_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00729_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19799_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00730_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19800_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00731_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19801_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00732_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19802_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00733_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19803_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00734_),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19804_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00735_),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19805_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00736_),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19806_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00737_),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19807_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00738_),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19808_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00739_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19809_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00740_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19810_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00741_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19811_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00742_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19812_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00743_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19813_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00744_),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _19814_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00745_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19815_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00746_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19816_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00747_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19817_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00748_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19818_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00749_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19819_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00750_),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19820_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00751_),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19821_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00752_),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19822_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00753_),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19823_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00754_),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19824_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00755_),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19825_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00756_),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19826_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00757_),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19827_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00758_),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19828_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00759_),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sky130_fd_sc_hd__dfxtp_2 _19829_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00760_),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _19830_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00761_),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19831_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00762_),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19832_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00763_),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19833_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00764_),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19834_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00765_),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19835_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00766_),
    .Q(\rbzero.map_overlay.i_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19836_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00767_),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19837_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00768_),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19838_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00769_),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19839_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00770_),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19840_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00771_),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19841_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00772_),
    .Q(\rbzero.map_overlay.i_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19842_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00773_),
    .Q(\rbzero.mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19843_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00774_),
    .Q(\rbzero.mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19844_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00775_),
    .Q(\rbzero.mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19845_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00776_),
    .Q(\rbzero.mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19846_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00777_),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19847_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00778_),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19848_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00779_),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19849_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00780_),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19850_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00781_),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19851_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00782_),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19852_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00783_),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19853_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00784_),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19854_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00785_),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19855_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00786_),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19856_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00787_),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19857_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00788_),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19858_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00789_),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19859_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00790_),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19860_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00791_),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19861_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00792_),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19862_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00793_),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19863_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00794_),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19864_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00795_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19865_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00796_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19866_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00797_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19867_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00798_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19868_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00799_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19869_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00800_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19870_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00801_),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _19871_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00802_),
    .Q(\rbzero.spi_registers.new_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19872_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00803_),
    .Q(\rbzero.spi_registers.new_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19873_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00804_),
    .Q(\rbzero.spi_registers.new_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19874_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00805_),
    .Q(\rbzero.spi_registers.new_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19875_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00806_),
    .Q(\rbzero.spi_registers.new_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19876_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00807_),
    .Q(\rbzero.spi_registers.new_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19877_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00808_),
    .Q(\rbzero.spi_registers.got_new_sky ));
 sky130_fd_sc_hd__dfxtp_1 _19878_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00809_),
    .Q(\rbzero.spi_registers.new_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19879_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00810_),
    .Q(\rbzero.spi_registers.new_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19880_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00811_),
    .Q(\rbzero.spi_registers.new_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19881_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00812_),
    .Q(\rbzero.spi_registers.new_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19882_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00813_),
    .Q(\rbzero.spi_registers.new_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19883_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00814_),
    .Q(\rbzero.spi_registers.new_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19884_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00815_),
    .Q(\rbzero.spi_registers.got_new_floor ));
 sky130_fd_sc_hd__dfxtp_1 _19885_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00816_),
    .Q(\rbzero.spi_registers.new_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19886_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00817_),
    .Q(\rbzero.spi_registers.new_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19887_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00818_),
    .Q(\rbzero.spi_registers.new_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19888_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00819_),
    .Q(\rbzero.spi_registers.new_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19889_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00820_),
    .Q(\rbzero.spi_registers.new_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19890_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00821_),
    .Q(\rbzero.spi_registers.new_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19891_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00822_),
    .Q(\rbzero.spi_registers.got_new_leak ));
 sky130_fd_sc_hd__dfxtp_1 _19892_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00823_),
    .Q(\rbzero.spi_registers.new_other[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19893_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00824_),
    .Q(\rbzero.spi_registers.new_other[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19894_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00825_),
    .Q(\rbzero.spi_registers.new_other[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19895_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00826_),
    .Q(\rbzero.spi_registers.new_other[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19896_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00827_),
    .Q(\rbzero.spi_registers.new_other[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19897_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00828_),
    .Q(\rbzero.spi_registers.new_other[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19898_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00829_),
    .Q(\rbzero.spi_registers.new_other[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19899_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00830_),
    .Q(\rbzero.spi_registers.new_other[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19900_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00831_),
    .Q(\rbzero.spi_registers.new_other[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19901_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00832_),
    .Q(\rbzero.spi_registers.new_other[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19902_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00833_),
    .Q(\rbzero.spi_registers.got_new_other ));
 sky130_fd_sc_hd__dfxtp_1 _19903_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00834_),
    .Q(\rbzero.spi_registers.new_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19904_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00835_),
    .Q(\rbzero.spi_registers.new_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19905_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00836_),
    .Q(\rbzero.spi_registers.new_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19906_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00837_),
    .Q(\rbzero.spi_registers.new_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19907_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00838_),
    .Q(\rbzero.spi_registers.new_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19908_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00839_),
    .Q(\rbzero.spi_registers.new_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19909_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00840_),
    .Q(\rbzero.spi_registers.got_new_vshift ));
 sky130_fd_sc_hd__dfxtp_1 _19910_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00841_),
    .Q(\rbzero.spi_registers.new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _19911_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00842_),
    .Q(\rbzero.spi_registers.got_new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _19912_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00843_),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _19913_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00844_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19914_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00845_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19915_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00846_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19916_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00847_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19917_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00848_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19918_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00849_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19919_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00850_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19920_ (.CLK(net149),
    .D(_00851_),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19921_ (.CLK(net150),
    .D(_00852_),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19922_ (.CLK(net151),
    .D(_00853_),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19923_ (.CLK(net152),
    .D(_00854_),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19924_ (.CLK(net153),
    .D(_00855_),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19925_ (.CLK(net154),
    .D(_00856_),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19926_ (.CLK(net155),
    .D(_00857_),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19927_ (.CLK(net156),
    .D(_00858_),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19928_ (.CLK(net157),
    .D(_00859_),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19929_ (.CLK(net158),
    .D(_00860_),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19930_ (.CLK(net159),
    .D(_00861_),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19931_ (.CLK(net160),
    .D(_00862_),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19932_ (.CLK(net161),
    .D(_00863_),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19933_ (.CLK(net162),
    .D(_00864_),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19934_ (.CLK(net163),
    .D(_00865_),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19935_ (.CLK(net164),
    .D(_00866_),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19936_ (.CLK(net165),
    .D(_00867_),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19937_ (.CLK(net166),
    .D(_00868_),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19938_ (.CLK(net167),
    .D(_00869_),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19939_ (.CLK(net168),
    .D(_00870_),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19940_ (.CLK(net169),
    .D(_00871_),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19941_ (.CLK(net170),
    .D(_00872_),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19942_ (.CLK(net171),
    .D(_00873_),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19943_ (.CLK(net172),
    .D(_00874_),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19944_ (.CLK(net173),
    .D(_00875_),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19945_ (.CLK(net174),
    .D(_00876_),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19946_ (.CLK(net175),
    .D(_00877_),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19947_ (.CLK(net176),
    .D(_00878_),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19948_ (.CLK(net177),
    .D(_00879_),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19949_ (.CLK(net178),
    .D(_00880_),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19950_ (.CLK(net179),
    .D(_00881_),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19951_ (.CLK(net180),
    .D(_00882_),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19952_ (.CLK(net181),
    .D(_00883_),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _19953_ (.CLK(net182),
    .D(_00884_),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _19954_ (.CLK(net183),
    .D(_00885_),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _19955_ (.CLK(net184),
    .D(_00886_),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _19956_ (.CLK(net185),
    .D(_00887_),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _19957_ (.CLK(net186),
    .D(_00888_),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _19958_ (.CLK(net187),
    .D(_00889_),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _19959_ (.CLK(net188),
    .D(_00890_),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _19960_ (.CLK(net189),
    .D(_00891_),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _19961_ (.CLK(net190),
    .D(_00892_),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _19962_ (.CLK(net191),
    .D(_00893_),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _19963_ (.CLK(net192),
    .D(_00894_),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _19964_ (.CLK(net193),
    .D(_00895_),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _19965_ (.CLK(net194),
    .D(_00896_),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _19966_ (.CLK(net195),
    .D(_00897_),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _19967_ (.CLK(net196),
    .D(_00898_),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _19968_ (.CLK(net197),
    .D(_00899_),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _19969_ (.CLK(net198),
    .D(_00900_),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _19970_ (.CLK(net199),
    .D(_00901_),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _19971_ (.CLK(net200),
    .D(_00902_),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _19972_ (.CLK(net201),
    .D(_00903_),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _19973_ (.CLK(net202),
    .D(_00904_),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _19974_ (.CLK(net203),
    .D(_00905_),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _19975_ (.CLK(net204),
    .D(_00906_),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _19976_ (.CLK(net205),
    .D(_00907_),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _19977_ (.CLK(net206),
    .D(_00908_),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _19978_ (.CLK(net207),
    .D(_00909_),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _19979_ (.CLK(net208),
    .D(_00910_),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _19980_ (.CLK(net209),
    .D(_00911_),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _19981_ (.CLK(net210),
    .D(_00912_),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _19982_ (.CLK(net211),
    .D(_00913_),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _19983_ (.CLK(net212),
    .D(_00914_),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _19984_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00915_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19985_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00916_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19986_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00917_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19987_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00918_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19988_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00919_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19989_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00920_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19990_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00921_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19991_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00922_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19992_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00923_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19993_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00924_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19994_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00925_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19995_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00926_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19996_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00927_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19997_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00928_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19998_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00929_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19999_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00930_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20000_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00931_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20001_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00932_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20002_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00933_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20003_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00934_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20004_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00935_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20005_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00936_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20006_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00937_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20007_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00938_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20008_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00939_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20009_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00940_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20010_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00941_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20011_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00942_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20012_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00943_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20013_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00944_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20014_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00945_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20015_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00946_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20016_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00947_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20017_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00948_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20018_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00949_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20019_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00950_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20020_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00951_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20021_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00952_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20022_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00953_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20023_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00954_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20024_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00955_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20025_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00956_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20026_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00957_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20027_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00958_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20028_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00959_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20029_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00960_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20030_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00961_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20031_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00962_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20032_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00963_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20033_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00964_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20034_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00965_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20035_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00966_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20036_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00967_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20037_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00968_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20038_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00969_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20039_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00970_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20040_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00971_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20041_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00972_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20042_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00973_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20043_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00974_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20044_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00975_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20045_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00976_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20046_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00977_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20047_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00978_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20048_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00979_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _20049_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00980_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _20050_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00981_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _20051_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00982_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _20052_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00983_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _20053_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00984_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _20054_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00985_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _20055_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00986_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _20056_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00987_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _20057_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00988_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _20058_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00989_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20059_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00990_),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _20060_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00991_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20061_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00992_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20062_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00993_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20063_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00994_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20064_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00995_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20065_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00996_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20066_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00997_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20067_ (.CLK(clknet_3_4_0_i_clk),
    .D(_00998_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20068_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00999_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _20069_ (.CLK(clknet_leaf_67_i_clk),
    .D(_01000_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20070_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01001_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_4 _20071_ (.CLK(clknet_leaf_64_i_clk),
    .D(_01002_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _20072_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01003_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _20073_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01004_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20074_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01005_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20075_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01006_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20076_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01007_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20077_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01008_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20078_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01009_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20079_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01010_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20080_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01011_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20081_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01012_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20082_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01013_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20083_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01014_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20084_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01015_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20085_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01016_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20086_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01017_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20087_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01018_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20088_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01019_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20089_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01020_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20090_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01021_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20091_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01022_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20092_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01023_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20093_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01024_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20094_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01025_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20095_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01026_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20096_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01027_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20097_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01028_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20098_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01029_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20099_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01030_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20100_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01031_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20101_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01032_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20102_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01033_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20103_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01034_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20104_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01035_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20105_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01036_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20106_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01037_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20107_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01038_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20108_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01039_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20109_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01040_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _20110_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01041_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20111_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01042_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20112_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01043_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20113_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01044_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20114_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01045_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20115_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01046_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20116_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01047_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20117_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01048_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20118_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01049_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20119_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01050_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20120_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01051_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20121_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01052_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20122_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01053_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20123_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01054_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _20124_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01055_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _20125_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01056_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20126_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01057_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20127_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01058_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20128_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01059_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20129_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01060_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20130_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01061_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20131_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01062_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _20132_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01063_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20133_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01064_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20134_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01065_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20135_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01066_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20136_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01067_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20137_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01068_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20138_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01069_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20139_ (.CLK(clknet_leaf_0_i_clk),
    .D(_01070_),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_2 _20140_ (.CLK(clknet_leaf_26_i_clk),
    .D(_01071_),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_2 _20141_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01072_),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_2 _20142_ (.CLK(clknet_leaf_12_i_clk),
    .D(_01073_),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20143_ (.CLK(clknet_leaf_12_i_clk),
    .D(_01074_),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20144_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01075_),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20145_ (.CLK(clknet_leaf_12_i_clk),
    .D(_01076_),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20146_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01077_),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20147_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01078_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20148_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01079_),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20149_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01080_),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20150_ (.CLK(clknet_leaf_20_i_clk),
    .D(_01081_),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20151_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01082_),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20152_ (.CLK(clknet_leaf_18_i_clk),
    .D(_01083_),
    .Q(\rbzero.spi_registers.got_new_mapd ));
 sky130_fd_sc_hd__dfxtp_1 _20153_ (.CLK(net213),
    .D(_01084_),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20154_ (.CLK(net214),
    .D(_01085_),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20155_ (.CLK(net215),
    .D(_01086_),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20156_ (.CLK(net216),
    .D(_01087_),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20157_ (.CLK(net217),
    .D(_01088_),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20158_ (.CLK(net218),
    .D(_01089_),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20159_ (.CLK(net219),
    .D(_01090_),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20160_ (.CLK(net220),
    .D(_01091_),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20161_ (.CLK(net221),
    .D(_01092_),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20162_ (.CLK(net222),
    .D(_01093_),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20163_ (.CLK(net223),
    .D(_01094_),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20164_ (.CLK(net224),
    .D(_01095_),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20165_ (.CLK(net225),
    .D(_01096_),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20166_ (.CLK(net226),
    .D(_01097_),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20167_ (.CLK(net227),
    .D(_01098_),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20168_ (.CLK(net228),
    .D(_01099_),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20169_ (.CLK(net229),
    .D(_01100_),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20170_ (.CLK(net230),
    .D(_01101_),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20171_ (.CLK(net231),
    .D(_01102_),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20172_ (.CLK(net232),
    .D(_01103_),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20173_ (.CLK(net233),
    .D(_01104_),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20174_ (.CLK(net234),
    .D(_01105_),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20175_ (.CLK(net235),
    .D(_01106_),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20176_ (.CLK(net236),
    .D(_01107_),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20177_ (.CLK(net237),
    .D(_01108_),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20178_ (.CLK(net238),
    .D(_01109_),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20179_ (.CLK(net239),
    .D(_01110_),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20180_ (.CLK(net240),
    .D(_01111_),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20181_ (.CLK(net241),
    .D(_01112_),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20182_ (.CLK(net242),
    .D(_01113_),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20183_ (.CLK(net243),
    .D(_01114_),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20184_ (.CLK(net244),
    .D(_01115_),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20185_ (.CLK(net245),
    .D(_01116_),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20186_ (.CLK(net246),
    .D(_01117_),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20187_ (.CLK(net247),
    .D(_01118_),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20188_ (.CLK(net248),
    .D(_01119_),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20189_ (.CLK(net249),
    .D(_01120_),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20190_ (.CLK(net250),
    .D(_01121_),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20191_ (.CLK(net251),
    .D(_01122_),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20192_ (.CLK(net252),
    .D(_01123_),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20193_ (.CLK(net253),
    .D(_01124_),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20194_ (.CLK(net254),
    .D(_01125_),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20195_ (.CLK(net255),
    .D(_01126_),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20196_ (.CLK(net256),
    .D(_01127_),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20197_ (.CLK(net257),
    .D(_01128_),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20198_ (.CLK(net258),
    .D(_01129_),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20199_ (.CLK(net259),
    .D(_01130_),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20200_ (.CLK(net260),
    .D(_01131_),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20201_ (.CLK(net261),
    .D(_01132_),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20202_ (.CLK(net262),
    .D(_01133_),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20203_ (.CLK(net263),
    .D(_01134_),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20204_ (.CLK(net264),
    .D(_01135_),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20205_ (.CLK(net265),
    .D(_01136_),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20206_ (.CLK(net266),
    .D(_01137_),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20207_ (.CLK(net267),
    .D(_01138_),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20208_ (.CLK(net268),
    .D(_01139_),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20209_ (.CLK(net269),
    .D(_01140_),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20210_ (.CLK(net270),
    .D(_01141_),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20211_ (.CLK(net271),
    .D(_01142_),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20212_ (.CLK(net272),
    .D(_01143_),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20213_ (.CLK(net273),
    .D(_01144_),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20214_ (.CLK(net274),
    .D(_01145_),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20215_ (.CLK(net275),
    .D(_01146_),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20216_ (.CLK(net276),
    .D(_01147_),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20217_ (.CLK(net277),
    .D(_01148_),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20218_ (.CLK(net278),
    .D(_01149_),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20219_ (.CLK(net279),
    .D(_01150_),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20220_ (.CLK(net280),
    .D(_01151_),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20221_ (.CLK(net281),
    .D(_01152_),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20222_ (.CLK(net282),
    .D(_01153_),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20223_ (.CLK(net283),
    .D(_01154_),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20224_ (.CLK(net284),
    .D(_01155_),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20225_ (.CLK(net285),
    .D(_01156_),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20226_ (.CLK(net286),
    .D(_01157_),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20227_ (.CLK(net287),
    .D(_01158_),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20228_ (.CLK(net288),
    .D(_01159_),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20229_ (.CLK(net289),
    .D(_01160_),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20230_ (.CLK(net290),
    .D(_01161_),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20231_ (.CLK(net291),
    .D(_01162_),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20232_ (.CLK(net292),
    .D(_01163_),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20233_ (.CLK(net293),
    .D(_01164_),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20234_ (.CLK(net294),
    .D(_01165_),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20235_ (.CLK(net295),
    .D(_01166_),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20236_ (.CLK(net296),
    .D(_01167_),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20237_ (.CLK(net297),
    .D(_01168_),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20238_ (.CLK(net298),
    .D(_01169_),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20239_ (.CLK(net299),
    .D(_01170_),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20240_ (.CLK(net300),
    .D(_01171_),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20241_ (.CLK(net301),
    .D(_01172_),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20242_ (.CLK(net302),
    .D(_01173_),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20243_ (.CLK(net303),
    .D(_01174_),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20244_ (.CLK(net304),
    .D(_01175_),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20245_ (.CLK(net305),
    .D(_01176_),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20246_ (.CLK(net306),
    .D(_01177_),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20247_ (.CLK(net307),
    .D(_01178_),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20248_ (.CLK(net308),
    .D(_01179_),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20249_ (.CLK(net309),
    .D(_01180_),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20250_ (.CLK(net310),
    .D(_01181_),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20251_ (.CLK(net311),
    .D(_01182_),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20252_ (.CLK(net312),
    .D(_01183_),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20253_ (.CLK(net313),
    .D(_01184_),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20254_ (.CLK(net314),
    .D(_01185_),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20255_ (.CLK(net315),
    .D(_01186_),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20256_ (.CLK(net316),
    .D(_01187_),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20257_ (.CLK(net317),
    .D(_01188_),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20258_ (.CLK(net318),
    .D(_01189_),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20259_ (.CLK(net319),
    .D(_01190_),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20260_ (.CLK(net320),
    .D(_01191_),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20261_ (.CLK(net321),
    .D(_01192_),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20262_ (.CLK(net322),
    .D(_01193_),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20263_ (.CLK(net323),
    .D(_01194_),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20264_ (.CLK(net324),
    .D(_01195_),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20265_ (.CLK(net325),
    .D(_01196_),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20266_ (.CLK(net326),
    .D(_01197_),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20267_ (.CLK(net327),
    .D(_01198_),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20268_ (.CLK(net328),
    .D(_01199_),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20269_ (.CLK(net329),
    .D(_01200_),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20270_ (.CLK(net330),
    .D(_01201_),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20271_ (.CLK(net331),
    .D(_01202_),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20272_ (.CLK(net332),
    .D(_01203_),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20273_ (.CLK(net333),
    .D(_01204_),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20274_ (.CLK(net334),
    .D(_01205_),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20275_ (.CLK(net335),
    .D(_01206_),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20276_ (.CLK(net336),
    .D(_01207_),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20277_ (.CLK(net337),
    .D(_01208_),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20278_ (.CLK(net338),
    .D(_01209_),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20279_ (.CLK(net339),
    .D(_01210_),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20280_ (.CLK(net340),
    .D(_01211_),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20281_ (.CLK(net341),
    .D(_01212_),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20282_ (.CLK(net342),
    .D(_01213_),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20283_ (.CLK(net343),
    .D(_01214_),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20284_ (.CLK(net344),
    .D(_01215_),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20285_ (.CLK(net345),
    .D(_01216_),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20286_ (.CLK(net346),
    .D(_01217_),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20287_ (.CLK(net347),
    .D(_01218_),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20288_ (.CLK(net348),
    .D(_01219_),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20289_ (.CLK(net349),
    .D(_01220_),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20290_ (.CLK(net350),
    .D(_01221_),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20291_ (.CLK(net351),
    .D(_01222_),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20292_ (.CLK(net352),
    .D(_01223_),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20293_ (.CLK(net353),
    .D(_01224_),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20294_ (.CLK(net354),
    .D(_01225_),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20295_ (.CLK(net355),
    .D(_01226_),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20296_ (.CLK(net356),
    .D(_01227_),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20297_ (.CLK(net357),
    .D(_01228_),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20298_ (.CLK(net358),
    .D(_01229_),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20299_ (.CLK(net359),
    .D(_01230_),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20300_ (.CLK(net360),
    .D(_01231_),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20301_ (.CLK(net361),
    .D(_01232_),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20302_ (.CLK(net362),
    .D(_01233_),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20303_ (.CLK(net363),
    .D(_01234_),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20304_ (.CLK(net364),
    .D(_01235_),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20305_ (.CLK(net365),
    .D(_01236_),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20306_ (.CLK(net366),
    .D(_01237_),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20307_ (.CLK(net367),
    .D(_01238_),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20308_ (.CLK(net368),
    .D(_01239_),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20309_ (.CLK(net369),
    .D(_01240_),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20310_ (.CLK(net370),
    .D(_01241_),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20311_ (.CLK(net371),
    .D(_01242_),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20312_ (.CLK(net372),
    .D(_01243_),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20313_ (.CLK(net373),
    .D(_01244_),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20314_ (.CLK(net374),
    .D(_01245_),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20315_ (.CLK(net375),
    .D(_01246_),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20316_ (.CLK(net376),
    .D(_01247_),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20317_ (.CLK(net377),
    .D(_01248_),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20318_ (.CLK(net378),
    .D(_01249_),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20319_ (.CLK(net379),
    .D(_01250_),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20320_ (.CLK(net380),
    .D(_01251_),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20321_ (.CLK(net381),
    .D(_01252_),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20322_ (.CLK(net382),
    .D(_01253_),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20323_ (.CLK(net383),
    .D(_01254_),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20324_ (.CLK(net384),
    .D(_01255_),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20325_ (.CLK(net385),
    .D(_01256_),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20326_ (.CLK(net386),
    .D(_01257_),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20327_ (.CLK(net387),
    .D(_01258_),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20328_ (.CLK(net388),
    .D(_01259_),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20329_ (.CLK(net389),
    .D(_01260_),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20330_ (.CLK(net390),
    .D(_01261_),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20331_ (.CLK(net391),
    .D(_01262_),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20332_ (.CLK(net392),
    .D(_01263_),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20333_ (.CLK(net393),
    .D(_01264_),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20334_ (.CLK(net394),
    .D(_01265_),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20335_ (.CLK(net395),
    .D(_01266_),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20336_ (.CLK(net396),
    .D(_01267_),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20337_ (.CLK(net397),
    .D(_01268_),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20338_ (.CLK(net398),
    .D(_01269_),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20339_ (.CLK(net399),
    .D(_01270_),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20340_ (.CLK(net400),
    .D(_01271_),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20341_ (.CLK(net401),
    .D(_01272_),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20342_ (.CLK(net402),
    .D(_01273_),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20343_ (.CLK(net403),
    .D(_01274_),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20344_ (.CLK(net404),
    .D(_01275_),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20345_ (.CLK(net405),
    .D(_01276_),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20346_ (.CLK(net406),
    .D(_01277_),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20347_ (.CLK(net407),
    .D(_01278_),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20348_ (.CLK(net408),
    .D(_01279_),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20349_ (.CLK(net409),
    .D(_01280_),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20350_ (.CLK(net410),
    .D(_01281_),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20351_ (.CLK(net411),
    .D(_01282_),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20352_ (.CLK(net412),
    .D(_01283_),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20353_ (.CLK(net413),
    .D(_01284_),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20354_ (.CLK(net414),
    .D(_01285_),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20355_ (.CLK(net415),
    .D(_01286_),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20356_ (.CLK(net416),
    .D(_01287_),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20357_ (.CLK(net417),
    .D(_01288_),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20358_ (.CLK(net418),
    .D(_01289_),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20359_ (.CLK(net419),
    .D(_01290_),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20360_ (.CLK(net420),
    .D(_01291_),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20361_ (.CLK(net421),
    .D(_01292_),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20362_ (.CLK(net422),
    .D(_01293_),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20363_ (.CLK(net423),
    .D(_01294_),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20364_ (.CLK(net424),
    .D(_01295_),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20365_ (.CLK(net425),
    .D(_01296_),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20366_ (.CLK(net426),
    .D(_01297_),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20367_ (.CLK(net427),
    .D(_01298_),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20368_ (.CLK(net428),
    .D(_01299_),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20369_ (.CLK(net429),
    .D(_01300_),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20370_ (.CLK(net430),
    .D(_01301_),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20371_ (.CLK(net431),
    .D(_01302_),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20372_ (.CLK(net432),
    .D(_01303_),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20373_ (.CLK(net433),
    .D(_01304_),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20374_ (.CLK(net434),
    .D(_01305_),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20375_ (.CLK(net435),
    .D(_01306_),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20376_ (.CLK(net436),
    .D(_01307_),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20377_ (.CLK(net437),
    .D(_01308_),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20378_ (.CLK(net438),
    .D(_01309_),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20379_ (.CLK(net439),
    .D(_01310_),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20380_ (.CLK(net440),
    .D(_01311_),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20381_ (.CLK(net441),
    .D(_01312_),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20382_ (.CLK(net442),
    .D(_01313_),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20383_ (.CLK(net443),
    .D(_01314_),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20384_ (.CLK(net444),
    .D(_01315_),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20385_ (.CLK(net445),
    .D(_01316_),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20386_ (.CLK(net446),
    .D(_01317_),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20387_ (.CLK(net447),
    .D(_01318_),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20388_ (.CLK(net448),
    .D(_01319_),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20389_ (.CLK(net449),
    .D(_01320_),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20390_ (.CLK(net450),
    .D(_01321_),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20391_ (.CLK(net451),
    .D(_01322_),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20392_ (.CLK(net452),
    .D(_01323_),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20393_ (.CLK(net453),
    .D(_01324_),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20394_ (.CLK(net454),
    .D(_01325_),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20395_ (.CLK(net455),
    .D(_01326_),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20396_ (.CLK(net456),
    .D(_01327_),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20397_ (.CLK(net457),
    .D(_01328_),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20398_ (.CLK(net458),
    .D(_01329_),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20399_ (.CLK(net459),
    .D(_01330_),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20400_ (.CLK(net460),
    .D(_01331_),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20401_ (.CLK(net461),
    .D(_01332_),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20402_ (.CLK(net462),
    .D(_01333_),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20403_ (.CLK(net463),
    .D(_01334_),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20404_ (.CLK(net464),
    .D(_01335_),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20405_ (.CLK(net465),
    .D(_01336_),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20406_ (.CLK(net466),
    .D(_01337_),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20407_ (.CLK(net467),
    .D(_01338_),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20408_ (.CLK(net468),
    .D(_01339_),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20409_ (.CLK(net469),
    .D(_01340_),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20410_ (.CLK(net470),
    .D(_01341_),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20411_ (.CLK(net471),
    .D(_01342_),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20412_ (.CLK(net472),
    .D(_01343_),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20413_ (.CLK(net473),
    .D(_01344_),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20414_ (.CLK(net474),
    .D(_01345_),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20415_ (.CLK(net475),
    .D(_01346_),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20416_ (.CLK(net476),
    .D(_01347_),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20417_ (.CLK(net477),
    .D(_01348_),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20418_ (.CLK(net478),
    .D(_01349_),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20419_ (.CLK(net479),
    .D(_01350_),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20420_ (.CLK(net480),
    .D(_01351_),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20421_ (.CLK(net481),
    .D(_01352_),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20422_ (.CLK(net482),
    .D(_01353_),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20423_ (.CLK(net483),
    .D(_01354_),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20424_ (.CLK(net484),
    .D(_01355_),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20425_ (.CLK(net485),
    .D(_01356_),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20426_ (.CLK(net486),
    .D(_01357_),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20427_ (.CLK(net487),
    .D(_01358_),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20428_ (.CLK(net488),
    .D(_01359_),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20429_ (.CLK(net489),
    .D(_01360_),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20430_ (.CLK(net490),
    .D(_01361_),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20431_ (.CLK(net491),
    .D(_01362_),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20432_ (.CLK(net492),
    .D(_01363_),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20433_ (.CLK(net493),
    .D(_01364_),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20434_ (.CLK(net494),
    .D(_01365_),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20435_ (.CLK(net495),
    .D(_01366_),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20436_ (.CLK(net496),
    .D(_01367_),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20437_ (.CLK(net497),
    .D(_01368_),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20438_ (.CLK(net498),
    .D(_01369_),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20439_ (.CLK(net499),
    .D(_01370_),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20440_ (.CLK(net500),
    .D(_01371_),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20441_ (.CLK(net501),
    .D(_01372_),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20442_ (.CLK(net502),
    .D(_01373_),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20443_ (.CLK(net503),
    .D(_01374_),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20444_ (.CLK(net504),
    .D(_01375_),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20445_ (.CLK(net505),
    .D(_01376_),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20446_ (.CLK(net506),
    .D(_01377_),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20447_ (.CLK(net507),
    .D(_01378_),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20448_ (.CLK(net508),
    .D(_01379_),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20449_ (.CLK(net129),
    .D(_01380_),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20450_ (.CLK(net130),
    .D(_01381_),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20451_ (.CLK(net131),
    .D(_01382_),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20452_ (.CLK(net132),
    .D(_01383_),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20453_ (.CLK(net133),
    .D(_01384_),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20454_ (.CLK(net134),
    .D(_01385_),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20455_ (.CLK(net135),
    .D(_01386_),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20456_ (.CLK(net136),
    .D(_01387_),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20457_ (.CLK(net137),
    .D(_01388_),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20458_ (.CLK(net138),
    .D(_01389_),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20459_ (.CLK(net139),
    .D(_01390_),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20460_ (.CLK(net140),
    .D(_01391_),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20461_ (.CLK(net141),
    .D(_01392_),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20462_ (.CLK(net142),
    .D(_01393_),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20463_ (.CLK(net143),
    .D(_01394_),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20464_ (.CLK(net144),
    .D(_01395_),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20465_ (.CLK(net145),
    .D(_01396_),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20466_ (.CLK(net146),
    .D(_01397_),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20467_ (.CLK(net147),
    .D(_01398_),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20468_ (.CLK(net148),
    .D(_01399_),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20469_ (.CLK(net125),
    .D(_01400_),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20470_ (.CLK(net126),
    .D(_01401_),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20471_ (.CLK(net127),
    .D(_01402_),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20472_ (.CLK(net128),
    .D(_01403_),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20473_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01404_),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20474_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01405_),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20475_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01406_),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20476_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01407_),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20477_ (.CLK(clknet_leaf_63_i_clk),
    .D(_01408_),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20478_ (.CLK(clknet_leaf_66_i_clk),
    .D(_01409_),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20479_ (.CLK(clknet_leaf_63_i_clk),
    .D(_01410_),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20480_ (.CLK(clknet_leaf_62_i_clk),
    .D(_01411_),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20481_ (.CLK(clknet_leaf_63_i_clk),
    .D(_01412_),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20482_ (.CLK(clknet_leaf_61_i_clk),
    .D(_01413_),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20483_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01414_),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20484_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01415_),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20485_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01416_),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20486_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01417_),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20487_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01418_),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20488_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01419_),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20489_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01420_),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20490_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01421_),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20491_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01422_),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20492_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01423_),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20493_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01424_),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20494_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01425_),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20495_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01426_),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20496_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01427_),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20497_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01428_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20498_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01429_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20499_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01430_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20500_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01431_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20501_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01432_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20502_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01433_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20503_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01434_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20504_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01435_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20505_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01436_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20506_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01437_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20507_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01438_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20508_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01439_),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20509_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01440_),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20510_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01441_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20511_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01442_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20512_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01443_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20513_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01444_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20514_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01445_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20515_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01446_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20516_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01447_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20517_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01448_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20518_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01449_),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20519_ (.CLK(clknet_leaf_24_i_clk),
    .D(_01450_),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20520_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01451_),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20521_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01452_),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20522_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01453_),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20523_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01454_),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20524_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01455_),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20525_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01456_),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.HI(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.HI(net109));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.HI(net110));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.HI(net111));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_122 (.HI(net122));
 sky130_fd_sc_hd__inv_2 _11708__1 (.A(clknet_1_1__leaf__04486_),
    .Y(net123));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.HI(net107));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(i_debug_map_overlay),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(i_debug_vec_overlay),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(i_gpout0_sel[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(i_gpout0_sel[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(i_gpout0_sel[2]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(i_gpout0_sel[3]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(i_gpout0_sel[4]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(i_gpout0_sel[5]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(i_gpout1_sel[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(i_gpout1_sel[1]),
    .X(net10));
 sky130_fd_sc_hd__buf_6 input11 (.A(i_gpout1_sel[2]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(i_gpout1_sel[3]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(i_gpout1_sel[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 input14 (.A(i_gpout1_sel[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 input15 (.A(i_gpout2_sel[0]),
    .X(net15));
 sky130_fd_sc_hd__buf_6 input16 (.A(i_gpout2_sel[1]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(i_gpout2_sel[2]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(i_gpout2_sel[3]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_8 input19 (.A(i_gpout2_sel[4]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(i_gpout2_sel[5]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(i_gpout3_sel[0]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(i_gpout3_sel[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(i_gpout3_sel[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(i_gpout3_sel[3]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_8 input25 (.A(i_gpout3_sel[4]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(i_gpout3_sel[5]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(i_gpout4_sel[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(i_gpout4_sel[1]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(i_gpout4_sel[2]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(i_gpout4_sel[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(i_gpout4_sel[4]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(i_gpout4_sel[5]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(i_gpout5_sel[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_6 input34 (.A(i_gpout5_sel[1]),
    .X(net34));
 sky130_fd_sc_hd__buf_6 input35 (.A(i_gpout5_sel[2]),
    .X(net35));
 sky130_fd_sc_hd__buf_6 input36 (.A(i_gpout5_sel[3]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_8 input37 (.A(i_gpout5_sel[4]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(i_gpout5_sel[5]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_16 input39 (.A(i_mode[0]),
    .X(net39));
 sky130_fd_sc_hd__buf_8 input40 (.A(i_mode[1]),
    .X(net40));
 sky130_fd_sc_hd__buf_4 input41 (.A(i_mode[2]),
    .X(net41));
 sky130_fd_sc_hd__buf_8 input42 (.A(i_reg_csb),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(i_reg_mosi),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(i_reg_sclk),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(i_reset_lock_a),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input46 (.A(i_reset_lock_b),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(i_tex_in[0]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_tex_in[1]),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(i_tex_in[2]),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input50 (.A(i_tex_in[3]),
    .X(net50));
 sky130_fd_sc_hd__buf_8 input51 (.A(i_vec_csb),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(i_vec_mosi),
    .X(net52));
 sky130_fd_sc_hd__buf_8 input53 (.A(i_vec_sclk),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(o_hsync));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(o_reset));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(o_tex_csb));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(o_tex_out0));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net123),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(o_vsync));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_73 (.LO(net73));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_1_0__leaf__04486_),
    .Y(net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04486_ (.A(_04486_),
    .X(clknet_0__04486_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04486_ (.A(clknet_0__04486_),
    .X(clknet_1_0__leaf__04486_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04486_ (.A(clknet_0__04486_),
    .X(clknet_1_1__leaf__04486_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02755_ (.A(_02755_),
    .X(clknet_0__02755_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02755_ (.A(clknet_0__02755_),
    .X(clknet_1_0__leaf__02755_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02755_ (.A(clknet_0__02755_),
    .X(clknet_1_1__leaf__02755_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02754_ (.A(_02754_),
    .X(clknet_0__02754_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02754_ (.A(clknet_0__02754_),
    .X(clknet_1_0__leaf__02754_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02754_ (.A(clknet_0__02754_),
    .X(clknet_1_1__leaf__02754_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02743_ (.A(_02743_),
    .X(clknet_0__02743_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02743_ (.A(clknet_0__02743_),
    .X(clknet_1_0__leaf__02743_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02743_ (.A(clknet_0__02743_),
    .X(clknet_1_1__leaf__02743_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02753_ (.A(_02753_),
    .X(clknet_0__02753_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02753_ (.A(clknet_0__02753_),
    .X(clknet_1_0__leaf__02753_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02753_ (.A(clknet_0__02753_),
    .X(clknet_1_1__leaf__02753_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02752_ (.A(_02752_),
    .X(clknet_0__02752_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02752_ (.A(clknet_0__02752_),
    .X(clknet_1_0__leaf__02752_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02752_ (.A(clknet_0__02752_),
    .X(clknet_1_1__leaf__02752_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02751_ (.A(_02751_),
    .X(clknet_0__02751_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02751_ (.A(clknet_0__02751_),
    .X(clknet_1_0__leaf__02751_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02751_ (.A(clknet_0__02751_),
    .X(clknet_1_1__leaf__02751_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02750_ (.A(_02750_),
    .X(clknet_0__02750_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02750_ (.A(clknet_0__02750_),
    .X(clknet_1_0__leaf__02750_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02750_ (.A(clknet_0__02750_),
    .X(clknet_1_1__leaf__02750_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02749_ (.A(_02749_),
    .X(clknet_0__02749_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02749_ (.A(clknet_0__02749_),
    .X(clknet_1_0__leaf__02749_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02749_ (.A(clknet_0__02749_),
    .X(clknet_1_1__leaf__02749_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02748_ (.A(_02748_),
    .X(clknet_0__02748_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02748_ (.A(clknet_0__02748_),
    .X(clknet_1_0__leaf__02748_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02748_ (.A(clknet_0__02748_),
    .X(clknet_1_1__leaf__02748_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02747_ (.A(_02747_),
    .X(clknet_0__02747_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02747_ (.A(clknet_0__02747_),
    .X(clknet_1_0__leaf__02747_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02747_ (.A(clknet_0__02747_),
    .X(clknet_1_1__leaf__02747_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02746_ (.A(_02746_),
    .X(clknet_0__02746_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02746_ (.A(clknet_0__02746_),
    .X(clknet_1_0__leaf__02746_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02746_ (.A(clknet_0__02746_),
    .X(clknet_1_1__leaf__02746_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02745_ (.A(_02745_),
    .X(clknet_0__02745_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02745_ (.A(clknet_0__02745_),
    .X(clknet_1_0__leaf__02745_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02745_ (.A(clknet_0__02745_),
    .X(clknet_1_1__leaf__02745_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02744_ (.A(_02744_),
    .X(clknet_0__02744_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02744_ (.A(clknet_0__02744_),
    .X(clknet_1_0__leaf__02744_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02744_ (.A(clknet_0__02744_),
    .X(clknet_1_1__leaf__02744_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02732_ (.A(_02732_),
    .X(clknet_0__02732_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02732_ (.A(clknet_0__02732_),
    .X(clknet_1_0__leaf__02732_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02732_ (.A(clknet_0__02732_),
    .X(clknet_1_1__leaf__02732_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02742_ (.A(_02742_),
    .X(clknet_0__02742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02742_ (.A(clknet_0__02742_),
    .X(clknet_1_0__leaf__02742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02742_ (.A(clknet_0__02742_),
    .X(clknet_1_1__leaf__02742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02741_ (.A(_02741_),
    .X(clknet_0__02741_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02741_ (.A(clknet_0__02741_),
    .X(clknet_1_0__leaf__02741_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02741_ (.A(clknet_0__02741_),
    .X(clknet_1_1__leaf__02741_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02740_ (.A(_02740_),
    .X(clknet_0__02740_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02740_ (.A(clknet_0__02740_),
    .X(clknet_1_0__leaf__02740_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02740_ (.A(clknet_0__02740_),
    .X(clknet_1_1__leaf__02740_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02739_ (.A(_02739_),
    .X(clknet_0__02739_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02739_ (.A(clknet_0__02739_),
    .X(clknet_1_0__leaf__02739_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02739_ (.A(clknet_0__02739_),
    .X(clknet_1_1__leaf__02739_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02738_ (.A(_02738_),
    .X(clknet_0__02738_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02738_ (.A(clknet_0__02738_),
    .X(clknet_1_0__leaf__02738_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02738_ (.A(clknet_0__02738_),
    .X(clknet_1_1__leaf__02738_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02737_ (.A(_02737_),
    .X(clknet_0__02737_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02737_ (.A(clknet_0__02737_),
    .X(clknet_1_0__leaf__02737_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02737_ (.A(clknet_0__02737_),
    .X(clknet_1_1__leaf__02737_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02736_ (.A(_02736_),
    .X(clknet_0__02736_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02736_ (.A(clknet_0__02736_),
    .X(clknet_1_0__leaf__02736_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02736_ (.A(clknet_0__02736_),
    .X(clknet_1_1__leaf__02736_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02735_ (.A(_02735_),
    .X(clknet_0__02735_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02735_ (.A(clknet_0__02735_),
    .X(clknet_1_0__leaf__02735_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02735_ (.A(clknet_0__02735_),
    .X(clknet_1_1__leaf__02735_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02734_ (.A(_02734_),
    .X(clknet_0__02734_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02734_ (.A(clknet_0__02734_),
    .X(clknet_1_0__leaf__02734_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02734_ (.A(clknet_0__02734_),
    .X(clknet_1_1__leaf__02734_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02733_ (.A(_02733_),
    .X(clknet_0__02733_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02733_ (.A(clknet_0__02733_),
    .X(clknet_1_0__leaf__02733_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02733_ (.A(clknet_0__02733_),
    .X(clknet_1_1__leaf__02733_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02440_ (.A(_02440_),
    .X(clknet_0__02440_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02440_ (.A(clknet_0__02440_),
    .X(clknet_1_0__leaf__02440_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02440_ (.A(clknet_0__02440_),
    .X(clknet_1_1__leaf__02440_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02731_ (.A(_02731_),
    .X(clknet_0__02731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02731_ (.A(clknet_0__02731_),
    .X(clknet_1_0__leaf__02731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02731_ (.A(clknet_0__02731_),
    .X(clknet_1_1__leaf__02731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02730_ (.A(_02730_),
    .X(clknet_0__02730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02730_ (.A(clknet_0__02730_),
    .X(clknet_1_0__leaf__02730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02730_ (.A(clknet_0__02730_),
    .X(clknet_1_1__leaf__02730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02729_ (.A(_02729_),
    .X(clknet_0__02729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02729_ (.A(clknet_0__02729_),
    .X(clknet_1_0__leaf__02729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02729_ (.A(clknet_0__02729_),
    .X(clknet_1_1__leaf__02729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02728_ (.A(_02728_),
    .X(clknet_0__02728_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02728_ (.A(clknet_0__02728_),
    .X(clknet_1_0__leaf__02728_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02728_ (.A(clknet_0__02728_),
    .X(clknet_1_1__leaf__02728_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02727_ (.A(_02727_),
    .X(clknet_0__02727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02727_ (.A(clknet_0__02727_),
    .X(clknet_1_0__leaf__02727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02727_ (.A(clknet_0__02727_),
    .X(clknet_1_1__leaf__02727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02726_ (.A(_02726_),
    .X(clknet_0__02726_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02726_ (.A(clknet_0__02726_),
    .X(clknet_1_0__leaf__02726_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02726_ (.A(clknet_0__02726_),
    .X(clknet_1_1__leaf__02726_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02725_ (.A(_02725_),
    .X(clknet_0__02725_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02725_ (.A(clknet_0__02725_),
    .X(clknet_1_0__leaf__02725_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02725_ (.A(clknet_0__02725_),
    .X(clknet_1_1__leaf__02725_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02724_ (.A(_02724_),
    .X(clknet_0__02724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02724_ (.A(clknet_0__02724_),
    .X(clknet_1_0__leaf__02724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02724_ (.A(clknet_0__02724_),
    .X(clknet_1_1__leaf__02724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02723_ (.A(_02723_),
    .X(clknet_0__02723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02723_ (.A(clknet_0__02723_),
    .X(clknet_1_0__leaf__02723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02723_ (.A(clknet_0__02723_),
    .X(clknet_1_1__leaf__02723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02441_ (.A(_02441_),
    .X(clknet_0__02441_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02441_ (.A(clknet_0__02441_),
    .X(clknet_1_0__leaf__02441_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02441_ (.A(clknet_0__02441_),
    .X(clknet_1_1__leaf__02441_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02433_ (.A(_02433_),
    .X(clknet_0__02433_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02433_ (.A(clknet_0__02433_),
    .X(clknet_1_0__leaf__02433_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02433_ (.A(clknet_0__02433_),
    .X(clknet_1_1__leaf__02433_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02439_ (.A(_02439_),
    .X(clknet_0__02439_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02439_ (.A(clknet_0__02439_),
    .X(clknet_1_0__leaf__02439_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02439_ (.A(clknet_0__02439_),
    .X(clknet_1_1__leaf__02439_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02438_ (.A(_02438_),
    .X(clknet_0__02438_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02438_ (.A(clknet_0__02438_),
    .X(clknet_1_0__leaf__02438_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02438_ (.A(clknet_0__02438_),
    .X(clknet_1_1__leaf__02438_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02437_ (.A(_02437_),
    .X(clknet_0__02437_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02437_ (.A(clknet_0__02437_),
    .X(clknet_1_0__leaf__02437_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02437_ (.A(clknet_0__02437_),
    .X(clknet_1_1__leaf__02437_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02436_ (.A(_02436_),
    .X(clknet_0__02436_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02436_ (.A(clknet_0__02436_),
    .X(clknet_1_0__leaf__02436_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02436_ (.A(clknet_0__02436_),
    .X(clknet_1_1__leaf__02436_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02435_ (.A(_02435_),
    .X(clknet_0__02435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02435_ (.A(clknet_0__02435_),
    .X(clknet_1_0__leaf__02435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02435_ (.A(clknet_0__02435_),
    .X(clknet_1_1__leaf__02435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02434_ (.A(_02434_),
    .X(clknet_0__02434_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02434_ (.A(clknet_0__02434_),
    .X(clknet_1_0__leaf__02434_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02434_ (.A(clknet_0__02434_),
    .X(clknet_1_1__leaf__02434_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rbzero.tex_r1[40] ),
    .X(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_04834_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_06855_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_06938_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_07052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_07147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_07817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_03688_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_06916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_06916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_07151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_08958_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net49));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1192 ();
 assign o_rgb[0] = net73;
 assign o_rgb[10] = net81;
 assign o_rgb[11] = net82;
 assign o_rgb[12] = net83;
 assign o_rgb[13] = net84;
 assign o_rgb[16] = net85;
 assign o_rgb[17] = net86;
 assign o_rgb[18] = net87;
 assign o_rgb[19] = net88;
 assign o_rgb[1] = net74;
 assign o_rgb[20] = net89;
 assign o_rgb[21] = net90;
 assign o_rgb[2] = net75;
 assign o_rgb[3] = net76;
 assign o_rgb[4] = net77;
 assign o_rgb[5] = net78;
 assign o_rgb[8] = net79;
 assign o_rgb[9] = net80;
 assign ones[0] = net107;
 assign ones[10] = net117;
 assign ones[11] = net118;
 assign ones[12] = net119;
 assign ones[13] = net120;
 assign ones[14] = net121;
 assign ones[15] = net122;
 assign ones[1] = net108;
 assign ones[2] = net109;
 assign ones[3] = net110;
 assign ones[4] = net111;
 assign ones[5] = net112;
 assign ones[6] = net113;
 assign ones[7] = net114;
 assign ones[8] = net115;
 assign ones[9] = net116;
 assign zeros[0] = net91;
 assign zeros[10] = net101;
 assign zeros[11] = net102;
 assign zeros[12] = net103;
 assign zeros[13] = net104;
 assign zeros[14] = net105;
 assign zeros[15] = net106;
 assign zeros[1] = net92;
 assign zeros[2] = net93;
 assign zeros[3] = net94;
 assign zeros[4] = net95;
 assign zeros[5] = net96;
 assign zeros[6] = net97;
 assign zeros[7] = net98;
 assign zeros[8] = net99;
 assign zeros[9] = net100;
endmodule

