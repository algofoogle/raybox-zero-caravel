magic
tech sky130A
magscale 1 2
timestamp 1699096299
<< nwell >>
rect 1066 116677 116786 117243
rect 1066 115589 116786 116155
rect 1066 114501 116786 115067
rect 1066 113413 116786 113979
rect 1066 112325 116786 112891
rect 1066 111237 116786 111803
rect 1066 110149 116786 110715
rect 1066 109061 116786 109627
rect 1066 107973 116786 108539
rect 1066 106885 116786 107451
rect 1066 105797 116786 106363
rect 1066 104709 116786 105275
rect 1066 103621 116786 104187
rect 1066 102533 116786 103099
rect 1066 101445 116786 102011
rect 1066 100357 116786 100923
rect 1066 99269 116786 99835
rect 1066 98181 116786 98747
rect 1066 97093 116786 97659
rect 1066 96005 116786 96571
rect 1066 94917 116786 95483
rect 1066 93829 116786 94395
rect 1066 92741 116786 93307
rect 1066 91653 116786 92219
rect 1066 90565 116786 91131
rect 1066 89477 116786 90043
rect 1066 88389 116786 88955
rect 1066 87301 116786 87867
rect 1066 86213 116786 86779
rect 1066 85125 116786 85691
rect 1066 84037 116786 84603
rect 1066 82949 116786 83515
rect 1066 81861 116786 82427
rect 1066 80773 116786 81339
rect 1066 79685 116786 80251
rect 1066 78597 116786 79163
rect 1066 77509 116786 78075
rect 1066 76421 116786 76987
rect 1066 75333 116786 75899
rect 1066 74245 116786 74811
rect 1066 73157 116786 73723
rect 1066 72069 116786 72635
rect 1066 70981 116786 71547
rect 1066 69893 116786 70459
rect 1066 68805 116786 69371
rect 1066 67717 116786 68283
rect 1066 66629 116786 67195
rect 1066 65541 116786 66107
rect 1066 64453 116786 65019
rect 1066 63365 116786 63931
rect 1066 62277 116786 62843
rect 1066 61189 116786 61755
rect 1066 60101 116786 60667
rect 1066 59013 116786 59579
rect 1066 57925 116786 58491
rect 1066 56837 116786 57403
rect 1066 55749 116786 56315
rect 1066 54661 116786 55227
rect 1066 53573 116786 54139
rect 1066 52485 116786 53051
rect 1066 51397 116786 51963
rect 1066 50309 116786 50875
rect 1066 49221 116786 49787
rect 1066 48133 116786 48699
rect 1066 47045 116786 47611
rect 1066 45957 116786 46523
rect 1066 44869 116786 45435
rect 1066 43781 116786 44347
rect 1066 42693 116786 43259
rect 1066 41605 116786 42171
rect 1066 40517 116786 41083
rect 1066 39429 116786 39995
rect 1066 38341 116786 38907
rect 1066 37253 116786 37819
rect 1066 36165 116786 36731
rect 1066 35077 116786 35643
rect 1066 33989 116786 34555
rect 1066 32901 116786 33467
rect 1066 31813 116786 32379
rect 1066 30725 116786 31291
rect 1066 29637 116786 30203
rect 1066 28549 116786 29115
rect 1066 27461 116786 28027
rect 1066 26373 116786 26939
rect 1066 25285 116786 25851
rect 1066 24197 116786 24763
rect 1066 23109 116786 23675
rect 1066 22021 116786 22587
rect 1066 20933 116786 21499
rect 1066 19845 116786 20411
rect 1066 18757 116786 19323
rect 1066 17669 116786 18235
rect 1066 16581 116786 17147
rect 1066 15493 116786 16059
rect 1066 14405 116786 14971
rect 1066 13317 116786 13883
rect 1066 12229 116786 12795
rect 1066 11141 116786 11707
rect 1066 10053 116786 10619
rect 1066 8965 116786 9531
rect 1066 7877 116786 8443
rect 1066 6789 116786 7355
rect 1066 5701 116786 6267
rect 1066 4613 116786 5179
rect 1066 3525 116786 4091
rect 1066 2437 116786 3003
<< obsli1 >>
rect 1104 2159 116748 117521
<< obsm1 >>
rect 1104 1912 116748 117552
<< metal2 >>
rect 1490 119265 1546 120065
rect 3882 119265 3938 120065
rect 6274 119265 6330 120065
rect 8666 119265 8722 120065
rect 11058 119265 11114 120065
rect 13450 119265 13506 120065
rect 15842 119265 15898 120065
rect 18234 119265 18290 120065
rect 20626 119265 20682 120065
rect 23018 119265 23074 120065
rect 25410 119265 25466 120065
rect 27802 119265 27858 120065
rect 30194 119265 30250 120065
rect 32586 119265 32642 120065
rect 34978 119265 35034 120065
rect 37370 119265 37426 120065
rect 39762 119265 39818 120065
rect 42154 119265 42210 120065
rect 44546 119265 44602 120065
rect 46938 119265 46994 120065
rect 49330 119265 49386 120065
rect 51722 119265 51778 120065
rect 54114 119265 54170 120065
rect 56506 119265 56562 120065
rect 58898 119265 58954 120065
rect 61290 119265 61346 120065
rect 63682 119265 63738 120065
rect 66074 119265 66130 120065
rect 68466 119265 68522 120065
rect 70858 119265 70914 120065
rect 73250 119265 73306 120065
rect 75642 119265 75698 120065
rect 78034 119265 78090 120065
rect 80426 119265 80482 120065
rect 82818 119265 82874 120065
rect 85210 119265 85266 120065
rect 87602 119265 87658 120065
rect 89994 119265 90050 120065
rect 92386 119265 92442 120065
rect 94778 119265 94834 120065
rect 97170 119265 97226 120065
rect 99562 119265 99618 120065
rect 101954 119265 102010 120065
rect 104346 119265 104402 120065
rect 106738 119265 106794 120065
rect 109130 119265 109186 120065
rect 111522 119265 111578 120065
rect 113914 119265 113970 120065
rect 116306 119265 116362 120065
rect 2962 0 3018 800
rect 5906 0 5962 800
rect 8850 0 8906 800
rect 11794 0 11850 800
rect 14738 0 14794 800
rect 17682 0 17738 800
rect 20626 0 20682 800
rect 23570 0 23626 800
rect 26514 0 26570 800
rect 29458 0 29514 800
rect 32402 0 32458 800
rect 35346 0 35402 800
rect 38290 0 38346 800
rect 41234 0 41290 800
rect 44178 0 44234 800
rect 47122 0 47178 800
rect 50066 0 50122 800
rect 53010 0 53066 800
rect 55954 0 56010 800
rect 58898 0 58954 800
rect 61842 0 61898 800
rect 64786 0 64842 800
rect 67730 0 67786 800
rect 70674 0 70730 800
rect 73618 0 73674 800
rect 76562 0 76618 800
rect 79506 0 79562 800
rect 82450 0 82506 800
rect 85394 0 85450 800
rect 88338 0 88394 800
rect 91282 0 91338 800
rect 94226 0 94282 800
rect 97170 0 97226 800
rect 100114 0 100170 800
rect 103058 0 103114 800
rect 106002 0 106058 800
rect 108946 0 109002 800
rect 111890 0 111946 800
rect 114834 0 114890 800
<< obsm2 >>
rect 1602 119209 3826 119265
rect 3994 119209 6218 119265
rect 6386 119209 8610 119265
rect 8778 119209 11002 119265
rect 11170 119209 13394 119265
rect 13562 119209 15786 119265
rect 15954 119209 18178 119265
rect 18346 119209 20570 119265
rect 20738 119209 22962 119265
rect 23130 119209 25354 119265
rect 25522 119209 27746 119265
rect 27914 119209 30138 119265
rect 30306 119209 32530 119265
rect 32698 119209 34922 119265
rect 35090 119209 37314 119265
rect 37482 119209 39706 119265
rect 39874 119209 42098 119265
rect 42266 119209 44490 119265
rect 44658 119209 46882 119265
rect 47050 119209 49274 119265
rect 49442 119209 51666 119265
rect 51834 119209 54058 119265
rect 54226 119209 56450 119265
rect 56618 119209 58842 119265
rect 59010 119209 61234 119265
rect 61402 119209 63626 119265
rect 63794 119209 66018 119265
rect 66186 119209 68410 119265
rect 68578 119209 70802 119265
rect 70970 119209 73194 119265
rect 73362 119209 75586 119265
rect 75754 119209 77978 119265
rect 78146 119209 80370 119265
rect 80538 119209 82762 119265
rect 82930 119209 85154 119265
rect 85322 119209 87546 119265
rect 87714 119209 89938 119265
rect 90106 119209 92330 119265
rect 92498 119209 94722 119265
rect 94890 119209 97114 119265
rect 97282 119209 99506 119265
rect 99674 119209 101898 119265
rect 102066 119209 104290 119265
rect 104458 119209 106682 119265
rect 106850 119209 109074 119265
rect 109242 119209 111466 119265
rect 111634 119209 113858 119265
rect 114026 119209 116250 119265
rect 116418 119209 116636 119265
rect 1584 856 116636 119209
rect 1584 800 2906 856
rect 3074 800 5850 856
rect 6018 800 8794 856
rect 8962 800 11738 856
rect 11906 800 14682 856
rect 14850 800 17626 856
rect 17794 800 20570 856
rect 20738 800 23514 856
rect 23682 800 26458 856
rect 26626 800 29402 856
rect 29570 800 32346 856
rect 32514 800 35290 856
rect 35458 800 38234 856
rect 38402 800 41178 856
rect 41346 800 44122 856
rect 44290 800 47066 856
rect 47234 800 50010 856
rect 50178 800 52954 856
rect 53122 800 55898 856
rect 56066 800 58842 856
rect 59010 800 61786 856
rect 61954 800 64730 856
rect 64898 800 67674 856
rect 67842 800 70618 856
rect 70786 800 73562 856
rect 73730 800 76506 856
rect 76674 800 79450 856
rect 79618 800 82394 856
rect 82562 800 85338 856
rect 85506 800 88282 856
rect 88450 800 91226 856
rect 91394 800 94170 856
rect 94338 800 97114 856
rect 97282 800 100058 856
rect 100226 800 103002 856
rect 103170 800 105946 856
rect 106114 800 108890 856
rect 109058 800 111834 856
rect 112002 800 114778 856
rect 114946 800 116636 856
<< metal3 >>
rect 117121 117104 117921 117224
rect 117121 114248 117921 114368
rect 117121 111392 117921 111512
rect 117121 108536 117921 108656
rect 117121 105680 117921 105800
rect 117121 102824 117921 102944
rect 117121 99968 117921 100088
rect 117121 97112 117921 97232
rect 117121 94256 117921 94376
rect 117121 91400 117921 91520
rect 117121 88544 117921 88664
rect 117121 85688 117921 85808
rect 117121 82832 117921 82952
rect 117121 79976 117921 80096
rect 117121 77120 117921 77240
rect 117121 74264 117921 74384
rect 117121 71408 117921 71528
rect 117121 68552 117921 68672
rect 117121 65696 117921 65816
rect 117121 62840 117921 62960
rect 117121 59984 117921 60104
rect 117121 57128 117921 57248
rect 117121 54272 117921 54392
rect 117121 51416 117921 51536
rect 117121 48560 117921 48680
rect 117121 45704 117921 45824
rect 117121 42848 117921 42968
rect 117121 39992 117921 40112
rect 117121 37136 117921 37256
rect 117121 34280 117921 34400
rect 117121 31424 117921 31544
rect 117121 28568 117921 28688
rect 117121 25712 117921 25832
rect 117121 22856 117921 22976
rect 117121 20000 117921 20120
rect 117121 17144 117921 17264
rect 117121 14288 117921 14408
rect 117121 11432 117921 11552
rect 117121 8576 117921 8696
rect 117121 5720 117921 5840
rect 117121 2864 117921 2984
<< obsm3 >>
rect 4210 117304 117121 117537
rect 4210 117024 117041 117304
rect 4210 114448 117121 117024
rect 4210 114168 117041 114448
rect 4210 111592 117121 114168
rect 4210 111312 117041 111592
rect 4210 108736 117121 111312
rect 4210 108456 117041 108736
rect 4210 105880 117121 108456
rect 4210 105600 117041 105880
rect 4210 103024 117121 105600
rect 4210 102744 117041 103024
rect 4210 100168 117121 102744
rect 4210 99888 117041 100168
rect 4210 97312 117121 99888
rect 4210 97032 117041 97312
rect 4210 94456 117121 97032
rect 4210 94176 117041 94456
rect 4210 91600 117121 94176
rect 4210 91320 117041 91600
rect 4210 88744 117121 91320
rect 4210 88464 117041 88744
rect 4210 85888 117121 88464
rect 4210 85608 117041 85888
rect 4210 83032 117121 85608
rect 4210 82752 117041 83032
rect 4210 80176 117121 82752
rect 4210 79896 117041 80176
rect 4210 77320 117121 79896
rect 4210 77040 117041 77320
rect 4210 74464 117121 77040
rect 4210 74184 117041 74464
rect 4210 71608 117121 74184
rect 4210 71328 117041 71608
rect 4210 68752 117121 71328
rect 4210 68472 117041 68752
rect 4210 65896 117121 68472
rect 4210 65616 117041 65896
rect 4210 63040 117121 65616
rect 4210 62760 117041 63040
rect 4210 60184 117121 62760
rect 4210 59904 117041 60184
rect 4210 57328 117121 59904
rect 4210 57048 117041 57328
rect 4210 54472 117121 57048
rect 4210 54192 117041 54472
rect 4210 51616 117121 54192
rect 4210 51336 117041 51616
rect 4210 48760 117121 51336
rect 4210 48480 117041 48760
rect 4210 45904 117121 48480
rect 4210 45624 117041 45904
rect 4210 43048 117121 45624
rect 4210 42768 117041 43048
rect 4210 40192 117121 42768
rect 4210 39912 117041 40192
rect 4210 37336 117121 39912
rect 4210 37056 117041 37336
rect 4210 34480 117121 37056
rect 4210 34200 117041 34480
rect 4210 31624 117121 34200
rect 4210 31344 117041 31624
rect 4210 28768 117121 31344
rect 4210 28488 117041 28768
rect 4210 25912 117121 28488
rect 4210 25632 117041 25912
rect 4210 23056 117121 25632
rect 4210 22776 117041 23056
rect 4210 20200 117121 22776
rect 4210 19920 117041 20200
rect 4210 17344 117121 19920
rect 4210 17064 117041 17344
rect 4210 14488 117121 17064
rect 4210 14208 117041 14488
rect 4210 11632 117121 14208
rect 4210 11352 117041 11632
rect 4210 8776 117121 11352
rect 4210 8496 117041 8776
rect 4210 5920 117121 8496
rect 4210 5640 117041 5920
rect 4210 3064 117121 5640
rect 4210 2784 117041 3064
rect 4210 1803 117121 2784
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 14963 2048 19488 117061
rect 19968 2048 34848 117061
rect 35328 2048 50208 117061
rect 50688 2048 65568 117061
rect 66048 2048 80928 117061
rect 81408 2048 96288 117061
rect 96768 2048 104637 117061
rect 14963 1803 104637 2048
<< labels >>
rlabel metal3 s 117121 2864 117921 2984 6 i_clk
port 1 nsew signal input
rlabel metal3 s 117121 71408 117921 71528 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 117121 51416 117921 51536 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 117121 17144 117921 17264 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 117121 20000 117921 20120 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 117121 22856 117921 22976 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 117121 25712 117921 25832 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 117121 28568 117921 28688 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 117121 31424 117921 31544 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 117121 34280 117921 34400 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 117121 37136 117921 37256 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 117121 39992 117921 40112 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 117121 42848 117921 42968 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 117121 45704 117921 45824 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 117121 48560 117921 48680 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 117121 54272 117921 54392 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 117121 57128 117921 57248 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 117121 59984 117921 60104 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 117121 62840 117921 62960 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 117121 65696 117921 65816 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 117121 68552 117921 68672 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 117121 74264 117921 74384 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 117121 77120 117921 77240 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 117121 79976 117921 80096 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 117121 82832 117921 82952 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 117121 85688 117921 85808 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 117121 88544 117921 88664 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 117121 91400 117921 91520 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 117121 94256 117921 94376 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 117121 97112 117921 97232 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 117121 99968 117921 100088 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 117121 102824 117921 102944 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 117121 105680 117921 105800 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 117121 108536 117921 108656 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 117121 111392 117921 111512 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 117121 114248 117921 114368 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 117121 5720 117921 5840 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 117121 8576 117921 8696 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 117121 11432 117921 11552 6 i_reg_outs_enb
port 47 nsew signal input
rlabel metal3 s 117121 14288 117921 14408 6 i_reg_sclk
port 48 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 i_reset_lock_a
port 49 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 i_reset_lock_b
port 50 nsew signal input
rlabel metal3 s 117121 117104 117921 117224 6 i_spare_0
port 51 nsew signal input
rlabel metal2 s 1490 119265 1546 120065 6 i_spare_1
port 52 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 i_test_wb_clk_i
port 53 nsew signal input
rlabel metal2 s 11058 119265 11114 120065 6 i_tex_in[0]
port 54 nsew signal input
rlabel metal2 s 8666 119265 8722 120065 6 i_tex_in[1]
port 55 nsew signal input
rlabel metal2 s 6274 119265 6330 120065 6 i_tex_in[2]
port 56 nsew signal input
rlabel metal2 s 3882 119265 3938 120065 6 i_tex_in[3]
port 57 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 i_vec_csb
port 58 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 i_vec_mosi
port 59 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 i_vec_sclk
port 60 nsew signal input
rlabel metal2 s 25410 119265 25466 120065 6 o_gpout[0]
port 61 nsew signal output
rlabel metal2 s 23018 119265 23074 120065 6 o_gpout[1]
port 62 nsew signal output
rlabel metal2 s 20626 119265 20682 120065 6 o_gpout[2]
port 63 nsew signal output
rlabel metal2 s 18234 119265 18290 120065 6 o_gpout[3]
port 64 nsew signal output
rlabel metal2 s 15842 119265 15898 120065 6 o_gpout[4]
port 65 nsew signal output
rlabel metal2 s 13450 119265 13506 120065 6 o_gpout[5]
port 66 nsew signal output
rlabel metal2 s 39762 119265 39818 120065 6 o_hsync
port 67 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 o_reset
port 68 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 o_rgb[0]
port 69 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 o_rgb[10]
port 70 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 o_rgb[11]
port 71 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 o_rgb[12]
port 72 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 o_rgb[13]
port 73 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 o_rgb[14]
port 74 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 o_rgb[15]
port 75 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 o_rgb[16]
port 76 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 o_rgb[17]
port 77 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 o_rgb[18]
port 78 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 o_rgb[19]
port 79 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 o_rgb[1]
port 80 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 o_rgb[20]
port 81 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 o_rgb[21]
port 82 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 o_rgb[22]
port 83 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 o_rgb[23]
port 84 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 o_rgb[2]
port 85 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 o_rgb[3]
port 86 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 o_rgb[4]
port 87 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 o_rgb[5]
port 88 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 o_rgb[6]
port 89 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 o_rgb[7]
port 90 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 o_rgb[8]
port 91 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 o_rgb[9]
port 92 nsew signal output
rlabel metal2 s 34978 119265 35034 120065 6 o_tex_csb
port 93 nsew signal output
rlabel metal2 s 32586 119265 32642 120065 6 o_tex_oeb0
port 94 nsew signal output
rlabel metal2 s 30194 119265 30250 120065 6 o_tex_out0
port 95 nsew signal output
rlabel metal2 s 27802 119265 27858 120065 6 o_tex_sclk
port 96 nsew signal output
rlabel metal2 s 37370 119265 37426 120065 6 o_vsync
port 97 nsew signal output
rlabel metal2 s 116306 119265 116362 120065 6 ones[0]
port 98 nsew signal output
rlabel metal2 s 92386 119265 92442 120065 6 ones[10]
port 99 nsew signal output
rlabel metal2 s 89994 119265 90050 120065 6 ones[11]
port 100 nsew signal output
rlabel metal2 s 87602 119265 87658 120065 6 ones[12]
port 101 nsew signal output
rlabel metal2 s 85210 119265 85266 120065 6 ones[13]
port 102 nsew signal output
rlabel metal2 s 82818 119265 82874 120065 6 ones[14]
port 103 nsew signal output
rlabel metal2 s 80426 119265 80482 120065 6 ones[15]
port 104 nsew signal output
rlabel metal2 s 113914 119265 113970 120065 6 ones[1]
port 105 nsew signal output
rlabel metal2 s 111522 119265 111578 120065 6 ones[2]
port 106 nsew signal output
rlabel metal2 s 109130 119265 109186 120065 6 ones[3]
port 107 nsew signal output
rlabel metal2 s 106738 119265 106794 120065 6 ones[4]
port 108 nsew signal output
rlabel metal2 s 104346 119265 104402 120065 6 ones[5]
port 109 nsew signal output
rlabel metal2 s 101954 119265 102010 120065 6 ones[6]
port 110 nsew signal output
rlabel metal2 s 99562 119265 99618 120065 6 ones[7]
port 111 nsew signal output
rlabel metal2 s 97170 119265 97226 120065 6 ones[8]
port 112 nsew signal output
rlabel metal2 s 94778 119265 94834 120065 6 ones[9]
port 113 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 115 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 115 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 115 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 115 nsew ground bidirectional
rlabel metal2 s 78034 119265 78090 120065 6 zeros[0]
port 116 nsew signal output
rlabel metal2 s 54114 119265 54170 120065 6 zeros[10]
port 117 nsew signal output
rlabel metal2 s 51722 119265 51778 120065 6 zeros[11]
port 118 nsew signal output
rlabel metal2 s 49330 119265 49386 120065 6 zeros[12]
port 119 nsew signal output
rlabel metal2 s 46938 119265 46994 120065 6 zeros[13]
port 120 nsew signal output
rlabel metal2 s 44546 119265 44602 120065 6 zeros[14]
port 121 nsew signal output
rlabel metal2 s 42154 119265 42210 120065 6 zeros[15]
port 122 nsew signal output
rlabel metal2 s 75642 119265 75698 120065 6 zeros[1]
port 123 nsew signal output
rlabel metal2 s 73250 119265 73306 120065 6 zeros[2]
port 124 nsew signal output
rlabel metal2 s 70858 119265 70914 120065 6 zeros[3]
port 125 nsew signal output
rlabel metal2 s 68466 119265 68522 120065 6 zeros[4]
port 126 nsew signal output
rlabel metal2 s 66074 119265 66130 120065 6 zeros[5]
port 127 nsew signal output
rlabel metal2 s 63682 119265 63738 120065 6 zeros[6]
port 128 nsew signal output
rlabel metal2 s 61290 119265 61346 120065 6 zeros[7]
port 129 nsew signal output
rlabel metal2 s 58898 119265 58954 120065 6 zeros[8]
port 130 nsew signal output
rlabel metal2 s 56506 119265 56562 120065 6 zeros[9]
port 131 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 117921 120065
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 33014132
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/top_ew_algofoogle/runs/23_11_04_21_36/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1418004
<< end >>

