magic
tech sky130A
magscale 1 2
timestamp 1699030802
<< nwell >>
rect 1066 116677 116326 116998
rect 1066 115589 116326 116155
rect 1066 114501 116326 115067
rect 1066 113413 116326 113979
rect 1066 112325 116326 112891
rect 1066 111237 116326 111803
rect 1066 110149 116326 110715
rect 1066 109061 116326 109627
rect 1066 107973 116326 108539
rect 1066 106885 116326 107451
rect 1066 105797 116326 106363
rect 1066 104709 116326 105275
rect 1066 103621 116326 104187
rect 1066 102533 116326 103099
rect 1066 101445 116326 102011
rect 1066 100357 116326 100923
rect 1066 99269 116326 99835
rect 1066 98181 116326 98747
rect 1066 97093 116326 97659
rect 1066 96005 116326 96571
rect 1066 94917 116326 95483
rect 1066 93829 116326 94395
rect 1066 92741 116326 93307
rect 1066 91653 116326 92219
rect 1066 90565 116326 91131
rect 1066 89477 116326 90043
rect 1066 88389 116326 88955
rect 1066 87301 116326 87867
rect 1066 86213 116326 86779
rect 1066 85125 116326 85691
rect 1066 84037 116326 84603
rect 1066 82949 116326 83515
rect 1066 81861 116326 82427
rect 1066 80773 116326 81339
rect 1066 79685 116326 80251
rect 1066 78597 116326 79163
rect 1066 77509 116326 78075
rect 1066 76421 116326 76987
rect 1066 75333 116326 75899
rect 1066 74245 116326 74811
rect 1066 73157 116326 73723
rect 1066 72069 116326 72635
rect 1066 70981 116326 71547
rect 1066 69893 116326 70459
rect 1066 68805 116326 69371
rect 1066 67717 116326 68283
rect 1066 66629 116326 67195
rect 1066 65541 116326 66107
rect 1066 64453 116326 65019
rect 1066 63365 116326 63931
rect 1066 62277 116326 62843
rect 1066 61189 116326 61755
rect 1066 60101 116326 60667
rect 1066 59013 116326 59579
rect 1066 57925 116326 58491
rect 1066 56837 116326 57403
rect 1066 55749 116326 56315
rect 1066 54661 116326 55227
rect 1066 53573 116326 54139
rect 1066 52485 116326 53051
rect 1066 51397 116326 51963
rect 1066 50309 116326 50875
rect 1066 49221 116326 49787
rect 1066 48133 116326 48699
rect 1066 47045 116326 47611
rect 1066 45957 116326 46523
rect 1066 44869 116326 45435
rect 1066 43781 116326 44347
rect 1066 42693 116326 43259
rect 1066 41605 116326 42171
rect 1066 40517 116326 41083
rect 1066 39429 116326 39995
rect 1066 38341 116326 38907
rect 1066 37253 116326 37819
rect 1066 36165 116326 36731
rect 1066 35077 116326 35643
rect 1066 33989 116326 34555
rect 1066 32901 116326 33467
rect 1066 31813 116326 32379
rect 1066 30725 116326 31291
rect 1066 29637 116326 30203
rect 1066 28549 116326 29115
rect 1066 27461 116326 28027
rect 1066 26373 116326 26939
rect 1066 25285 116326 25851
rect 1066 24197 116326 24763
rect 1066 23109 116326 23675
rect 1066 22021 116326 22587
rect 1066 20933 116326 21499
rect 1066 19845 116326 20411
rect 1066 18757 116326 19323
rect 1066 17669 116326 18235
rect 1066 16581 116326 17147
rect 1066 15493 116326 16059
rect 1066 14405 116326 14971
rect 1066 13317 116326 13883
rect 1066 12229 116326 12795
rect 1066 11141 116326 11707
rect 1066 10053 116326 10619
rect 1066 8965 116326 9531
rect 1066 7877 116326 8443
rect 1066 6789 116326 7355
rect 1066 5701 116326 6267
rect 1066 4613 116326 5179
rect 1066 3525 116326 4091
rect 1066 2437 116326 3003
<< obsli1 >>
rect 1104 2159 116288 116977
<< obsm1 >>
rect 1104 1844 116288 117008
<< metal2 >>
rect 1306 118814 1362 119614
rect 3698 118814 3754 119614
rect 6090 118814 6146 119614
rect 8482 118814 8538 119614
rect 10874 118814 10930 119614
rect 13266 118814 13322 119614
rect 15658 118814 15714 119614
rect 18050 118814 18106 119614
rect 20442 118814 20498 119614
rect 22834 118814 22890 119614
rect 25226 118814 25282 119614
rect 27618 118814 27674 119614
rect 30010 118814 30066 119614
rect 32402 118814 32458 119614
rect 34794 118814 34850 119614
rect 37186 118814 37242 119614
rect 39578 118814 39634 119614
rect 41970 118814 42026 119614
rect 44362 118814 44418 119614
rect 46754 118814 46810 119614
rect 49146 118814 49202 119614
rect 51538 118814 51594 119614
rect 53930 118814 53986 119614
rect 56322 118814 56378 119614
rect 58714 118814 58770 119614
rect 61106 118814 61162 119614
rect 63498 118814 63554 119614
rect 65890 118814 65946 119614
rect 68282 118814 68338 119614
rect 70674 118814 70730 119614
rect 73066 118814 73122 119614
rect 75458 118814 75514 119614
rect 77850 118814 77906 119614
rect 80242 118814 80298 119614
rect 82634 118814 82690 119614
rect 85026 118814 85082 119614
rect 87418 118814 87474 119614
rect 89810 118814 89866 119614
rect 92202 118814 92258 119614
rect 94594 118814 94650 119614
rect 96986 118814 97042 119614
rect 99378 118814 99434 119614
rect 101770 118814 101826 119614
rect 104162 118814 104218 119614
rect 106554 118814 106610 119614
rect 108946 118814 109002 119614
rect 111338 118814 111394 119614
rect 113730 118814 113786 119614
rect 116122 118814 116178 119614
rect 2778 0 2834 800
rect 5722 0 5778 800
rect 8666 0 8722 800
rect 11610 0 11666 800
rect 14554 0 14610 800
rect 17498 0 17554 800
rect 20442 0 20498 800
rect 23386 0 23442 800
rect 26330 0 26386 800
rect 29274 0 29330 800
rect 32218 0 32274 800
rect 35162 0 35218 800
rect 38106 0 38162 800
rect 41050 0 41106 800
rect 43994 0 44050 800
rect 46938 0 46994 800
rect 49882 0 49938 800
rect 52826 0 52882 800
rect 55770 0 55826 800
rect 58714 0 58770 800
rect 61658 0 61714 800
rect 64602 0 64658 800
rect 67546 0 67602 800
rect 70490 0 70546 800
rect 73434 0 73490 800
rect 76378 0 76434 800
rect 79322 0 79378 800
rect 82266 0 82322 800
rect 85210 0 85266 800
rect 88154 0 88210 800
rect 91098 0 91154 800
rect 94042 0 94098 800
rect 96986 0 97042 800
rect 99930 0 99986 800
rect 102874 0 102930 800
rect 105818 0 105874 800
rect 108762 0 108818 800
rect 111706 0 111762 800
rect 114650 0 114706 800
<< obsm2 >>
rect 1860 118758 3642 118946
rect 3810 118758 6034 118946
rect 6202 118758 8426 118946
rect 8594 118758 10818 118946
rect 10986 118758 13210 118946
rect 13378 118758 15602 118946
rect 15770 118758 17994 118946
rect 18162 118758 20386 118946
rect 20554 118758 22778 118946
rect 22946 118758 25170 118946
rect 25338 118758 27562 118946
rect 27730 118758 29954 118946
rect 30122 118758 32346 118946
rect 32514 118758 34738 118946
rect 34906 118758 37130 118946
rect 37298 118758 39522 118946
rect 39690 118758 41914 118946
rect 42082 118758 44306 118946
rect 44474 118758 46698 118946
rect 46866 118758 49090 118946
rect 49258 118758 51482 118946
rect 51650 118758 53874 118946
rect 54042 118758 56266 118946
rect 56434 118758 58658 118946
rect 58826 118758 61050 118946
rect 61218 118758 63442 118946
rect 63610 118758 65834 118946
rect 66002 118758 68226 118946
rect 68394 118758 70618 118946
rect 70786 118758 73010 118946
rect 73178 118758 75402 118946
rect 75570 118758 77794 118946
rect 77962 118758 80186 118946
rect 80354 118758 82578 118946
rect 82746 118758 84970 118946
rect 85138 118758 87362 118946
rect 87530 118758 89754 118946
rect 89922 118758 92146 118946
rect 92314 118758 94538 118946
rect 94706 118758 96930 118946
rect 97098 118758 99322 118946
rect 99490 118758 101714 118946
rect 101882 118758 104106 118946
rect 104274 118758 106498 118946
rect 106666 118758 108890 118946
rect 109058 118758 111282 118946
rect 111450 118758 113674 118946
rect 113842 118758 116066 118946
rect 1860 856 116176 118758
rect 1860 800 2722 856
rect 2890 800 5666 856
rect 5834 800 8610 856
rect 8778 800 11554 856
rect 11722 800 14498 856
rect 14666 800 17442 856
rect 17610 800 20386 856
rect 20554 800 23330 856
rect 23498 800 26274 856
rect 26442 800 29218 856
rect 29386 800 32162 856
rect 32330 800 35106 856
rect 35274 800 38050 856
rect 38218 800 40994 856
rect 41162 800 43938 856
rect 44106 800 46882 856
rect 47050 800 49826 856
rect 49994 800 52770 856
rect 52938 800 55714 856
rect 55882 800 58658 856
rect 58826 800 61602 856
rect 61770 800 64546 856
rect 64714 800 67490 856
rect 67658 800 70434 856
rect 70602 800 73378 856
rect 73546 800 76322 856
rect 76490 800 79266 856
rect 79434 800 82210 856
rect 82378 800 85154 856
rect 85322 800 88098 856
rect 88266 800 91042 856
rect 91210 800 93986 856
rect 94154 800 96930 856
rect 97098 800 99874 856
rect 100042 800 102818 856
rect 102986 800 105762 856
rect 105930 800 108706 856
rect 108874 800 111650 856
rect 111818 800 114594 856
rect 114762 800 116176 856
<< metal3 >>
rect 116670 116832 117470 116952
rect 116670 113976 117470 114096
rect 116670 111120 117470 111240
rect 116670 108264 117470 108384
rect 116670 105408 117470 105528
rect 116670 102552 117470 102672
rect 116670 99696 117470 99816
rect 116670 96840 117470 96960
rect 116670 93984 117470 94104
rect 116670 91128 117470 91248
rect 116670 88272 117470 88392
rect 116670 85416 117470 85536
rect 116670 82560 117470 82680
rect 116670 79704 117470 79824
rect 116670 76848 117470 76968
rect 116670 73992 117470 74112
rect 116670 71136 117470 71256
rect 116670 68280 117470 68400
rect 116670 65424 117470 65544
rect 116670 62568 117470 62688
rect 116670 59712 117470 59832
rect 116670 56856 117470 56976
rect 116670 54000 117470 54120
rect 116670 51144 117470 51264
rect 116670 48288 117470 48408
rect 116670 45432 117470 45552
rect 116670 42576 117470 42696
rect 116670 39720 117470 39840
rect 116670 36864 117470 36984
rect 116670 34008 117470 34128
rect 116670 31152 117470 31272
rect 116670 28296 117470 28416
rect 116670 25440 117470 25560
rect 116670 22584 117470 22704
rect 116670 19728 117470 19848
rect 116670 16872 117470 16992
rect 116670 14016 117470 14136
rect 116670 11160 117470 11280
rect 116670 8304 117470 8424
rect 116670 5448 117470 5568
rect 116670 2592 117470 2712
<< obsm3 >>
rect 4210 116752 116590 116993
rect 4210 114176 116670 116752
rect 4210 113896 116590 114176
rect 4210 111320 116670 113896
rect 4210 111040 116590 111320
rect 4210 108464 116670 111040
rect 4210 108184 116590 108464
rect 4210 105608 116670 108184
rect 4210 105328 116590 105608
rect 4210 102752 116670 105328
rect 4210 102472 116590 102752
rect 4210 99896 116670 102472
rect 4210 99616 116590 99896
rect 4210 97040 116670 99616
rect 4210 96760 116590 97040
rect 4210 94184 116670 96760
rect 4210 93904 116590 94184
rect 4210 91328 116670 93904
rect 4210 91048 116590 91328
rect 4210 88472 116670 91048
rect 4210 88192 116590 88472
rect 4210 85616 116670 88192
rect 4210 85336 116590 85616
rect 4210 82760 116670 85336
rect 4210 82480 116590 82760
rect 4210 79904 116670 82480
rect 4210 79624 116590 79904
rect 4210 77048 116670 79624
rect 4210 76768 116590 77048
rect 4210 74192 116670 76768
rect 4210 73912 116590 74192
rect 4210 71336 116670 73912
rect 4210 71056 116590 71336
rect 4210 68480 116670 71056
rect 4210 68200 116590 68480
rect 4210 65624 116670 68200
rect 4210 65344 116590 65624
rect 4210 62768 116670 65344
rect 4210 62488 116590 62768
rect 4210 59912 116670 62488
rect 4210 59632 116590 59912
rect 4210 57056 116670 59632
rect 4210 56776 116590 57056
rect 4210 54200 116670 56776
rect 4210 53920 116590 54200
rect 4210 51344 116670 53920
rect 4210 51064 116590 51344
rect 4210 48488 116670 51064
rect 4210 48208 116590 48488
rect 4210 45632 116670 48208
rect 4210 45352 116590 45632
rect 4210 42776 116670 45352
rect 4210 42496 116590 42776
rect 4210 39920 116670 42496
rect 4210 39640 116590 39920
rect 4210 37064 116670 39640
rect 4210 36784 116590 37064
rect 4210 34208 116670 36784
rect 4210 33928 116590 34208
rect 4210 31352 116670 33928
rect 4210 31072 116590 31352
rect 4210 28496 116670 31072
rect 4210 28216 116590 28496
rect 4210 25640 116670 28216
rect 4210 25360 116590 25640
rect 4210 22784 116670 25360
rect 4210 22504 116590 22784
rect 4210 19928 116670 22504
rect 4210 19648 116590 19928
rect 4210 17072 116670 19648
rect 4210 16792 116590 17072
rect 4210 14216 116670 16792
rect 4210 13936 116590 14216
rect 4210 11360 116670 13936
rect 4210 11080 116590 11360
rect 4210 8504 116670 11080
rect 4210 8224 116590 8504
rect 4210 5648 116670 8224
rect 4210 5368 116590 5648
rect 4210 2792 116670 5368
rect 4210 2512 116590 2792
rect 4210 2143 116670 2512
<< metal4 >>
rect 4208 2128 4528 117008
rect 19568 2128 19888 117008
rect 34928 2128 35248 117008
rect 50288 2128 50608 117008
rect 65648 2128 65968 117008
rect 81008 2128 81328 117008
rect 96368 2128 96688 117008
rect 111728 2128 112048 117008
<< obsm4 >>
rect 9259 2347 19488 116109
rect 19968 2347 34848 116109
rect 35328 2347 50208 116109
rect 50688 2347 65568 116109
rect 66048 2347 80928 116109
rect 81408 2347 96288 116109
rect 96768 2347 111648 116109
rect 112128 2347 115309 116109
<< labels >>
rlabel metal3 s 116670 2592 117470 2712 6 i_clk
port 1 nsew signal input
rlabel metal3 s 116670 71136 117470 71256 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 116670 51144 117470 51264 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 116670 16872 117470 16992 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 116670 19728 117470 19848 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 116670 22584 117470 22704 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 116670 25440 117470 25560 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 116670 28296 117470 28416 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 116670 31152 117470 31272 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 116670 34008 117470 34128 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 116670 36864 117470 36984 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 116670 39720 117470 39840 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 116670 42576 117470 42696 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 116670 45432 117470 45552 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 116670 48288 117470 48408 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 116670 54000 117470 54120 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 116670 56856 117470 56976 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 116670 59712 117470 59832 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 116670 62568 117470 62688 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 116670 65424 117470 65544 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 116670 68280 117470 68400 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 116670 73992 117470 74112 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 116670 76848 117470 76968 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 116670 79704 117470 79824 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 116670 82560 117470 82680 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 116670 85416 117470 85536 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 116670 88272 117470 88392 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 116670 91128 117470 91248 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 116670 93984 117470 94104 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 116670 96840 117470 96960 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 116670 99696 117470 99816 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 116670 102552 117470 102672 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 116670 105408 117470 105528 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 116670 108264 117470 108384 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 116670 111120 117470 111240 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 116670 113976 117470 114096 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 116670 5448 117470 5568 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 116670 8304 117470 8424 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 116670 11160 117470 11280 6 i_reg_outs_enb
port 47 nsew signal input
rlabel metal3 s 116670 14016 117470 14136 6 i_reg_sclk
port 48 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 i_reset_lock_a
port 49 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 i_reset_lock_b
port 50 nsew signal input
rlabel metal3 s 116670 116832 117470 116952 6 i_spare_0
port 51 nsew signal input
rlabel metal2 s 1306 118814 1362 119614 6 i_spare_1
port 52 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 i_test_wb_clk_i
port 53 nsew signal input
rlabel metal2 s 10874 118814 10930 119614 6 i_tex_in[0]
port 54 nsew signal input
rlabel metal2 s 8482 118814 8538 119614 6 i_tex_in[1]
port 55 nsew signal input
rlabel metal2 s 6090 118814 6146 119614 6 i_tex_in[2]
port 56 nsew signal input
rlabel metal2 s 3698 118814 3754 119614 6 i_tex_in[3]
port 57 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 i_vec_csb
port 58 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 i_vec_mosi
port 59 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 i_vec_sclk
port 60 nsew signal input
rlabel metal2 s 25226 118814 25282 119614 6 o_gpout[0]
port 61 nsew signal output
rlabel metal2 s 22834 118814 22890 119614 6 o_gpout[1]
port 62 nsew signal output
rlabel metal2 s 20442 118814 20498 119614 6 o_gpout[2]
port 63 nsew signal output
rlabel metal2 s 18050 118814 18106 119614 6 o_gpout[3]
port 64 nsew signal output
rlabel metal2 s 15658 118814 15714 119614 6 o_gpout[4]
port 65 nsew signal output
rlabel metal2 s 13266 118814 13322 119614 6 o_gpout[5]
port 66 nsew signal output
rlabel metal2 s 39578 118814 39634 119614 6 o_hsync
port 67 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 o_reset
port 68 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 o_rgb[0]
port 69 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 o_rgb[10]
port 70 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 o_rgb[11]
port 71 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 o_rgb[12]
port 72 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 o_rgb[13]
port 73 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 o_rgb[14]
port 74 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 o_rgb[15]
port 75 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 o_rgb[16]
port 76 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 o_rgb[17]
port 77 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 o_rgb[18]
port 78 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 o_rgb[19]
port 79 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 o_rgb[1]
port 80 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 o_rgb[20]
port 81 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 o_rgb[21]
port 82 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 o_rgb[22]
port 83 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 o_rgb[23]
port 84 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 o_rgb[2]
port 85 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 o_rgb[3]
port 86 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 o_rgb[4]
port 87 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 o_rgb[5]
port 88 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 o_rgb[6]
port 89 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 o_rgb[7]
port 90 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 o_rgb[8]
port 91 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 o_rgb[9]
port 92 nsew signal output
rlabel metal2 s 34794 118814 34850 119614 6 o_tex_csb
port 93 nsew signal output
rlabel metal2 s 32402 118814 32458 119614 6 o_tex_oeb0
port 94 nsew signal output
rlabel metal2 s 30010 118814 30066 119614 6 o_tex_out0
port 95 nsew signal output
rlabel metal2 s 27618 118814 27674 119614 6 o_tex_sclk
port 96 nsew signal output
rlabel metal2 s 37186 118814 37242 119614 6 o_vsync
port 97 nsew signal output
rlabel metal2 s 116122 118814 116178 119614 6 ones[0]
port 98 nsew signal output
rlabel metal2 s 92202 118814 92258 119614 6 ones[10]
port 99 nsew signal output
rlabel metal2 s 89810 118814 89866 119614 6 ones[11]
port 100 nsew signal output
rlabel metal2 s 87418 118814 87474 119614 6 ones[12]
port 101 nsew signal output
rlabel metal2 s 85026 118814 85082 119614 6 ones[13]
port 102 nsew signal output
rlabel metal2 s 82634 118814 82690 119614 6 ones[14]
port 103 nsew signal output
rlabel metal2 s 80242 118814 80298 119614 6 ones[15]
port 104 nsew signal output
rlabel metal2 s 113730 118814 113786 119614 6 ones[1]
port 105 nsew signal output
rlabel metal2 s 111338 118814 111394 119614 6 ones[2]
port 106 nsew signal output
rlabel metal2 s 108946 118814 109002 119614 6 ones[3]
port 107 nsew signal output
rlabel metal2 s 106554 118814 106610 119614 6 ones[4]
port 108 nsew signal output
rlabel metal2 s 104162 118814 104218 119614 6 ones[5]
port 109 nsew signal output
rlabel metal2 s 101770 118814 101826 119614 6 ones[6]
port 110 nsew signal output
rlabel metal2 s 99378 118814 99434 119614 6 ones[7]
port 111 nsew signal output
rlabel metal2 s 96986 118814 97042 119614 6 ones[8]
port 112 nsew signal output
rlabel metal2 s 94594 118814 94650 119614 6 ones[9]
port 113 nsew signal output
rlabel metal4 s 4208 2128 4528 117008 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117008 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117008 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117008 6 vccd1
port 114 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117008 6 vssd1
port 115 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117008 6 vssd1
port 115 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117008 6 vssd1
port 115 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117008 6 vssd1
port 115 nsew ground bidirectional
rlabel metal2 s 77850 118814 77906 119614 6 zeros[0]
port 116 nsew signal output
rlabel metal2 s 53930 118814 53986 119614 6 zeros[10]
port 117 nsew signal output
rlabel metal2 s 51538 118814 51594 119614 6 zeros[11]
port 118 nsew signal output
rlabel metal2 s 49146 118814 49202 119614 6 zeros[12]
port 119 nsew signal output
rlabel metal2 s 46754 118814 46810 119614 6 zeros[13]
port 120 nsew signal output
rlabel metal2 s 44362 118814 44418 119614 6 zeros[14]
port 121 nsew signal output
rlabel metal2 s 41970 118814 42026 119614 6 zeros[15]
port 122 nsew signal output
rlabel metal2 s 75458 118814 75514 119614 6 zeros[1]
port 123 nsew signal output
rlabel metal2 s 73066 118814 73122 119614 6 zeros[2]
port 124 nsew signal output
rlabel metal2 s 70674 118814 70730 119614 6 zeros[3]
port 125 nsew signal output
rlabel metal2 s 68282 118814 68338 119614 6 zeros[4]
port 126 nsew signal output
rlabel metal2 s 65890 118814 65946 119614 6 zeros[5]
port 127 nsew signal output
rlabel metal2 s 63498 118814 63554 119614 6 zeros[6]
port 128 nsew signal output
rlabel metal2 s 61106 118814 61162 119614 6 zeros[7]
port 129 nsew signal output
rlabel metal2 s 58714 118814 58770 119614 6 zeros[8]
port 130 nsew signal output
rlabel metal2 s 56322 118814 56378 119614 6 zeros[9]
port 131 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 117470 119614
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32892248
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/top_ew_algofoogle/runs/23_11_04_03_24/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1402734
<< end >>

