* NGSPICE file created from top_ew_algofoogle.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt top_ew_algofoogle i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout0_sel[4]
+ i_gpout0_sel[5] i_gpout1_sel[0] i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3]
+ i_gpout1_sel[4] i_gpout1_sel[5] i_gpout2_sel[0] i_gpout2_sel[1] i_gpout2_sel[2]
+ i_gpout2_sel[3] i_gpout2_sel[4] i_gpout2_sel[5] i_gpout3_sel[0] i_gpout3_sel[1]
+ i_gpout3_sel[2] i_gpout3_sel[3] i_gpout3_sel[4] i_gpout3_sel[5] i_gpout4_sel[0]
+ i_gpout4_sel[1] i_gpout4_sel[2] i_gpout4_sel[3] i_gpout4_sel[4] i_gpout4_sel[5]
+ i_gpout5_sel[0] i_gpout5_sel[1] i_gpout5_sel[2] i_gpout5_sel[3] i_gpout5_sel[4]
+ i_gpout5_sel[5] i_la_invalid i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_sclk i_reset_lock_a i_reset_lock_b i_tex_in[0] i_tex_in[1] i_tex_in[2] i_tex_in[3]
+ i_vec_csb i_vec_mosi i_vec_sclk o_gpout[0] o_gpout[1] o_gpout[2] o_gpout[3] o_gpout[4]
+ o_gpout[5] o_hsync o_reset o_rgb[0] o_rgb[10] o_rgb[11] o_rgb[12] o_rgb[13] o_rgb[14]
+ o_rgb[15] o_rgb[16] o_rgb[17] o_rgb[18] o_rgb[19] o_rgb[1] o_rgb[20] o_rgb[21] o_rgb[22]
+ o_rgb[23] o_rgb[2] o_rgb[3] o_rgb[4] o_rgb[5] o_rgb[6] o_rgb[7] o_rgb[8] o_rgb[9]
+ o_tex_csb o_tex_oeb0 o_tex_out0 o_tex_sclk o_vsync ones[0] ones[10] ones[11] ones[12]
+ ones[13] ones[14] ones[15] ones[1] ones[2] ones[3] ones[4] ones[5] ones[6] ones[7]
+ ones[8] ones[9] vccd1 vssd1 zeros[0] zeros[10] zeros[11] zeros[12] zeros[13] zeros[14]
+ zeros[15] zeros[1] zeros[2] zeros[3] zeros[4] zeros[5] zeros[6] zeros[7] zeros[8]
+ zeros[9]
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18869_ rbzero.wall_tracer.trackDistY\[9\] _02542_ _02398_ vssd1 vssd1 vccd1 vccd1
+ _02543_ sky130_fd_sc_hd__mux2_1
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20900_ clknet_leaf_81_i_clk _00669_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20831_ clknet_leaf_91_i_clk _00600_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20762_ clknet_leaf_32_i_clk _00531_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20693_ clknet_leaf_7_i_clk _00477_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21314_ net235 _01083_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21245_ clknet_leaf_64_i_clk _01014_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21176_ clknet_leaf_74_i_clk _00945_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20127_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__buf_1
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11900_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _04290_ vssd1 vssd1 vccd1 vccd1 _04676_
+ sky130_fd_sc_hd__mux2_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ rbzero.wall_tracer.visualWallDist\[-1\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05617_ sky130_fd_sc_hd__a21o_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _04605_ _04606_ _04607_ _04266_ _04229_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__o221a_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _07259_ _07266_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _04129_ vssd1 vssd1 vccd1 vccd1 _04540_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _06201_ _06204_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__or2_1
XFILLER_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ rbzero.tex_g1\[1\] rbzero.tex_g1\[2\] _03691_ vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14481_ _07216_ _07217_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__nor2_2
XFILLER_159_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ rbzero.debug_overlay.vplaneY\[-4\] _04464_ _04460_ rbzero.debug_overlay.vplaneY\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a22o_1
XFILLER_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16220_ _08860_ _08864_ vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__or2_1
X_13432_ _06156_ _06167_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__and2_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ rbzero.tex_g1\[34\] rbzero.tex_g1\[35\] _03658_ vssd1 vssd1 vccd1 vccd1 _03662_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _08795_ _08792_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__xnor2_1
X_13363_ _05823_ _05973_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__or2_1
X_10575_ _03625_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15102_ _07757_ _07758_ _07759_ _07760_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__nand4_2
X_12314_ net27 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16082_ _08283_ _08491_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__or2_1
X_13294_ _05975_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15033_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__nor2_1
X_19910_ rbzero.pov.ready_buffer\[50\] _03141_ _03192_ _03210_ vssd1 vssd1 vccd1 vccd1
+ _03211_ sky130_fd_sc_hd__a211o_1
XFILLER_108_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12245_ net41 _04962_ _04978_ net43 net17 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a221o_1
XFILLER_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12176_ _04907_ net10 _04944_ _04946_ net11 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a311o_1
X_19841_ rbzero.pov.ready_buffer\[64\] _07948_ _03146_ vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11127_ rbzero.wall_tracer.visualWallDist\[8\] rbzero.wall_tracer.visualWallDist\[7\]
+ rbzero.wall_tracer.visualWallDist\[6\] rbzero.wall_tracer.visualWallDist\[5\] vssd1
+ vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or4_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16984_ _09620_ _09623_ vssd1 vssd1 vccd1 vccd1 _09624_ sky130_fd_sc_hd__nand2_1
X_19772_ rbzero.pov.spi_buffer\[59\] rbzero.pov.spi_buffer\[60\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ rbzero.tex_b0\[30\] rbzero.tex_b0\[29\] _03876_ vssd1 vssd1 vccd1 vccd1 _03879_
+ sky130_fd_sc_hd__mux2_1
X_18723_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__nand2_1
X_15935_ _08129_ _08579_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__or2_1
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18654_ _02330_ _02349_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__xnor2_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _08510_ _08466_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__xnor2_4
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14817_ _07487_ _07456_ _07544_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__a21o_1
X_17605_ _10167_ _10170_ vssd1 vssd1 vccd1 vccd1 _10171_ sky130_fd_sc_hd__xnor2_4
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18585_ _02269_ _02270_ _02281_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a21oi_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _08382_ _08388_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__xnor2_2
Xtop_ew_algofoogle_120 vssd1 vssd1 vccd1 vccd1 ones[14] top_ew_algofoogle_120/LO sky130_fd_sc_hd__conb_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17536_ _09126_ _09674_ vssd1 vssd1 vccd1 vccd1 _10102_ sky130_fd_sc_hd__nor2_1
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748_ _05814_ _07472_ _07482_ _07459_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__o211a_1
XFILLER_83_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17467_ _10030_ _10031_ _10029_ _09902_ vssd1 vssd1 vccd1 vccd1 _10034_ sky130_fd_sc_hd__o211a_1
X_14679_ _07343_ _07344_ _07346_ _07378_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__o211a_1
XFILLER_149_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20140__170 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__inv_2
X_16418_ rbzero.debug_overlay.playerY\[-6\] rbzero.debug_overlay.playerX\[-6\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__mux2_1
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19206_ _02750_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17398_ _09670_ _09964_ vssd1 vssd1 vccd1 vccd1 _09965_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19137_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _02704_ sky130_fd_sc_hd__and3_1
XFILLER_160_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ _08991_ _08993_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__xnor2_2
XFILLER_146_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19068_ _02666_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18019_ _10094_ _08423_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_1
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21030_ clknet_leaf_51_i_clk _00799_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20223__245 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__inv_2
X_20814_ clknet_leaf_25_i_clk _00583_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189__389 _04959_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__inv_2
X_20745_ clknet_leaf_36_i_clk _00514_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20676_ clknet_leaf_3_i_clk _00460_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03292_ clknet_0__03292_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03292_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _03510_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ _04140_ _04754_ _04771_ _04787_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o32a_1
X_21228_ clknet_leaf_73_i_clk _00997_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21159_ clknet_leaf_84_i_clk _00928_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13981_ _06716_ _06717_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__nand2_1
XFILLER_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15720_ _08363_ _08364_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__xor2_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12932_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__inv_2
XFILLER_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15651_ _08288_ _08295_ vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__xnor2_2
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _05584_ _05586_ _05587_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__or4b_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _07149_ _07324_ _06176_ _07116_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__a2bb2o_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ rbzero.color_sky\[2\] rbzero.color_floor\[2\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04592_ sky130_fd_sc_hd__mux2_1
X_18370_ _01462_ _09703_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__nand2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _05207_ _08226_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__nor2_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12794_ _05534_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__or2_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_67_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20198__222 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__inv_2
X_17321_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09890_ sky130_fd_sc_hd__nor2_1
X_14533_ _07258_ _07050_ _07052_ _07269_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__o31ai_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ rbzero.tex_g0\[14\] _04356_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__and2_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ rbzero.wall_tracer.trackDistX\[-10\] _09828_ _05414_ vssd1 vssd1 vccd1 vccd1
+ _09829_ sky130_fd_sc_hd__mux2_1
X_14464_ _07151_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__inv_2
X_11676_ _04428_ _04447_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__and2_2
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16203_ _08799_ _08798_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__and2b_1
XFILLER_70_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13415_ _06051_ _06090_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__a21oi_1
XFILLER_168_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17183_ rbzero.traced_texa\[10\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a22o_1
X_10627_ rbzero.tex_g1\[42\] rbzero.tex_g1\[43\] _03647_ vssd1 vssd1 vccd1 vccd1 _03653_
+ sky130_fd_sc_hd__mux2_1
X_14395_ _07130_ _07131_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__nand2_1
XFILLER_167_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _08741_ _08753_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__xnor2_1
X_13346_ _06061_ _06067_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__or2_1
X_10558_ _03616_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16065_ _08701_ _08708_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__nor2_1
XFILLER_115_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13277_ _05986_ _06013_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__xnor2_2
X_10489_ _03557_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15016_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__nand2_1
XFILLER_68_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ net50 _04978_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a21oi_2
XFILLER_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19824_ _02728_ _02820_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__nor2_1
X_12159_ net11 net10 _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and3b_1
XFILLER_64_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19755_ rbzero.pov.spi_buffer\[51\] rbzero.pov.spi_buffer\[52\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
X_16967_ _09516_ _09477_ vssd1 vssd1 vccd1 vccd1 _09607_ sky130_fd_sc_hd__or2b_1
XFILLER_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18706_ _02400_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15918_ _08558_ _08562_ vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__or2b_1
X_19686_ _03069_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16898_ _09410_ _09412_ _09270_ _09409_ vssd1 vssd1 vccd1 vccd1 _09539_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18637_ _02275_ _02276_ _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15849_ _08047_ _08135_ _08491_ _08493_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__o22ai_4
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18568_ _02263_ _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17519_ _10051_ _10052_ _10084_ vssd1 vssd1 vccd1 vccd1 _10085_ sky130_fd_sc_hd__a21o_1
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18499_ _02184_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__xor2_1
X_20530_ _03421_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20461_ _03362_ _03363_ _03364_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__or3_1
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21013_ clknet_leaf_67_i_clk _00782_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11530_ _04244_ _04281_ _04289_ _04309_ _04140_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__a311o_1
XFILLER_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20728_ clknet_leaf_85_i_clk _00497_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ _04142_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__buf_4
X_20659_ clknet_leaf_25_i_clk _00443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13200_ _05930_ _05933_ _05936_ _05871_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a31o_1
X_10412_ _03537_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
X_14180_ _06914_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__nand2_1
X_11392_ rbzero.row_render.size\[6\] gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04172_
+ sky130_fd_sc_hd__or2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _05867_ _05697_ _05688_ _05783_ _05826_ _05801_ vssd1 vssd1 vccd1 vccd1 _05868_
+ sky130_fd_sc_hd__mux4_1
X_10343_ _03501_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13062_ _05794_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__nand2_1
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12013_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _04392_ vssd1 vssd1 vccd1 vccd1 _04788_
+ sky130_fd_sc_hd__mux2_1
X_17870_ _01471_ _01489_ _01487_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a21o_1
XFILLER_94_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16821_ _09461_ _09462_ vssd1 vssd1 vccd1 vccd1 _09463_ sky130_fd_sc_hd__or2_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19540_ _03002_ _03000_ _03011_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__or3_1
X_16752_ _09254_ _09255_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__or2_1
X_13964_ _06696_ _06690_ _06672_ _06698_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o22ai_1
XFILLER_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15703_ _08345_ _08346_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__03040_ clknet_0__03040_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03040_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12915_ _04031_ _05372_ _05651_ _04001_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a211o_1
X_16683_ _09186_ _09187_ _09325_ vssd1 vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19471_ rbzero.wall_tracer.rayAddendY\[4\] rbzero.wall_tracer.rayAddendY\[3\] _02904_
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__o21ai_2
XFILLER_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _06620_ _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__or2_1
XFILLER_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18422_ _02118_ _02119_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nand2_1
X_15634_ _08252_ _08261_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__nor2_1
XFILLER_179_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ rbzero.wall_tracer.visualWallDist\[-7\] _05351_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _02049_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__xor2_1
XFILLER_61_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _08208_ _08209_ _05194_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__o21ai_1
X_12777_ _05519_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _09864_ _09866_ _09865_ vssd1 vssd1 vccd1 vccd1 _09875_ sky130_fd_sc_hd__a21boi_1
XFILLER_14_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14516_ _07067_ _07069_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__nor2_1
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18284_ _01982_ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ rbzero.debug_overlay.playerY\[-7\] _04455_ _04501_ _04504_ _04506_ vssd1
+ vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a2111o_1
XFILLER_202_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15496_ _08097_ _08128_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__or2_1
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _09813_ sky130_fd_sc_hd__or2_1
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _07168_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__xnor2_1
X_11659_ _04424_ _04426_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17166_ rbzero.traced_texa\[-4\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__a22o_1
X_14378_ _06724_ _06740_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__or2_1
XFILLER_122_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _08739_ _08760_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13329_ _05752_ _06053_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
XFILLER_142_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17097_ _09735_ _09736_ vssd1 vssd1 vccd1 vccd1 _09737_ sky130_fd_sc_hd__nor2_2
XFILLER_116_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20252__271 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__inv_2
XFILLER_192_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16048_ _08654_ _08663_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__xnor2_2
XFILLER_142_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19628__80 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__inv_2
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19807_ _03132_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17999_ _09526_ _09480_ _09484_ _09391_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__o22a_1
Xclkbuf_1_1__f__03307_ clknet_0__03307_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03307_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19738_ rbzero.pov.spi_buffer\[43\] rbzero.pov.spi_buffer\[44\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
XFILLER_84_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19669_ rbzero.pov.spi_buffer\[10\] rbzero.pov.spi_buffer\[11\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
XFILLER_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21631_ clknet_leaf_37_i_clk _01400_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21562_ net483 _01331_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20513_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__and2b_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21493_ net414 _01262_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20335__346 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__inv_2
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20444_ rbzero.texV\[-7\] _03175_ _03332_ _03350_ vssd1 vssd1 vccd1 vccd1 _01389_
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20381__388 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__inv_2
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _03481_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__clkbuf_4
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20080__116 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__inv_2
XFILLER_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12700_ rbzero.wall_tracer.rayAddendX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__or2_1
XFILLER_204_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13680_ _06395_ _06415_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__or2_1
X_10892_ rbzero.tex_b1\[44\] rbzero.tex_b1\[45\] _03784_ vssd1 vssd1 vccd1 vccd1 _03792_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12631_ rbzero.map_rom.d6 _05377_ _05375_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15350_ _07990_ rbzero.wall_tracer.stepDistX\[-3\] _07994_ vssd1 vssd1 vccd1 vccd1
+ _07995_ sky130_fd_sc_hd__o21bai_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__nor2_1
XFILLER_197_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14301_ _07034_ _07036_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__and3_1
XFILLER_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11513_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _04291_ vssd1 vssd1 vccd1 vccd1 _04293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15281_ _05346_ _05468_ _07893_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ rbzero.wall_tracer.trackDistY\[-7\] _05238_ _05239_ rbzero.wall_tracer.trackDistY\[-8\]
+ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__o221a_1
X_17020_ _09539_ _09548_ _09547_ vssd1 vssd1 vccd1 vccd1 _09660_ sky130_fd_sc_hd__a21o_1
X_14232_ _06942_ _06943_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__or2_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11444_ _04138_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__buf_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14163_ _06893_ _06898_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__nor2_1
X_11375_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] rbzero.row_render.size\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__a21o_1
XFILLER_152_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ _05820_ _05849_ _05850_ _05798_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__o211a_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10326_ _03492_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
X_14094_ _06827_ _06829_ _06830_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__a21oi_1
X_18971_ _02615_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13045_ _05781_ _05702_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__or2_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _09103_ _09552_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__or2_1
XFILLER_65_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17853_ _10179_ _10181_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__or2_1
XFILLER_152_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16804_ _09309_ _09311_ vssd1 vssd1 vccd1 vccd1 _09446_ sky130_fd_sc_hd__and2_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17784_ _01485_ _01486_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__and2_1
XFILLER_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14996_ _07668_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19523_ _02979_ _02989_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__or2_1
X_13947_ _06673_ _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16735_ _09375_ _09376_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__nor2_1
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19454_ _02923_ _02925_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__or3_1
X_16666_ _09305_ _09306_ _09308_ vssd1 vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__nand3_1
XFILLER_207_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13878_ _06598_ _06599_ _06614_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__a21oi_4
XFILLER_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18405_ _01966_ _02000_ _02103_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a21oi_2
X_15617_ _08252_ _08261_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__xor2_2
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__buf_2
X_16597_ _09098_ _09108_ _09106_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__a21o_1
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19385_ _02870_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18336_ _01987_ _01994_ _02034_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a21o_1
X_15548_ _08179_ _08190_ _08192_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__a21o_1
XFILLER_124_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18267_ _08895_ _08767_ _01524_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__or3_1
X_15479_ _07951_ _08123_ _08062_ _05207_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__a211o_4
XFILLER_147_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _09792_ _09796_ _09797_ vssd1 vssd1 vccd1 vccd1 _09799_ sky130_fd_sc_hd__o21ai_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18198_ _01697_ _01780_ _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17149_ rbzero.row_render.texu\[0\] _09762_ _07728_ rbzero.wall_tracer.texu\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__a22o_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20160_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__buf_1
XFILLER_171_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ clknet_leaf_51_i_clk _00762_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21614_ clknet_leaf_43_i_clk _01383_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21545_ net466 _01314_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21476_ net397 _01245_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20427_ _03333_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_0__f__03043_ clknet_0__03043_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03043_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ rbzero.wall_tracer.mapX\[8\] _03947_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_
+ sky130_fd_sc_hd__or3b_1
XFILLER_175_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11091_ rbzero.tex_b0\[14\] rbzero.tex_b0\[13\] _03887_ vssd1 vssd1 vccd1 vccd1 _03896_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19607__61 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14850_ _07569_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__clkbuf_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _05824_ _06535_ _06536_ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__or4_1
X_19622__75 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14781_ _07487_ _07456_ _07513_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__a21oi_4
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11993_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _04250_ vssd1 vssd1 vccd1 vccd1 _04768_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16520_ _09163_ vssd1 vssd1 vccd1 vccd1 _09164_ sky130_fd_sc_hd__buf_2
XFILLER_84_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13732_ _06057_ _06045_ _05945_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__or3_1
XFILLER_147_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ _03819_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _08821_ _08059_ _09094_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__or3_1
X_13663_ _06357_ _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10875_ rbzero.tex_b1\[52\] rbzero.tex_b1\[53\] _03773_ vssd1 vssd1 vccd1 vccd1 _03783_
+ sky130_fd_sc_hd__mux2_1
X_15402_ _08046_ vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__buf_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ gpout0.vpos\[9\] _04315_ _02703_ _02706_ vssd1 vssd1 vccd1 vccd1 _02727_
+ sky130_fd_sc_hd__or4_1
X_12614_ _05315_ _05366_ _05314_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or3_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ rbzero.wall_tracer.visualWallDist\[6\] _08148_ vssd1 vssd1 vccd1 vccd1 _09027_
+ sky130_fd_sc_hd__nand2_4
X_13594_ _06302_ _06329_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__o21ba_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _01462_ _09480_ _09484_ _09526_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__o22a_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15333_ rbzero.wall_tracer.visualWallDist\[-9\] _07903_ vssd1 vssd1 vccd1 vccd1 _07978_
+ sky130_fd_sc_hd__or2_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12545_ _05297_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__and2_1
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20318__330 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__inv_2
XFILLER_177_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18052_ _10125_ _10136_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__nand2_1
XFILLER_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15264_ _07908_ rbzero.debug_overlay.playerY\[-6\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _07909_ sky130_fd_sc_hd__mux2_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12476_ _05214_ rbzero.wall_tracer.trackDistX\[10\] _05230_ vssd1 vssd1 vccd1 vccd1
+ _05231_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17003_ _07994_ _08705_ _08058_ _08150_ vssd1 vssd1 vccd1 vccd1 _09643_ sky130_fd_sc_hd__or4_1
X_14215_ _06852_ _06950_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__and2b_1
XANTENNA_5 _04374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _04143_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__buf_6
X_15195_ _07820_ _07730_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__and2_1
XFILLER_153_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _06842_ _06881_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__and2_1
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11358_ _04089_ _04114_ _04124_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__nor3b_2
XFILLER_125_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ rbzero.tex_r1\[63\] net46 _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux2_1
XFILLER_98_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14077_ _06800_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__xnor2_1
X_18954_ rbzero.pov.spi_buffer\[10\] rbzero.pov.ready_buffer\[10\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
X_11289_ _04065_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nor2_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _05567_ _05575_ _05656_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__o21a_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17905_ _01575_ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__xor2_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18885_ rbzero.spi_registers.new_vinf rbzero.spi_registers.spi_buffer\[0\] _02555_
+ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__mux2_1
XFILLER_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _10277_ _10279_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__or2b_1
XFILLER_187_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20364__372 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__inv_2
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17767_ _01461_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__xor2_1
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20063__100 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__inv_2
XFILLER_130_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14979_ _07659_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__clkbuf_1
X_19506_ _02963_ _02966_ _02964_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a21boi_1
X_16718_ _08162_ _09214_ _09359_ _09212_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__o31a_1
XFILLER_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17698_ _10258_ _10262_ vssd1 vssd1 vccd1 vccd1 _10263_ sky130_fd_sc_hd__xor2_2
XFILLER_74_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19437_ _02920_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__clkbuf_1
X_16649_ _09288_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__03037_ _03037_ vssd1 vssd1 vccd1 vccd1 clknet_0__03037_ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19368_ _07676_ _02856_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__nor2_1
XFILLER_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _01909_ _01911_ _01910_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__o21bai_1
XFILLER_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19299_ _02805_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21330_ net251 _01099_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21261_ clknet_leaf_62_i_clk _01030_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21192_ clknet_leaf_75_i_clk _00961_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ clknet_leaf_53_i_clk _00745_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _03670_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10591_ _03633_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12330_ net29 _05089_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__o21a_1
X_20192__217 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__inv_2
X_21528_ net449 _01297_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ net21 net22 _05027_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__and4_1
XFILLER_108_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21459_ net380 _01228_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[38\] sky130_fd_sc_hd__dfxtp_1
X_14000_ _06735_ _06736_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__nor2_1
X_11212_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__buf_2
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12192_ _04960_ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__nor2_1
XFILLER_162_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 o_gpout[0] sky130_fd_sc_hd__clkbuf_1
X_11143_ rbzero.debug_overlay.playerX\[2\] _03929_ rbzero.map_rom.d6 _03930_ _03931_
+ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a221o_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 o_rgb[23] sky130_fd_sc_hd__buf_2
XFILLER_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11074_ _03717_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15951_ _08591_ _08592_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__nand2_1
XFILLER_153_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14902_ _07591_ _07608_ _07609_ _04039_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__o211a_1
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15882_ _08476_ _08473_ vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__nand2_1
X_18670_ _08445_ _09704_ _02256_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__o31a_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _09912_ _10047_ _10045_ vssd1 vssd1 vccd1 vccd1 _10186_ sky130_fd_sc_hd__a21o_1
X_14833_ _07459_ _07439_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__nor2_1
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14764_ _07420_ _07347_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__nand2_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _10116_ _10117_ vssd1 vssd1 vccd1 vccd1 _10118_ sky130_fd_sc_hd__xnor2_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ rbzero.tex_b1\[30\] _04272_ _04265_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a21o_1
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13715_ _06441_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__or2_1
XFILLER_147_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16503_ _08976_ _08990_ _09146_ vssd1 vssd1 vccd1 vccd1 _09147_ sky130_fd_sc_hd__a21oi_2
X_10927_ _03810_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17483_ _09947_ _09949_ vssd1 vssd1 vccd1 vccd1 _10049_ sky130_fd_sc_hd__nor2_1
XFILLER_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14695_ _07418_ _07422_ _07424_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__or4b_1
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19222_ rbzero.color_floor\[5\] _02751_ _02760_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__a21o_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13646_ _06382_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__and3_1
X_16434_ _09077_ _09078_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__nand2_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10858_ _03774_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16365_ _07995_ _08109_ _08084_ _07931_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__o22a_1
X_19153_ rbzero.spi_registers.new_other\[9\] _02712_ vssd1 vssd1 vccd1 vccd1 _02717_
+ sky130_fd_sc_hd__or2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _06312_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__xnor2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ rbzero.tex_g0\[30\] rbzero.tex_g0\[29\] _03729_ vssd1 vssd1 vccd1 vccd1 _03738_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15316_ rbzero.wall_tracer.state\[3\] _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__nand2_1
X_18104_ _01700_ _01731_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__or2_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12528_ _05203_ _05211_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__o21ai_4
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16296_ _08719_ _08763_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__nor2_1
XFILLER_121_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19084_ _02674_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18035_ _08493_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__buf_2
X_15247_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__clkbuf_4
X_12459_ rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__inv_2
XFILLER_126_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15178_ _07816_ _07824_ _07828_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__a31o_1
XFILLER_114_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ _06769_ _06662_ _06667_ _06776_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__o22a_1
XFILLER_154_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19986_ _02721_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18937_ rbzero.pov.spi_buffer\[2\] rbzero.pov.ready_buffer\[2\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
XFILLER_97_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18868_ _02540_ _02541_ _02228_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17819_ _01516_ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__xor2_1
XFILLER_54_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18799_ _02479_ _02476_ _02480_ _02481_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a211o_1
XFILLER_48_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19601__56 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
X_20830_ clknet_leaf_1_i_clk _00599_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20761_ clknet_leaf_32_i_clk _00530_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20692_ clknet_leaf_7_i_clk _00476_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21313_ net234 _01082_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21244_ clknet_leaf_63_i_clk _01013_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_102_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21175_ clknet_leaf_74_i_clk _00944_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ rbzero.tex_g1\[59\] rbzero.tex_g1\[58\] _04337_ vssd1 vssd1 vccd1 vccd1 _04607_
+ sky130_fd_sc_hd__mux2_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04119_ _04526_ _04530_ _04538_ _04121_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__o311a_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ clknet_leaf_59_i_clk _00728_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13500_ _06160_ _06202_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nand2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _03697_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14480_ _07200_ _07215_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__nor2_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__buf_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20200__224 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__inv_2
XFILLER_202_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _06156_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__nor2_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10643_ _03661_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16150_ _08780_ _08781_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__nand2_1
X_13362_ _06025_ _06027_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10574_ rbzero.tex_r0\[4\] rbzero.tex_r0\[3\] _03624_ vssd1 vssd1 vccd1 vccd1 _03625_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15101_ _07741_ _07744_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__or2_1
X_12313_ net30 net31 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nor2_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16081_ _08723_ _08724_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__xnor2_1
X_13293_ _06024_ _06028_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__xor2_1
XFILLER_154_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15032_ rbzero.debug_overlay.vplaneX\[-9\] _03914_ _07679_ _07694_ _07696_ vssd1
+ vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a221o_1
XFILLER_182_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ net48 net39 net38 net40 net15 _04961_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__mux4_1
XFILLER_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19840_ _03139_ _03154_ _03156_ _03157_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__o211a_1
X_12175_ _04892_ _04909_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__o21a_1
XFILLER_150_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11126_ rbzero.wall_tracer.visualWallDist\[0\] rbzero.wall_tracer.visualWallDist\[-1\]
+ rbzero.wall_tracer.visualWallDist\[-2\] rbzero.wall_tracer.visualWallDist\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__or4_1
X_19771_ _03046_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__buf_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16983_ _08331_ _09621_ _09488_ _09622_ vssd1 vssd1 vccd1 vccd1 _09623_ sky130_fd_sc_hd__a31oi_1
XFILLER_89_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20407__8 clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
X_18722_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__or2_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _03878_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15934_ _08572_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__buf_2
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18653_ _02331_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__xnor2_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _08467_ _08464_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__and2b_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _09906_ _10168_ _10169_ vssd1 vssd1 vccd1 vccd1 _10170_ sky130_fd_sc_hd__o21a_1
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14816_ _07486_ _07399_ _07543_ _07527_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__a22o_1
XFILLER_97_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18584_ _02271_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _08391_ _08397_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__xnor2_1
Xtop_ew_algofoogle_110 vssd1 vssd1 vccd1 vccd1 ones[4] top_ew_algofoogle_110/LO sky130_fd_sc_hd__conb_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_121 vssd1 vssd1 vccd1 vccd1 ones[15] top_ew_algofoogle_121/LO sky130_fd_sc_hd__conb_1
XFILLER_92_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17535_ _09670_ _10099_ _10100_ vssd1 vssd1 vccd1 vccd1 _10101_ sky130_fd_sc_hd__a21o_1
X_11959_ _04206_ _04700_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__and3b_1
X_14747_ _07473_ _07478_ _07481_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__o21bai_1
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14678_ _07378_ _07413_ _07414_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__nor3_1
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17466_ _10032_ vssd1 vssd1 vccd1 vccd1 _10033_ sky130_fd_sc_hd__inv_2
XFILLER_177_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19205_ _09753_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__and2_1
X_13629_ _06355_ _06359_ _06365_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__o21ba_1
X_16417_ _08549_ _08957_ _09060_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__nand3_4
XFILLER_60_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17397_ _09126_ _08570_ vssd1 vssd1 vccd1 vccd1 _09964_ sky130_fd_sc_hd__nor2_1
X_20175__201 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__inv_2
XFILLER_125_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19136_ _04891_ _04887_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__nand3_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16348_ _08206_ _08248_ _08992_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__a21o_1
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19067_ rbzero.pov.spi_buffer\[64\] rbzero.pov.ready_buffer\[64\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
X_16279_ _08876_ _08923_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__nand2_1
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18018_ _01718_ _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19969_ rbzero.pov.ready_buffer\[42\] _03240_ _03243_ rbzero.debug_overlay.facingX\[0\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__o221a_1
XFILLER_80_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20813_ clknet_leaf_24_i_clk _00582_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20744_ clknet_leaf_35_i_clk _00513_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20675_ clknet_leaf_3_i_clk _00459_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[4\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0__f__03291_ clknet_0__03291_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03291_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21227_ clknet_leaf_73_i_clk _00996_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21158_ clknet_leaf_84_i_clk _00927_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13980_ _06245_ _06678_ _06715_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__o21bai_1
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21089_ net179 _00858_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12931_ _05628_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nand2_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15650_ _08289_ _08294_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__xnor2_1
X_12862_ _05594_ _05596_ _05598_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nor3_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _07327_ _07326_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__and2b_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _04205_ _04556_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__and3b_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ rbzero.wall_tracer.visualWallDist\[-11\] _04012_ vssd1 vssd1 vccd1 vccd1
+ _08226_ sky130_fd_sc_hd__nand2_2
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ rbzero.wall_tracer.mapY\[5\] _05397_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_
+ sky130_fd_sc_hd__o21a_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14532_ _07254_ _07257_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__nand2_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _05394_ vssd1 vssd1 vccd1 vccd1 _09889_ sky130_fd_sc_hd__clkbuf_4
X_11744_ _04522_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_8
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14463_ _07160_ _07199_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__nor2_1
X_17251_ _09824_ _09825_ _09827_ vssd1 vssd1 vccd1 vccd1 _09828_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11675_ _04433_ _04447_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and2_2
XFILLER_144_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13414_ _06021_ _06050_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__and2b_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16202_ _08840_ _08846_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__nand2_1
XFILLER_179_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17182_ rbzero.traced_texa\[9\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__a22o_1
X_10626_ _03652_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_1
X_14394_ _07111_ _07128_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__nand2_1
XFILLER_155_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16133_ _08660_ _08777_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__xnor2_1
X_13345_ _06063_ _06081_ _06073_ _06070_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a2bb2o_1
X_10557_ rbzero.tex_r0\[12\] rbzero.tex_r0\[11\] _03613_ vssd1 vssd1 vccd1 vccd1 _03616_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16064_ _08701_ _08708_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__xor2_1
X_13276_ _05978_ _05981_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__nor2_1
XFILLER_182_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ _03579_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15015_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__nor2_1
X_12227_ net49 _04962_ _04980_ net52 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a22o_1
XFILLER_97_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20170__197 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__inv_2
X_19823_ _03139_ _03142_ _03144_ _02765_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__o211a_1
XFILLER_190_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12158_ _04323_ _04903_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a21o_1
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11109_ _03905_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19754_ _03105_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12089_ _04858_ _04860_ net5 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__mux2_1
X_16966_ _09345_ _09590_ vssd1 vssd1 vccd1 vccd1 _09606_ sky130_fd_sc_hd__and2_1
X_18705_ rbzero.wall_tracer.trackDistY\[-12\] _02397_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02400_ sky130_fd_sc_hd__mux2_1
XFILLER_110_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15917_ _08482_ _08559_ _08560_ _08561_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__a2bb2o_1
X_19685_ rbzero.pov.spi_buffer\[18\] rbzero.pov.spi_buffer\[19\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
XFILLER_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16897_ _09518_ _09537_ vssd1 vssd1 vccd1 vccd1 _09538_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18636_ _02273_ _02274_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__and2_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _08129_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__buf_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18567_ _01498_ _09215_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15779_ _05208_ _08423_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__or2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17518_ _10069_ _10083_ vssd1 vssd1 vccd1 vccd1 _10084_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18498_ _02193_ _02195_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__xor2_1
XFILLER_127_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17449_ _09722_ _09724_ vssd1 vssd1 vccd1 vccd1 _10016_ sky130_fd_sc_hd__nor2_1
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20460_ _03357_ _03359_ _03358_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a21boi_1
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19119_ rbzero.spi_registers.spi_cmd\[2\] rbzero.spi_registers.spi_cmd\[3\] _02690_
+ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_106_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21012_ clknet_leaf_67_i_clk _00781_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20147__177 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__inv_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20727_ clknet_leaf_86_i_clk _00496_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _04237_ _04238_ _04239_ _04226_ _04210_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__o221a_1
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20658_ clknet_leaf_4_i_clk _00442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10411_ rbzero.tex_r1\[14\] rbzero.tex_r1\[15\] _03527_ vssd1 vssd1 vccd1 vccd1 _03537_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ rbzero.row_render.size\[6\] gpout0.hpos\[6\] _04004_ _04160_ _04170_ vssd1
+ vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__a221o_1
X_20589_ _03456_ _03457_ rbzero.wall_tracer.rayAddendX\[-6\] _09762_ vssd1 vssd1 vccd1
+ vccd1 _01427_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13130_ _05710_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__inv_2
XFILLER_87_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10342_ rbzero.tex_r1\[47\] rbzero.tex_r1\[48\] _03494_ vssd1 vssd1 vccd1 vccd1 _03501_
+ sky130_fd_sc_hd__mux2_1
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20312__325 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__inv_2
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13061_ _05754_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__nand2_2
XFILLER_139_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _04242_ _04778_ _04786_ _04207_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__o211a_1
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16820_ _09458_ _09460_ vssd1 vssd1 vccd1 vccd1 _09462_ sky130_fd_sc_hd__and2_1
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16751_ _09390_ _09392_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__and2_1
X_13963_ _06697_ _06699_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__nand2_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15702_ _08345_ _08346_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__xor2_1
XFILLER_189_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19470_ _02925_ _02935_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__nand2_1
X_12914_ rbzero.wall_tracer.visualWallDist\[6\] _04031_ vssd1 vssd1 vccd1 vccd1 _05651_
+ sky130_fd_sc_hd__nor2_1
X_13894_ _06629_ _06630_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__nand2_1
X_16682_ _09183_ _09185_ vssd1 vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__or2_1
XFILLER_47_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421_ _02118_ _02119_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__or2_1
XFILLER_59_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ _08268_ _08277_ vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__xnor2_2
X_12845_ _05561_ _05469_ _05580_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__o22a_2
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _10248_ _09977_ _01990_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__o31a_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _07560_ _07562_ _08171_ _07564_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__o31a_1
X_12776_ _05513_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__nand2_1
XFILLER_187_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17303_ _09872_ _09873_ vssd1 vssd1 vccd1 vccd1 _09874_ sky130_fd_sc_hd__or2b_1
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _07235_ _07251_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__xnor2_1
X_11727_ rbzero.debug_overlay.playerY\[3\] _04452_ _04464_ rbzero.debug_overlay.playerY\[-4\]
+ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a221o_1
X_15495_ _08109_ _08104_ _08042_ _08084_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__o22a_1
X_18283_ _09141_ _10238_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__nor2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17234_ _04016_ vssd1 vssd1 vccd1 vccd1 _09812_ sky130_fd_sc_hd__clkbuf_4
X_14446_ _07170_ _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__xor2_1
X_11658_ _04422_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__nor2_1
XFILLER_127_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ rbzero.tex_g1\[50\] rbzero.tex_g1\[51\] _03635_ vssd1 vssd1 vccd1 vccd1 _03643_
+ sky130_fd_sc_hd__mux2_1
X_14377_ _07112_ _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__nor2_1
X_17165_ rbzero.traced_texa\[-5\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__a22o_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ rbzero.tex_r1\[31\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__and3_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13328_ _05852_ _05853_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nand2_4
X_16116_ _08739_ _08760_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__xor2_2
XFILLER_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17096_ _09605_ _09606_ _09734_ vssd1 vssd1 vccd1 vccd1 _09736_ sky130_fd_sc_hd__o21a_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13259_ _05988_ _05989_ _05992_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a22o_1
X_16047_ _08682_ _08689_ _08691_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__a21oi_4
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20287__302 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__inv_2
XFILLER_69_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19806_ rbzero.pov.ss_buffer\[1\] rbzero.pov.ss_buffer\[0\] _05189_ vssd1 vssd1 vccd1
+ vccd1 _03132_ sky130_fd_sc_hd__mux2_1
XFILLER_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17998_ _01613_ _01631_ _01699_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19737_ _03096_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03306_ clknet_0__03306_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03306_
+ sky130_fd_sc_hd__clkbuf_16
X_16949_ _09587_ _09589_ vssd1 vssd1 vccd1 vccd1 _09590_ sky130_fd_sc_hd__xor2_1
X_20402__27 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19668_ _03060_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18619_ _02313_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__or2_1
X_21630_ clknet_leaf_36_i_clk _01399_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21561_ net482 _01330_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20512_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__nand2_1
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21492_ net413 _01261_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20443_ _03348_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_66_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10960_ _03827_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ _03791_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12630_ _05381_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__nor2_1
XFILLER_188_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__and2_1
XFILLER_196_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ _06911_ _06914_ _06884_ _06885_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__a211oi_2
X_11512_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _04291_ vssd1 vssd1 vccd1 vccd1 _04292_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15280_ _04013_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__buf_6
XFILLER_141_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12492_ _05239_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.trackDistY\[-9\]
+ _05240_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a221o_1
XFILLER_180_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _06888_ _06966_ _06963_ _06940_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__o211ai_1
XFILLER_138_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11443_ rbzero.tex_r0\[57\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_19_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14162_ _06893_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__nand2_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11374_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__clkbuf_4
XFILLER_153_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ _05797_ _05809_ _05839_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a21o_1
X_10325_ rbzero.tex_r1\[55\] rbzero.tex_r1\[56\] _03483_ vssd1 vssd1 vccd1 vccd1 _03492_
+ sky130_fd_sc_hd__mux2_1
X_14093_ _06804_ _06828_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__and2b_1
X_18970_ rbzero.pov.spi_buffer\[18\] rbzero.pov.ready_buffer\[18\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XFILLER_124_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13044_ _05695_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__clkinv_2
X_17921_ _01503_ _01623_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__xnor2_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ _01554_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__nand2_1
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _09405_ _09444_ vssd1 vssd1 vccd1 vccd1 _09445_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17783_ _01485_ _01486_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__nor2_1
XFILLER_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ rbzero.wall_tracer.stepDistX\[4\] _07566_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07668_ sky130_fd_sc_hd__mux2_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19522_ rbzero.wall_tracer.rayAddendY\[8\] _00013_ _02992_ _02999_ vssd1 vssd1 vccd1
+ vccd1 _00818_ sky130_fd_sc_hd__o22a_1
X_16734_ _09372_ _09374_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__and2_1
X_13946_ _06674_ _06679_ _06682_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20282__298 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__inv_2
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _02904_ rbzero.wall_tracer.rayAddendY\[4\] vssd1 vssd1 vccd1 vccd1 _02935_
+ sky130_fd_sc_hd__xor2_1
X_16665_ _09125_ _09148_ _09307_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__a21o_1
X_13877_ _06563_ _06600_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o21ai_2
XFILLER_179_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18404_ _01998_ _01999_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__nor2_1
X_15616_ _08256_ _08258_ _08260_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__a21boi_2
X_19384_ _02860_ _02863_ _02861_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a21bo_1
X_12828_ _04030_ _05327_ _05371_ _05564_ _04001_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a311o_1
X_16596_ _09209_ _09238_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18335_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__nor2_1
XFILLER_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _08170_ _08189_ _08191_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__o21ba_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12759_ _05504_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_175_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18266_ _01929_ _01965_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15478_ rbzero.wall_tracer.stepDistY\[-11\] vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__inv_2
XFILLER_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17217_ _09792_ _09796_ _09797_ vssd1 vssd1 vccd1 vccd1 _09798_ sky130_fd_sc_hd__or3_1
X_14429_ _06696_ _06663_ _06708_ _06698_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__o22a_1
XFILLER_190_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18197_ _01777_ _01779_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__nor2_1
XFILLER_129_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17148_ rbzero.row_render.size\[10\] _09762_ _07562_ _07756_ vssd1 vssd1 vccd1 vccd1
+ _00538_ sky130_fd_sc_hd__a22o_1
XFILLER_196_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17079_ _09571_ _09573_ vssd1 vssd1 vccd1 vccd1 _09719_ sky130_fd_sc_hd__and2b_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20992_ clknet_leaf_50_i_clk _00761_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20341__351 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__inv_2
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21613_ clknet_3_7_0_i_clk _01382_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21544_ net465 _01313_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20259__278 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__inv_2
XFILLER_194_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21475_ net396 _01244_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20426_ _03334_ _03335_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__and2b_1
XFILLER_135_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03042_ clknet_0__03042_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03042_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11090_ _03895_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _06529_ _06533_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__nor2_1
XFILLER_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14780_ _07459_ _07505_ _07510_ _07512_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__a31o_1
X_11992_ rbzero.tex_b1\[2\] _04272_ _04265_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a21o_1
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13731_ _06448_ _06450_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__xor2_1
X_10943_ rbzero.tex_b1\[20\] rbzero.tex_b1\[21\] _03817_ vssd1 vssd1 vccd1 vccd1 _03819_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16450_ _09092_ _09093_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__nand2_1
X_13662_ _06313_ _06356_ _06358_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__o21bai_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10874_ _03782_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15401_ _08045_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__buf_2
X_12613_ _05315_ _05366_ _05314_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__o21ai_1
X_13593_ _06303_ _06328_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _08369_ _08349_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__or2b_1
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _01735_ _01752_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12544_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or2_1
X_15332_ _05208_ rbzero.wall_tracer.stepDistX\[-2\] _07976_ vssd1 vssd1 vccd1 vccd1
+ _07977_ sky130_fd_sc_hd__a21boi_4
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18051_ _01735_ _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__xor2_1
XFILLER_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ _05212_ rbzero.wall_tracer.trackDistY\[11\] vssd1 vssd1 vccd1 vccd1 _05230_
+ sky130_fd_sc_hd__nor2_1
X_15263_ _07906_ _07907_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__and2_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03309_ clknet_0__03309_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03309_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17002_ _07994_ _08058_ _08151_ _08705_ vssd1 vssd1 vccd1 vccd1 _09642_ sky130_fd_sc_hd__o22a_1
X_14214_ _06950_ _06852_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__and2b_1
X_11426_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__buf_4
XANTENNA_6 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15194_ _07820_ _07730_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__nor2_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _06842_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__nor2_2
XFILLER_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11357_ _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14076_ _06802_ _06811_ _06812_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a21oi_1
X_18953_ _02606_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__clkbuf_1
X_11288_ rbzero.texV\[5\] _04066_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__a21boi_1
X_13027_ _05574_ _05662_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__xor2_2
X_17904_ _01591_ _01606_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__xnor2_1
X_18884_ rbzero.spi_registers.spi_done _03480_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_
+ sky130_fd_sc_hd__and3_1
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17835_ _01492_ _01538_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17766_ _01468_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nor2_1
XFILLER_82_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ rbzero.wall_tracer.stepDistX\[-4\] _07541_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07659_ sky130_fd_sc_hd__mux2_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19505_ _02982_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nand2_1
X_16717_ _09217_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__clkbuf_4
X_13929_ _05982_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__clkbuf_4
X_17697_ _10260_ _10261_ vssd1 vssd1 vccd1 vccd1 _10262_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19436_ rbzero.wall_tracer.rayAddendY\[2\] _02919_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _02920_ sky130_fd_sc_hd__mux2_1
X_16648_ _08239_ _09288_ _09289_ _09290_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__or4bb_1
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19367_ _02853_ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16579_ _09220_ _09221_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__and2_1
XFILLER_128_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__nand2_1
XFILLER_175_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19298_ rbzero.spi_registers.new_other\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__mux2_1
X_18249_ _01938_ _01948_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__nand2_1
XFILLER_175_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21260_ clknet_leaf_61_i_clk _01029_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21191_ clknet_leaf_75_i_clk _00960_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20975_ clknet_leaf_53_i_clk _00744_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10590_ rbzero.tex_g1\[59\] rbzero.tex_g1\[60\] _03549_ vssd1 vssd1 vccd1 vccd1 _03633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21527_ net448 _01296_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12260_ _05021_ net66 _05028_ net24 vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a211o_1
X_21458_ net379 _01227_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _03914_ _03999_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_1
X_20409_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__nand2_1
XFILLER_107_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12191_ net14 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__clkbuf_4
X_21389_ net310 _01158_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ rbzero.debug_overlay.playerY\[5\] rbzero.wall_tracer.mapY\[5\] vssd1 vssd1
+ vccd1 vccd1 _03931_ sky130_fd_sc_hd__xor2_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput54 net510 vssd1 vssd1 vccd1 vccd1 o_gpout[1] sky130_fd_sc_hd__clkbuf_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 o_rgb[6] sky130_fd_sc_hd__buf_2
XFILLER_150_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11073_ _03886_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15950_ _07974_ _08594_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__or2_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14901_ rbzero.wall_tracer.visualWallDist\[-7\] _07595_ vssd1 vssd1 vccd1 vccd1 _07609_
+ sky130_fd_sc_hd__or2_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _08517_ _08525_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__xor2_2
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _10169_ _10166_ _10165_ vssd1 vssd1 vccd1 vccd1 _10185_ sky130_fd_sc_hd__a21oi_2
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _00004_ _07555_ _07556_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a21oi_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _09114_ _09552_ vssd1 vssd1 vccd1 vccd1 _10117_ sky130_fd_sc_hd__nor2_1
X_14763_ _07419_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__clkinv_2
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ rbzero.tex_b1\[31\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__and3_1
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _08989_ _08987_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__and2b_1
X_13714_ _06442_ _06447_ _06448_ _06450_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_204_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10926_ rbzero.tex_b1\[28\] rbzero.tex_b1\[29\] _03806_ vssd1 vssd1 vccd1 vccd1 _03810_
+ sky130_fd_sc_hd__mux2_1
X_17482_ _09912_ _10047_ vssd1 vssd1 vccd1 vccd1 _10048_ sky130_fd_sc_hd__xor2_1
XFILLER_189_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14694_ _05742_ _07426_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__a21o_1
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19221_ rbzero.spi_registers.new_floor\[5\] rbzero.spi_registers.got_new_floor _02711_
+ _03911_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a31o_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16433_ _09074_ _09075_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__or2_1
XFILLER_72_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13645_ _06065_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__inv_2
X_10857_ rbzero.tex_b1\[61\] rbzero.tex_b1\[62\] _03773_ vssd1 vssd1 vccd1 vccd1 _03774_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19152_ rbzero.otherx\[2\] _02710_ _02716_ _02714_ vssd1 vssd1 vccd1 vccd1 _00731_
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ _07995_ _08570_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__nor2_1
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13576_ _05946_ _05939_ _06007_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__or3_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _03737_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _01563_ _01565_ _01696_ _01694_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a31o_1
X_15315_ _05360_ _05472_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__mux2_1
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19083_ rbzero.pov.spi_buffer\[72\] rbzero.pov.ready_buffer\[72\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
X_12527_ _04017_ _05279_ _05281_ _03970_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o211a_1
XFILLER_158_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16295_ _08851_ _08936_ _08937_ _08939_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__o211a_1
X_18034_ _01634_ _01642_ _01641_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a21bo_1
XFILLER_145_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15246_ _07892_ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12458_ _05212_ rbzero.wall_tracer.trackDistY\[11\] vssd1 vssd1 vccd1 vccd1 _05213_
+ sky130_fd_sc_hd__and2_1
XFILLER_193_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11409_ _04150_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__nand2_1
X_12389_ net38 _05142_ _05139_ net48 _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a221o_1
XFILLER_125_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15177_ _07830_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__buf_6
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ _06805_ _06707_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__or2_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19985_ rbzero.pov.ready_buffer\[12\] _03252_ _03253_ rbzero.debug_overlay.vplaneX\[-8\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__o221a_1
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14059_ _06786_ _06794_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18936_ _02597_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18867_ _02537_ _02538_ _02539_ _04016_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a31o_1
X_19598__53 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17818_ _01517_ _01521_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__xor2_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18798_ _05257_ _08200_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__nor2_1
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17749_ _01451_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__nor2_1
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20760_ clknet_leaf_32_i_clk _00529_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19419_ _07756_ _02896_ _02897_ _02903_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__a31o_1
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20691_ clknet_leaf_26_i_clk _00475_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21312_ net233 _01081_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21243_ clknet_leaf_63_i_clk _01012_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21174_ clknet_leaf_79_i_clk _00943_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11760_ _04208_ _04533_ _04537_ _04142_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a211o_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ clknet_leaf_52_i_clk _00727_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ rbzero.tex_g1\[2\] rbzero.tex_g1\[3\] _03691_ vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11691_ rbzero.debug_overlay.vplaneX\[10\] _04453_ _04457_ _04469_ vssd1 vssd1 vccd1
+ vccd1 _04470_ sky130_fd_sc_hd__a211o_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20889_ clknet_leaf_83_i_clk _00658_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13430_ _06157_ _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10642_ rbzero.tex_g1\[35\] rbzero.tex_g1\[36\] _03658_ vssd1 vssd1 vccd1 vccd1 _03661_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ _06094_ _06095_ _06096_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a21o_1
XFILLER_210_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _03557_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__buf_4
XFILLER_107_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15100_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__or2_1
X_12312_ _05031_ _05041_ _05079_ _05080_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__o31a_2
XFILLER_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13292_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__inv_2
XFILLER_154_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16080_ _08723_ _08724_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__nand2_1
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12243_ net46 _04980_ _05012_ _05010_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15031_ rbzero.wall_tracer.rayAddendX\[-5\] _07695_ vssd1 vssd1 vccd1 vccd1 _07696_
+ sky130_fd_sc_hd__and2_1
XFILLER_170_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12174_ gpout0.vpos\[0\] net8 net10 net9 vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__o211a_1
XFILLER_150_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11125_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__buf_4
X_19770_ _03113_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16982_ _08329_ _09216_ _09351_ _08054_ vssd1 vssd1 vccd1 vccd1 _09622_ sky130_fd_sc_hd__o22a_1
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18721_ _02413_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _03876_ vssd1 vssd1 vccd1 vccd1 _03878_
+ sky130_fd_sc_hd__mux2_1
X_15933_ _08569_ _08577_ vssd1 vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18652_ _02342_ _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _08487_ _08506_ _08508_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__a21oi_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17603_ _10023_ _10025_ vssd1 vssd1 vccd1 vccd1 _10169_ sky130_fd_sc_hd__or2_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _05894_ _07413_ _07516_ _07473_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__a22o_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18583_ _02278_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__and2b_1
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_100 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_100/HI zeros[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_184_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15795_ _08400_ _08409_ vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__xnor2_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_111 vssd1 vssd1 vccd1 vccd1 ones[5] top_ew_algofoogle_111/LO sky130_fd_sc_hd__conb_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _09276_ _08570_ _09417_ _08111_ vssd1 vssd1 vccd1 vccd1 _10100_ sky130_fd_sc_hd__o22a_1
X_14746_ _05844_ _07477_ _07479_ _07480_ _05800_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__a311o_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11958_ _04207_ _04708_ _04716_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a31o_1
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10909_ rbzero.tex_b1\[36\] rbzero.tex_b1\[37\] _03795_ vssd1 vssd1 vccd1 vccd1 _03801_
+ sky130_fd_sc_hd__mux2_1
X_17465_ _10029_ _09902_ _10030_ _10031_ vssd1 vssd1 vccd1 vccd1 _10032_ sky130_fd_sc_hd__a211o_1
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14677_ _07407_ _07409_ _07412_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__and3b_1
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11889_ _04663_ _04665_ _04521_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a21bo_4
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19204_ rbzero.spi_registers.new_sky\[5\] rbzero.color_sky\[5\] _02740_ vssd1 vssd1
+ vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
XFILLER_189_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16416_ _08549_ _08957_ _09060_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__a21o_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ _06360_ _06363_ _06364_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__and3_1
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17396_ _09961_ _09962_ vssd1 vssd1 vccd1 vccd1 _09963_ sky130_fd_sc_hd__and2_1
XFILLER_158_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19135_ _02702_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__clkbuf_1
X_16347_ _08241_ _08247_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__nor2_1
X_13559_ _06294_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19066_ _02665_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16278_ _08867_ _08875_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__or2_1
X_18017_ _08259_ _08157_ _08149_ _08188_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__o22ai_1
X_15229_ _07821_ _04033_ _07878_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__or3_1
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19968_ rbzero.pov.ready_buffer\[41\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-1\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__a221o_1
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18919_ _02585_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19899_ _07908_ _03141_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__nor2_1
XFILLER_110_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20812_ clknet_leaf_29_i_clk _00581_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20743_ clknet_leaf_35_i_clk _00512_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20674_ clknet_leaf_3_i_clk _00458_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03290_ clknet_0__03290_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03290_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21226_ clknet_leaf_73_i_clk _00995_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_160_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21157_ clknet_leaf_84_i_clk _00926_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21088_ net178 _00857_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20039_ _02741_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__nor2_1
X_12930_ _05652_ _05659_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nand2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19577__34 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _05481_ _05597_ _05561_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__mux2_2
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _07107_ _07335_ _07336_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__or3b_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04207_ _04564_ _04572_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a31o_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _08219_ _08221_ _08224_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__a21oi_2
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ rbzero.wall_tracer.mapY\[5\] _05397_ _05406_ vssd1 vssd1 vccd1 vccd1 _05535_
+ sky130_fd_sc_hd__a21o_1
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14531_ _07252_ _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__xnor2_1
X_19592__48 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
X_20124__156 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__inv_2
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _04411_ _04413_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__o21a_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17250_ _08944_ _08948_ _09826_ vssd1 vssd1 vccd1 vccd1 _09827_ sky130_fd_sc_hd__a21o_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _07162_ _07194_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__o21a_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11674_ _04445_ _04449_ _04451_ _04452_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__or4_4
XFILLER_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16201_ _08812_ _08844_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__xor2_1
X_13413_ _06145_ _06149_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__nor2_1
XFILLER_174_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17181_ rbzero.traced_texa\[8\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__a22o_1
X_10625_ rbzero.tex_g1\[43\] rbzero.tex_g1\[44\] _03647_ vssd1 vssd1 vccd1 vccd1 _03652_
+ sky130_fd_sc_hd__mux2_1
X_14393_ _06689_ _07072_ _07110_ _07108_ _06675_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__o32ai_1
X_16132_ _08767_ _08579_ _08727_ _08776_ _08774_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__o41a_1
X_13344_ _06078_ _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__or2_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10556_ _03615_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16063_ _08704_ _08706_ _08707_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__a21oi_1
X_10487_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _03569_ vssd1 vssd1 vccd1 vccd1 _03579_
+ sky130_fd_sc_hd__mux2_1
X_13275_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__inv_2
XFILLER_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15014_ _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__buf_4
X_12226_ _04977_ net16 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nand2_2
XFILLER_155_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12157_ _04907_ _04910_ net68 _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a31o_1
XFILLER_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19822_ _03140_ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__nand2_1
XFILLER_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ rbzero.tex_b0\[6\] rbzero.tex_b0\[5\] _03898_ vssd1 vssd1 vccd1 vccd1 _03905_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12088_ net40 _04855_ _04853_ net39 _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a221o_1
X_16965_ _09587_ _09589_ vssd1 vssd1 vccd1 vccd1 _09605_ sky130_fd_sc_hd__nor2_1
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19753_ rbzero.pov.spi_buffer\[50\] rbzero.pov.spi_buffer\[51\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03105_ sky130_fd_sc_hd__mux2_1
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11039_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _03865_ vssd1 vssd1 vccd1 vccd1 _03869_
+ sky130_fd_sc_hd__mux2_1
X_15916_ _08482_ _08559_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__xor2_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _02398_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__buf_4
X_19684_ _03068_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__clkbuf_1
X_16896_ _09520_ _09536_ vssd1 vssd1 vccd1 vccd1 _09537_ sky130_fd_sc_hd__xor2_1
XFILLER_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18635_ _09429_ _09433_ _08356_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a21o_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _08129_ _08047_ _08135_ _08491_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__or4_4
XFILLER_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18566_ _02261_ _02262_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__and2_1
XFILLER_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ rbzero.wall_tracer.visualWallDist\[5\] _04014_ vssd1 vssd1 vccd1 vccd1 _08423_
+ sky130_fd_sc_hd__nand2_4
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17517_ _10080_ _10082_ vssd1 vssd1 vccd1 vccd1 _10083_ sky130_fd_sc_hd__xor2_1
XFILLER_166_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14729_ _07456_ _07464_ _07459_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__mux2_2
XFILLER_162_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18497_ _02084_ _02092_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20099__133 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__inv_2
XFILLER_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ _09955_ _10014_ vssd1 vssd1 vccd1 vccd1 _10015_ sky130_fd_sc_hd__xnor2_2
XFILLER_178_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17379_ _09940_ _09945_ vssd1 vssd1 vccd1 vccd1 _09946_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19118_ _02693_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19049_ _02656_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21011_ clknet_leaf_67_i_clk _00780_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20726_ clknet_leaf_87_i_clk _00495_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20657_ clknet_leaf_0_i_clk _00441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10410_ _03536_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _04160_ gpout0.hpos\[5\] _04022_ _04161_ _04169_ vssd1 vssd1 vccd1 vccd1
+ _04170_ sky130_fd_sc_hd__o221a_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20588_ _07683_ _07692_ _07691_ _07831_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a31o_1
XFILLER_165_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10341_ _03500_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13060_ _05795_ _05796_ _05743_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a21o_1
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12011_ _04210_ _04781_ _04785_ _04371_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a211o_1
X_21209_ clknet_leaf_17_i_clk _00978_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_132_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16750_ _09391_ _08356_ _09389_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__o21ai_1
X_13962_ _06698_ _06690_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__nor2_1
XFILLER_150_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15701_ _08076_ _08085_ _08106_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__o21ba_1
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12913_ _05601_ _05606_ _05638_ _05649_ _05628_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__o41a_2
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16681_ _09321_ _09323_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__xnor2_1
X_13893_ _06579_ _06628_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__nand2_1
X_18420_ _01807_ _01810_ _01927_ _01925_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a31oi_4
XFILLER_59_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _08276_ _08008_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__nor2_1
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12844_ rbzero.wall_tracer.visualWallDist\[-5\] _05570_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05581_ sky130_fd_sc_hd__a21o_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18351_ _01988_ _01989_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__nand2_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _07560_ _07562_ _07564_ _08171_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__nor4_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _05511_ _05515_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or2_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09873_ sky130_fd_sc_hd__nand2_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14514_ _07245_ _07244_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__and2b_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18282_ _01737_ _09693_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__nor2_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ rbzero.debug_overlay.playerY\[5\] _04444_ _04439_ _04465_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__a32o_1
X_15494_ _08109_ _08042_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__or2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17233_ _05243_ _09781_ _09811_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14445_ _07175_ _07180_ _07181_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__o21a_1
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11657_ _04415_ _04430_ _04417_ _04022_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or4b_2
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17164_ rbzero.traced_texa\[-6\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a22o_1
XFILLER_70_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10608_ _03642_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ _06689_ _06760_ _07110_ _07108_ _06675_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__o32a_1
X_11588_ rbzero.tex_r1\[29\] rbzero.tex_r1\[28\] _04342_ vssd1 vssd1 vccd1 vccd1 _04367_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16115_ _08756_ _08758_ _08759_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__a21oi_2
X_13327_ _06058_ _06062_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__xnor2_1
X_10539_ _03606_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17095_ _09605_ _09606_ _09734_ vssd1 vssd1 vccd1 vccd1 _09735_ sky130_fd_sc_hd__nor3_1
XFILLER_182_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16046_ _08662_ _08690_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__nand2_1
X_13258_ _05994_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__buf_2
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12209_ _04323_ _04962_ _04978_ net68 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a22o_1
XFILLER_124_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13189_ _05807_ _05858_ _05871_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19805_ _03131_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17997_ _01615_ _01630_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nor2_1
X_20399__24 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
XFILLER_78_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03305_ clknet_0__03305_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03305_
+ sky130_fd_sc_hd__clkbuf_16
X_19736_ rbzero.pov.spi_buffer\[42\] rbzero.pov.spi_buffer\[43\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03096_ sky130_fd_sc_hd__mux2_1
X_16948_ _09347_ _09450_ _09588_ vssd1 vssd1 vccd1 vccd1 _09589_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19667_ rbzero.pov.spi_buffer\[9\] rbzero.pov.spi_buffer\[10\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
X_16879_ _09407_ _09414_ _09519_ vssd1 vssd1 vccd1 vccd1 _09520_ sky130_fd_sc_hd__a21o_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18618_ _02312_ _02314_ _05204_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a21o_1
XFILLER_198_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20107__140 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__inv_2
X_18549_ _02241_ _02245_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__xor2_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21560_ net481 _01329_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20511_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03407_
+ sky130_fd_sc_hd__nor2_1
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21491_ net412 _01260_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20442_ _03343_ _03345_ _03344_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o21bai_1
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20153__182 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__inv_2
XFILLER_115_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10890_ rbzero.tex_b1\[45\] rbzero.tex_b1\[46\] _03784_ vssd1 vssd1 vccd1 vccd1 _03791_
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12560_ _05313_ _05287_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__nor2_1
XFILLER_93_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11511_ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20709_ clknet_leaf_12_i_clk _00000_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12491_ rbzero.wall_tracer.trackDistY\[-9\] _05240_ rbzero.wall_tracer.trackDistY\[-10\]
+ _05241_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__o221a_1
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14230_ _06888_ _06966_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nand2_1
XFILLER_184_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ _04136_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__buf_4
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20236__257 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__inv_2
X_14161_ _06894_ _06896_ _06897_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__a21oi_1
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ rbzero.row_render.size\[7\] _04152_ rbzero.row_render.size\[8\] vssd1 vssd1
+ vccd1 vccd1 _04153_ sky130_fd_sc_hd__o21a_1
XFILLER_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10324_ _03491_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
X_13112_ _05718_ _05734_ _05803_ _05721_ _05777_ _05801_ vssd1 vssd1 vccd1 vccd1 _05849_
+ sky130_fd_sc_hd__mux4_1
XFILLER_180_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ _06804_ _06828_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13043_ _05695_ _05702_ _05677_ _05762_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__or4_1
XFILLER_140_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17920_ _08802_ _09693_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__nor2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17851_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__or2_1
XFILLER_121_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16802_ _09442_ _09443_ vssd1 vssd1 vccd1 vccd1 _09444_ sky130_fd_sc_hd__xor2_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17782_ _10215_ _10224_ _10222_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a21oi_1
X_14994_ _07667_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19521_ _03913_ _02997_ _02998_ _07695_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a31o_1
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16733_ _09372_ _09374_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__nor2_1
X_13945_ _06675_ _06668_ _06681_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__o21ba_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19452_ _07831_ _02925_ _02926_ _02934_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__o31ai_1
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16664_ _09145_ _09147_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__nor2_1
X_13876_ _06560_ _06601_ _06603_ _06612_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__a211oi_2
XFILLER_90_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18403_ _02060_ _02101_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__xnor2_1
X_15615_ _08259_ _08226_ _08244_ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__or3_1
XFILLER_37_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19383_ _02868_ _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_1
X_12827_ _03953_ _04030_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__nor2_1
XFILLER_188_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16595_ _09210_ _09237_ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _02031_ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nor2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15546_ _08177_ _07989_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__nor2_1
XFILLER_203_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12758_ rbzero.map_rom.f2 _05496_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__nor2_1
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18265_ _01932_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__xor2_1
X_11709_ rbzero.debug_overlay.facingY\[10\] _04453_ _04487_ vssd1 vssd1 vccd1 vccd1
+ _04488_ sky130_fd_sc_hd__a21oi_1
X_15477_ _08120_ _08121_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__nand2_1
X_12689_ _05420_ _05431_ _05419_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a21o_1
XFILLER_204_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17216_ rbzero.wall_tracer.mapX\[10\] _05525_ vssd1 vssd1 vccd1 vccd1 _09797_ sky130_fd_sc_hd__xor2_1
X_14428_ _06067_ _06668_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__or2_1
XFILLER_175_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18196_ _01817_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ rbzero.row_render.size\[9\] _09762_ _07560_ _07756_ vssd1 vssd1 vccd1 vccd1
+ _00537_ sky130_fd_sc_hd__a22o_1
X_14359_ _07031_ _07033_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nor2_1
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _09692_ _09717_ vssd1 vssd1 vccd1 vccd1 _09718_ sky130_fd_sc_hd__xnor2_2
XFILLER_118_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16029_ _08019_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19719_ rbzero.pov.spi_buffer\[34\] rbzero.pov.spi_buffer\[35\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
X_20991_ clknet_leaf_38_i_clk _00760_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03319_ _03319_ vssd1 vssd1 vccd1 vccd1 clknet_0__03319_ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21612_ net129 _01381_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21543_ net464 _01312_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21474_ net395 _01243_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20425_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0__f__03041_ clknet_0__03041_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03041_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ rbzero.tex_b1\[3\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and3_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13730_ _06440_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__xor2_1
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10942_ _03818_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13661_ _06365_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__or2_1
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ rbzero.tex_b1\[53\] rbzero.tex_b1\[54\] _03773_ vssd1 vssd1 vccd1 vccd1 _03782_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15400_ _07945_ _08044_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__or2_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _05308_ _05312_ _05318_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__o21a_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _09022_ _09024_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__xor2_2
X_13592_ _06303_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__xnor2_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15331_ _07925_ _07974_ _07975_ _05207_ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__a211o_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__nand2_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18050_ _01736_ _01751_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__xnor2_1
X_15262_ rbzero.debug_overlay.playerY\[-6\] _07905_ vssd1 vssd1 vccd1 vccd1 _07907_
+ sky130_fd_sc_hd__nand2_1
XFILLER_185_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _05219_ _05227_ _05228_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__o21a_1
XFILLER_126_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03308_ clknet_0__03308_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03308_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17001_ _09245_ _08159_ vssd1 vssd1 vccd1 vccd1 _09641_ sky130_fd_sc_hd__nor2_1
X_14213_ _06666_ _06690_ _06921_ _06919_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__o31a_1
X_11425_ rbzero.floor_leak\[5\] _04116_ _04133_ _04134_ _04204_ vssd1 vssd1 vccd1
+ vccd1 _04205_ sky130_fd_sc_hd__a221o_1
X_15193_ _07843_ _07844_ _07841_ _07842_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__a211o_1
XANTENNA_7 _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14144_ _06856_ _06879_ _06880_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__a21oi_2
X_11356_ _04127_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10307_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__buf_4
XFILLER_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14075_ _06803_ _06810_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nor2_1
X_18952_ rbzero.pov.spi_buffer\[9\] rbzero.pov.ready_buffer\[9\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
X_11287_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _04067_ sky130_fd_sc_hd__nand2_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13026_ _05761_ _05762_ _05748_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and3_1
X_17903_ _01604_ _01605_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__nor2_1
X_18883_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\]
+ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__and4bb_1
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17834_ _01535_ _01537_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__xor2_1
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14977_ _00008_ _07536_ _07658_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17765_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__and2_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19504_ rbzero.debug_overlay.vplaneY\[-1\] _02961_ vssd1 vssd1 vccd1 vccd1 _02983_
+ sky130_fd_sc_hd__nand2_1
X_13928_ _06659_ _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nand2_1
X_16716_ _09356_ _09357_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__xnor2_1
X_17696_ _10110_ _09973_ vssd1 vssd1 vccd1 vccd1 _10261_ sky130_fd_sc_hd__nor2_1
XFILLER_90_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19435_ _02908_ _02909_ _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__o21ai_1
X_16647_ _08215_ _08519_ _08985_ _09138_ vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__or4_1
X_13859_ _06564_ _06594_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__or2_1
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19366_ _02854_ _02842_ _02841_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a21oi_2
X_16578_ _09161_ _09219_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__or2_1
XFILLER_50_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18317_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__or2_1
X_15529_ _07894_ _05342_ _08173_ _07970_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__o211a_1
X_19297_ _02804_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _01946_ _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__and2_1
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20219__241 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__inv_2
XFILLER_204_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18179_ _10110_ _10266_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__nor2_1
XFILLER_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21190_ clknet_leaf_77_i_clk _00959_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20072_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__buf_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20265__283 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__inv_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20974_ clknet_leaf_53_i_clk _00743_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21526_ net447 _01295_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21457_ net378 _01226_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ _03970_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__and2_1
X_20408_ gpout5.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__nor2_1
X_12190_ net15 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21388_ net309 _01157_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ rbzero.debug_overlay.playerY\[0\] vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__inv_2
XFILLER_134_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 o_gpout[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 o_rgb[7] sky130_fd_sc_hd__buf_2
X_11072_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _03876_ vssd1 vssd1 vccd1 vccd1 _03886_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14900_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.trackDistX\[-7\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20348__358 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__inv_2
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15880_ _08522_ _08523_ _08524_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__o21ba_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ rbzero.wall_tracer.stepDistY\[0\] _07461_ vssd1 vssd1 vccd1 vccd1 _07556_
+ sky130_fd_sc_hd__nor2_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _09980_ _10115_ vssd1 vssd1 vccd1 vccd1 _10116_ sky130_fd_sc_hd__xnor2_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _05884_ _07492_ _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__a21o_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _04342_ vssd1 vssd1 vccd1 vccd1 _04749_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16501_ _09132_ _09144_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__xnor2_2
XFILLER_189_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13713_ _06041_ _06449_ _06407_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__mux2_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _03809_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__clkbuf_1
X_17481_ _10045_ _10046_ vssd1 vssd1 vccd1 vccd1 _10047_ sky130_fd_sc_hd__nor2_1
X_14693_ _05779_ _07428_ _07429_ _05892_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__o211a_1
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16432_ _09074_ _09075_ _09076_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__a21o_1
X_19220_ _02759_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13644_ _05988_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__xnor2_1
X_10856_ _03646_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__clkbuf_4
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ rbzero.spi_registers.new_other\[8\] _02712_ vssd1 vssd1 vccd1 vccd1 _02716_
+ sky130_fd_sc_hd__or2_1
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _09006_ _09007_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__and2_1
X_13575_ _05823_ _05961_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__or2_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _03729_ vssd1 vssd1 vccd1 vccd1 _03737_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18102_ _01784_ _01686_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__or2b_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ _07958_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__buf_4
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ _02673_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
X_12526_ _03912_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nor2_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16294_ _08803_ _08804_ _08807_ _08938_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__a211oi_1
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20093__128 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__inv_2
X_18033_ _01622_ _01629_ _01734_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a21o_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _04035_ _07891_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__and2_1
X_12457_ rbzero.wall_tracer.trackDistX\[11\] vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__inv_2
XFILLER_67_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ rbzero.row_render.size\[3\] _04149_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__nand2_1
X_15176_ _04033_ _04027_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__nand2_4
X_12388_ net40 _05145_ _05143_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__and3_1
XFILLER_126_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _06769_ _06667_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__nor2_1
XFILLER_181_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11339_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__clkbuf_4
XFILLER_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19984_ rbzero.pov.ready_buffer\[11\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-9\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__a221o_1
XFILLER_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ _06789_ _06793_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__or2b_1
X_18935_ rbzero.pov.spi_buffer\[1\] rbzero.pov.ready_buffer\[1\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13009_ _05690_ _05702_ _05683_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__or4_1
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18866_ _02537_ _02538_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17817_ _01519_ _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18797_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__nor2_1
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17748_ _01443_ _01444_ _01450_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__and3_1
XFILLER_78_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17679_ _08802_ _09552_ vssd1 vssd1 vccd1 vccd1 _10244_ sky130_fd_sc_hd__nor2_1
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19418_ rbzero.wall_tracer.rayAddendY\[1\] _07695_ _02902_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _02903_ sky130_fd_sc_hd__a22o_1
XFILLER_165_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20690_ clknet_leaf_26_i_clk _00474_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19349_ _07728_ _02838_ _02839_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a21o_1
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21311_ net232 _01080_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21242_ clknet_leaf_80_i_clk _01011_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21173_ clknet_leaf_79_i_clk _00942_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ clknet_leaf_41_i_clk _00726_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _03696_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__clkbuf_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11690_ rbzero.debug_overlay.vplaneX\[-9\] _04458_ _04461_ _04468_ vssd1 vssd1 vccd1
+ vccd1 _04469_ sky130_fd_sc_hd__a211o_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ clknet_leaf_82_i_clk _00657_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _03660_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13360_ _06094_ _06095_ _06096_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__nand3_1
X_10572_ _03623_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12311_ net24 net25 net66 _05068_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__or4_1
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21509_ net430 _01278_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _05855_ _06010_ _06025_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a22o_1
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ _04028_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__buf_4
X_12242_ _04867_ _04964_ net47 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12173_ _04154_ _03477_ net8 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__mux2_1
XFILLER_135_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__buf_4
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16981_ _05211_ _09350_ vssd1 vssd1 vccd1 vccd1 _09621_ sky130_fd_sc_hd__nor2_1
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18720_ rbzero.wall_tracer.trackDistY\[-10\] _02412_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _03877_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__clkbuf_1
X_15932_ _08570_ _08128_ _08571_ _08576_ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__o31a_1
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15863_ _08154_ _08507_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__nand2_1
X_18651_ _02345_ _02346_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14814_ _07542_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__clkbuf_1
X_17602_ _10023_ _10025_ vssd1 vssd1 vccd1 vccd1 _10168_ sky130_fd_sc_hd__and2_1
XFILLER_91_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _08412_ _08438_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__xnor2_1
X_18582_ _02272_ _02277_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__or2_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_101 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_101/HI zeros[11]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_112 vssd1 vssd1 vccd1 vccd1 ones[6] top_ew_algofoogle_112/LO sky130_fd_sc_hd__conb_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _07384_ _07401_ _05844_ _05952_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__o211a_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _09668_ _09417_ vssd1 vssd1 vccd1 vccd1 _10099_ sky130_fd_sc_hd__nor2_1
X_11957_ _04244_ _04724_ _04732_ _04116_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a31o_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10908_ _03800_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17464_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _10031_ sky130_fd_sc_hd__and2_1
X_14676_ _07407_ _07410_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__o21ba_2
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ _04206_ _04664_ _04314_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a21oi_1
XFILLER_189_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16415_ _09059_ _08547_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__xnor2_2
X_19203_ rbzero.color_sky\[4\] _02740_ _02748_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__a21o_1
X_13627_ _06078_ _05982_ _06361_ _06362_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__o211ai_1
XFILLER_60_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10839_ _03764_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
X_17395_ _09661_ _08356_ _09960_ vssd1 vssd1 vccd1 vccd1 _09962_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20101__135 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__inv_2
XFILLER_73_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19134_ rbzero.spi_registers.sclk_buffer\[1\] rbzero.spi_registers.sclk_buffer\[2\]
+ _02695_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
X_16346_ _08976_ _08990_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__xnor2_2
XFILLER_186_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13558_ _05888_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__and3_1
XFILLER_185_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ rbzero.wall_tracer.trackDistX\[3\] vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__inv_2
X_19065_ rbzero.pov.spi_buffer\[63\] rbzero.pov.ready_buffer\[63\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
X_16277_ _08912_ _08913_ _08920_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__and4b_1
X_13489_ _06197_ _06198_ _06224_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or3_1
XFILLER_121_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15228_ _07730_ _07854_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__nor2_1
X_18016_ _08259_ _08188_ _08157_ _08149_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__or4_1
XFILLER_173_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15159_ _07803_ _07808_ _07813_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__o21a_1
XFILLER_99_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19967_ rbzero.pov.ready_buffer\[40\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-2\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__o221a_1
XFILLER_102_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18918_ _02583_ _02584_ _02574_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__and3b_1
X_19898_ rbzero.debug_overlay.playerY\[-7\] _03198_ _03202_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00991_ sky130_fd_sc_hd__o211a_1
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18849_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__nand2_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20811_ clknet_leaf_28_i_clk _00580_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20742_ clknet_leaf_33_i_clk _00511_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20673_ clknet_leaf_3_i_clk _00457_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20377__384 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__inv_2
XFILLER_177_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20076__112 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__inv_2
XFILLER_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21225_ clknet_leaf_73_i_clk _00994_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_117_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21156_ clknet_leaf_85_i_clk _00925_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21087_ net177 _00856_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20038_ _04990_ _04989_ _04037_ _02705_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__and4_1
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12860_ rbzero.wall_tracer.visualWallDist\[-8\] _05353_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__mux2_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _04121_ _04580_ _04588_ _04116_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__a31o_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ rbzero.wall_tracer.mapY\[6\] _05397_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__xor2_1
XFILLER_183_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _07259_ _07266_ _07264_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__a21oi_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11742_ _04519_ _04520_ _04021_ _04323_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a211oi_2
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14461_ _07195_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__or2b_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11673_ _04432_ _04448_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nor2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16200_ _08812_ _08844_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__or2_1
X_13412_ _06147_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__and2b_1
X_17180_ _07679_ vssd1 vssd1 vccd1 vccd1 _09771_ sky130_fd_sc_hd__clkbuf_4
X_10624_ _03651_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__clkbuf_1
X_14392_ _07111_ _07128_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__or2_1
XFILLER_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16131_ _08774_ _08775_ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__nand2_1
X_13343_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10555_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _03613_ vssd1 vssd1 vccd1 vccd1 _03615_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16062_ _08702_ _08703_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__and2_1
X_13274_ _05946_ _05877_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__xnor2_1
X_10486_ _03578_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15013_ _07676_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__nor2_1
X_12225_ _04986_ _04994_ net19 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__and3b_1
XFILLER_154_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ _03138_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__clkbuf_4
X_12156_ net46 _04918_ _04922_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a22o_1
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03321_ clknet_0__03321_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03321_
+ sky130_fd_sc_hd__clkbuf_16
X_11107_ _03904_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19752_ _03104_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12087_ net38 _04857_ _04838_ net48 vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a22o_1
X_16964_ rbzero.wall_tracer.texu\[4\] _09085_ _04035_ _09604_ vssd1 vssd1 vccd1 vccd1
+ _00515_ sky130_fd_sc_hd__o211a_1
XFILLER_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18703_ _05203_ _09283_ _05282_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__o21a_2
X_11038_ _03868_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__clkbuf_1
X_15915_ _07959_ _08042_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__nor2_1
X_19683_ rbzero.pov.spi_buffer\[17\] rbzero.pov.spi_buffer\[18\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16895_ _09528_ _09535_ vssd1 vssd1 vccd1 vccd1 _09536_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _02326_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__xnor2_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _08124_ _08490_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__and2_2
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ _01739_ _09027_ _02260_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__o21ai_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _05657_ _05658_ _05663_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__or4b_1
XFILLER_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15777_ _08416_ _08420_ _08421_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__a21o_1
XFILLER_166_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ _09939_ _09946_ _10081_ vssd1 vssd1 vccd1 vccd1 _10082_ sky130_fd_sc_hd__a21oi_2
X_14728_ _07463_ _07424_ _07433_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__mux2_1
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18496_ _02085_ _01985_ _02091_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14659_ _07103_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__clkinv_2
X_17447_ _10011_ _10013_ vssd1 vssd1 vccd1 vccd1 _10014_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17378_ _09943_ _09944_ vssd1 vssd1 vccd1 vccd1 _09945_ sky130_fd_sc_hd__xor2_1
XFILLER_203_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19117_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[2\] _02690_
+ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_173_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16329_ _08972_ _08973_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__or2b_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ rbzero.pov.spi_buffer\[55\] rbzero.pov.ready_buffer\[55\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21010_ clknet_leaf_67_i_clk _00779_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20725_ clknet_leaf_86_i_clk _00494_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20656_ clknet_leaf_93_i_clk _00440_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20587_ _07683_ _07692_ _07691_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10340_ rbzero.tex_r1\[48\] rbzero.tex_r1\[49\] _03494_ vssd1 vssd1 vccd1 vccd1 _03500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _04782_ _04783_ _04784_ _04266_ _04229_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__o221a_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21208_ clknet_leaf_16_i_clk _00977_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21139_ clknet_leaf_60_i_clk _00908_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_20130__161 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__inv_2
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13961_ _06134_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12912_ _05640_ _05642_ _05645_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__or4_2
X_15700_ _08343_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__or2_1
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16680_ _09160_ _09180_ _09322_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__a21boi_1
X_13892_ _06579_ _06628_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__or2_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _08269_ _08275_ _07990_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__mux2_2
X_12843_ rbzero.wall_tracer.rcp_sel\[2\] _05347_ _05348_ vssd1 vssd1 vccd1 vccd1 _05580_
+ sky130_fd_sc_hd__and3_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18350_ _02047_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ rbzero.wall_tracer.stepDistY\[3\] vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__inv_2
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ rbzero.map_rom.i_col\[4\] _05512_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__xor2_1
XFILLER_203_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14513_ _07233_ _07249_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__xnor2_1
X_17301_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09872_ sky130_fd_sc_hd__nor2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ rbzero.debug_overlay.playerY\[-3\] _04463_ _04502_ _04503_ vssd1 vssd1 vccd1
+ vccd1 _04504_ sky130_fd_sc_hd__a211o_1
X_15493_ _08115_ _08116_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18281_ _01756_ _01881_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a21o_1
XFILLER_203_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14444_ _07172_ _07174_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__nand2_1
X_17232_ _05413_ _09808_ _09810_ vssd1 vssd1 vccd1 vccd1 _09811_ sky130_fd_sc_hd__and3_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ _04420_ _04428_ _04433_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__or4_1
XFILLER_168_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17163_ rbzero.traced_texa\[-7\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a22o_1
XFILLER_122_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ rbzero.tex_g1\[51\] rbzero.tex_g1\[52\] _03635_ vssd1 vssd1 vccd1 vccd1 _03642_
+ sky130_fd_sc_hd__mux2_1
X_14375_ _07110_ _07111_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__xor2_1
XFILLER_156_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11587_ _04364_ _04365_ _04329_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16114_ _08740_ _08755_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__nor2_1
X_13326_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__inv_2
X_10538_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _03602_ vssd1 vssd1 vccd1 vccd1 _03606_
+ sky130_fd_sc_hd__mux2_1
X_17094_ _09474_ _09733_ vssd1 vssd1 vccd1 vccd1 _09734_ sky130_fd_sc_hd__xor2_1
XFILLER_171_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16045_ _08659_ _08661_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__or2_1
X_13257_ _05979_ _05909_ _05900_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__or3b_1
X_10469_ rbzero.tex_r0\[54\] rbzero.tex_r0\[53\] _03569_ vssd1 vssd1 vccd1 vccd1 _03570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20213__236 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__inv_2
XFILLER_142_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12208_ net15 net14 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and2b_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13188_ _05807_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__nand2_1
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ net50 rbzero.pov.ss_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
X_12139_ net8 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17996_ _01591_ _01606_ _01604_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a21o_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03304_ clknet_0__03304_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03304_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19735_ _03095_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16947_ _09448_ _09449_ vssd1 vssd1 vccd1 vccd1 _09588_ sky130_fd_sc_hd__nor2_1
XFILLER_93_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19666_ _03047_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16878_ _09408_ _09413_ vssd1 vssd1 vccd1 vccd1 _09519_ sky130_fd_sc_hd__and2b_1
XFILLER_93_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18617_ _02125_ _02128_ _02222_ _02223_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a31o_1
X_15829_ _08008_ _07941_ vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__nor2_1
XFILLER_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18548_ _02242_ _02244_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18479_ _01939_ _02071_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__nand2_1
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20510_ _03401_ _03403_ _03402_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__a21boi_1
XFILLER_178_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21490_ net411 _01259_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20441_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _03348_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_140_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19619__72 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20188__213 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__inv_2
XFILLER_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19634__86 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__inv_2
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11510_ _04129_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__buf_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20708_ clknet_leaf_3_i_clk _00015_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12490_ rbzero.wall_tracer.trackDistY\[-10\] _05241_ rbzero.wall_tracer.trackDistY\[-11\]
+ _05242_ _05244_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a221o_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ _04135_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__buf_4
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20639_ clknet_leaf_25_i_clk _00423_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14160_ _06864_ _06895_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__and2_1
XFILLER_109_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11372_ rbzero.row_render.size\[6\] _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__and2_1
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ _05838_ _05843_ _05820_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__mux2_1
X_10323_ rbzero.tex_r1\[56\] rbzero.tex_r1\[57\] _03483_ vssd1 vssd1 vccd1 vccd1 _03491_
+ sky130_fd_sc_hd__mux2_1
X_14091_ _06776_ _06662_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__nor2_1
XFILLER_140_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__buf_2
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17850_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nand2_1
XFILLER_117_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16801_ _09303_ _09305_ vssd1 vssd1 vccd1 vccd1 _09443_ sky130_fd_sc_hd__and2_1
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17781_ _01472_ _01484_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14993_ rbzero.wall_tracer.stepDistX\[3\] _07564_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07667_ sky130_fd_sc_hd__mux2_1
XFILLER_94_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19520_ _02983_ _02987_ _02996_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a21o_1
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16732_ _09223_ _09230_ _09373_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__a21oi_1
X_13944_ _06680_ _06677_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__nor2_1
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19451_ rbzero.wall_tracer.rayAddendY\[3\] _07855_ _02932_ _02933_ vssd1 vssd1 vccd1
+ vccd1 _02934_ sky130_fd_sc_hd__a22oi_1
X_13875_ _06605_ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_4
XFILLER_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _09303_ _09304_ _09275_ vssd1 vssd1 vccd1 vccd1 _09306_ sky130_fd_sc_hd__a21o_1
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18402_ _02062_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12826_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__buf_2
X_15614_ _08175_ _08176_ vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__nand2_4
X_19382_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nand2_1
XFILLER_188_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16594_ _09222_ _09236_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__xor2_1
XFILLER_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18333_ _02030_ _02029_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__and2b_1
XFILLER_72_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _08180_ _08189_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__nor2_1
X_12757_ _03929_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__nor2_1
XFILLER_188_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11708_ rbzero.debug_overlay.facingY\[-7\] _04455_ _04482_ _04486_ vssd1 vssd1 vccd1
+ vccd1 _04487_ sky130_fd_sc_hd__a211o_1
X_15476_ _08012_ _08026_ _08119_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__nand3_1
XFILLER_124_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18264_ _01951_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and2_1
XFILLER_187_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14427_ _07139_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__or2_1
X_17215_ rbzero.wall_tracer.mapX\[9\] _05525_ _09791_ vssd1 vssd1 vccd1 vccd1 _09796_
+ sky130_fd_sc_hd__o21a_1
X_11639_ _04415_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__nor2_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18195_ _01894_ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14358_ _07093_ _07094_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__nor2_1
X_17146_ _07555_ _09763_ rbzero.row_render.size\[8\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00536_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _06041_ _06045_ _05991_ _05978_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__or4_1
X_17077_ _09714_ _09716_ vssd1 vssd1 vccd1 vccd1 _09717_ sky130_fd_sc_hd__xor2_2
XFILLER_196_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14289_ _07023_ _07025_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__xor2_2
XFILLER_157_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16028_ _08617_ _08672_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__nor2_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17979_ _01678_ _01679_ _01680_ _09889_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__o31a_1
XFILLER_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19718_ _03086_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
X_20990_ clknet_leaf_38_i_clk _00759_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03318_ _03318_ vssd1 vssd1 vccd1 vccd1 clknet_0__03318_ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19649_ _03050_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21611_ net128 _01380_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21542_ net463 _01311_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21473_ net394 _01242_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20424_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03334_
+ sky130_fd_sc_hd__nor2_1
XFILLER_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03040_ clknet_0__03040_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03040_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_175_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _04763_ _04764_ _04345_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__mux2_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ rbzero.tex_b1\[21\] rbzero.tex_b1\[22\] _03817_ vssd1 vssd1 vccd1 vccd1 _03818_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13660_ _06363_ _06364_ _06360_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10872_ _03781_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20242__262 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__inv_2
XFILLER_204_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _05346_ _05349_ _05361_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__or4_1
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13591_ _06324_ _06326_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a21oi_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _07925_ rbzero.wall_tracer.stepDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _07975_
+ sky130_fd_sc_hd__nor2_1
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12542_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__xor2_1
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ rbzero.debug_overlay.playerY\[-6\] _07905_ vssd1 vssd1 vccd1 vccd1 _07906_
+ sky130_fd_sc_hd__or2_1
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ rbzero.wall_tracer.trackDistY\[9\] _05215_ _05217_ rbzero.wall_tracer.trackDistY\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__o22a_1
XFILLER_138_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03307_ clknet_0__03307_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03307_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14212_ _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__or2b_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17000_ _09521_ _09525_ vssd1 vssd1 vccd1 vccd1 _09640_ sky130_fd_sc_hd__nand2_1
XFILLER_172_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11424_ _04146_ _04203_ rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15192_ _07841_ _07842_ _07843_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__o211ai_2
XANTENNA_8 _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _06857_ _06878_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__nor2_1
XFILLER_137_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11355_ _04088_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _03474_ _03475_ _03478_ _03480_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__and4_1
X_14074_ _06803_ _06810_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__xor2_1
XFILLER_153_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18951_ _02594_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__clkbuf_4
XFILLER_180_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _04066_ sky130_fd_sc_hd__or2_1
XFILLER_152_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13025_ _05605_ _05604_ _05680_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__mux2_1
X_17902_ _01602_ _01603_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__and2_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18882_ _02553_ _02390_ rbzero.wall_tracer.trackDistY\[11\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00624_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17833_ _10254_ _10276_ _01536_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19613__67 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
X_17764_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__nor2_1
X_14976_ rbzero.wall_tracer.stepDistX\[-5\] _07650_ vssd1 vssd1 vccd1 vccd1 _07658_
+ sky130_fd_sc_hd__nor2_1
XFILLER_94_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20325__337 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__inv_2
XFILLER_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19503_ _02980_ _02981_ _02961_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a21o_1
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16715_ _08062_ _09217_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__nor2_1
X_13927_ _06031_ _06663_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__nor2_2
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17695_ _10255_ _10259_ vssd1 vssd1 vccd1 vccd1 _10260_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19434_ _02899_ _02914_ _02915_ _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a31o_1
X_16646_ _08215_ _08985_ _09138_ _08519_ vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__o22ai_1
X_13858_ _06564_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nand2_2
XFILLER_90_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19365_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or2_1
XFILLER_76_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ rbzero.wall_tracer.mapY\[9\] _05404_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__nor2_1
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16577_ _09161_ _09219_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__nand2_1
XFILLER_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13789_ _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__nor2_1
XFILLER_163_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18316_ _09889_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__or2_1
XFILLER_163_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15528_ _07894_ _05490_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__nand2_1
XFILLER_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19296_ rbzero.spi_registers.new_other\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
XFILLER_175_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18247_ _01943_ _01945_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__nand2_1
XFILLER_175_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15459_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__or2_2
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18178_ _08895_ _07916_ _07921_ _10134_ _01878_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__o311a_2
XFILLER_190_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17129_ _09759_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20070__107 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__inv_2
XFILLER_132_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20973_ clknet_leaf_53_i_clk _00742_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21525_ net446 _01294_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21456_ net377 _01225_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21387_ net308 _01156_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11140_ rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__inv_2
XFILLER_190_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20338_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__buf_1
XFILLER_123_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 o_gpout[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 o_tex_csb sky130_fd_sc_hd__buf_2
XFILLER_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _03885_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _07486_ _07455_ _07554_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a21boi_4
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _07473_ _07477_ _07493_ _07494_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__a31o_1
X_11973_ _04746_ _04747_ _04218_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__mux2_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20166__193 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__inv_2
XFILLER_205_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _09140_ _09143_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__xnor2_2
X_13712_ _06057_ _05982_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nor2_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ rbzero.tex_b1\[29\] rbzero.tex_b1\[30\] _03806_ vssd1 vssd1 vccd1 vccd1 _03809_
+ sky130_fd_sc_hd__mux2_1
X_14692_ _07379_ _07380_ _05931_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__a21o_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17480_ _09952_ _10040_ _10044_ vssd1 vssd1 vccd1 vccd1 _10046_ sky130_fd_sc_hd__and3_1
XFILLER_189_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _08549_ _08957_ vssd1 vssd1 vccd1 vccd1 _09076_ sky130_fd_sc_hd__xor2_4
XFILLER_60_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ _06340_ _06342_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__xnor2_1
X_10855_ _03772_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19150_ rbzero.otherx\[1\] _02710_ _02715_ _02714_ vssd1 vssd1 vccd1 vccd1 _00730_
+ sky130_fd_sc_hd__o211a_1
XFILLER_198_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13574_ _05920_ _06016_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__or2_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _08823_ _08059_ _09005_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__o21ai_1
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _03736_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18101_ _01781_ _01783_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__or2_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _03968_ _03998_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__nor2_1
X_15313_ _07945_ _07950_ _07956_ _07957_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__a22o_4
XFILLER_200_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16293_ _08806_ _08801_ _08805_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__a21bo_1
X_19081_ rbzero.pov.spi_buffer\[71\] rbzero.pov.ready_buffer\[71\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02673_ sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18032_ _01626_ _01628_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__nor2_1
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12456_ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__buf_4
X_15244_ rbzero.wall_tracer.wall\[1\] _03999_ _05280_ _03996_ vssd1 vssd1 vccd1 vccd1
+ _07891_ sky130_fd_sc_hd__a22o_1
XFILLER_173_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11407_ rbzero.row_render.size\[4\] _04150_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__xnor2_1
X_15175_ _07816_ _07824_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__a21oi_1
X_12387_ _03474_ _04814_ _04317_ _04809_ _05146_ _05145_ vssd1 vssd1 vccd1 vccd1 _05154_
+ sky130_fd_sc_hd__mux4_1
XFILLER_181_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _06827_ _06829_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11338_ _04097_ _04114_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__or3_1
XFILLER_125_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19983_ rbzero.pov.ready_buffer\[32\] _03247_ _03249_ rbzero.debug_overlay.facingY\[10\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__a221o_1
XFILLER_153_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ _06789_ _06793_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__xnor2_1
X_18934_ _02596_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11269_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _04049_
+ sky130_fd_sc_hd__nand2_1
XFILLER_141_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13008_ _05642_ _05744_ _05634_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18865_ _02530_ _02532_ _02531_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__o21bai_1
XFILLER_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17816_ _09114_ _09693_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__nor2_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18796_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__nand2_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17747_ _01443_ _01444_ _01450_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a21oi_1
X_14959_ rbzero.wall_tracer.trackDistX\[11\] rbzero.wall_tracer.trackDistY\[11\] _04019_
+ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__a21o_1
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17678_ _10241_ _10242_ vssd1 vssd1 vccd1 vccd1 _10243_ sky130_fd_sc_hd__xnor2_2
XFILLER_63_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19417_ _02885_ _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16629_ _09114_ _08204_ vssd1 vssd1 vccd1 vccd1 _09272_ sky130_fd_sc_hd__nor2_1
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19348_ rbzero.debug_overlay.vplaneY\[-9\] _07703_ _07855_ rbzero.wall_tracer.rayAddendY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a22o_1
XFILLER_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19279_ _02794_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21310_ net231 _01079_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21241_ clknet_leaf_81_i_clk _01010_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21172_ clknet_leaf_79_i_clk _00941_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20054_ rbzero.spi_registers.got_new_vinf _09753_ _02728_ _02555_ vssd1 vssd1 vccd1
+ vccd1 _01061_ sky130_fd_sc_hd__a31o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20308__321 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__inv_2
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ clknet_leaf_48_i_clk _00725_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20887_ clknet_leaf_83_i_clk _00656_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10640_ rbzero.tex_g1\[36\] rbzero.tex_g1\[37\] _03658_ vssd1 vssd1 vccd1 vccd1 _03660_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _03613_ vssd1 vssd1 vccd1 vccd1 _03623_
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _05034_ net25 _05051_ _05061_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__a311o_2
XFILLER_194_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21508_ net429 _01277_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[23\] sky130_fd_sc_hd__dfxtp_1
X_13290_ _05855_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20354__363 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__inv_2
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ net19 _04996_ _05010_ _04867_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__or4b_1
XFILLER_177_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21439_ net360 _01208_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _04813_ _04811_ _04006_ _03475_ _04910_ net9 vssd1 vssd1 vccd1 vccd1 _04943_
+ sky130_fd_sc_hd__mux4_1
XFILLER_162_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ net71 _03480_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__nand2_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16980_ _08160_ _09483_ vssd1 vssd1 vccd1 vccd1 _09620_ sky130_fd_sc_hd__nor2_1
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11054_ rbzero.tex_b0\[32\] rbzero.tex_b0\[31\] _03876_ vssd1 vssd1 vccd1 vccd1 _03877_
+ sky130_fd_sc_hd__mux2_1
X_15931_ _08573_ _08575_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_64_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18650_ _01739_ _09162_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__nor2_1
XFILLER_67_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _08152_ _08153_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__nand2_1
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17601_ _10165_ _10166_ vssd1 vssd1 vccd1 vccd1 _10167_ sky130_fd_sc_hd__or2b_2
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ rbzero.wall_tracer.stepDistY\[-4\] _07541_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07542_ sky130_fd_sc_hd__mux2_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18581_ _02272_ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__and2_1
XFILLER_64_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15793_ _08413_ _08437_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__xnor2_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_102 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_102/HI zeros[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_123_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17532_ _10096_ _10097_ vssd1 vssd1 vccd1 vccd1 _10098_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_79_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xtop_ew_algofoogle_113 vssd1 vssd1 vccd1 vccd1 ones[7] top_ew_algofoogle_113/LO sky130_fd_sc_hd__conb_1
X_14744_ _07385_ _07387_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__or2b_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _04726_ _04728_ _04731_ _04332_ _04241_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__a221o_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ rbzero.tex_b1\[37\] rbzero.tex_b1\[38\] _03795_ vssd1 vssd1 vccd1 vccd1 _03800_
+ sky130_fd_sc_hd__mux2_1
X_17463_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _10030_ sky130_fd_sc_hd__nor2_1
X_14675_ _06724_ _06761_ _07411_ _07340_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o211a_1
X_11887_ rbzero.color_sky\[3\] rbzero.color_floor\[3\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04664_ sky130_fd_sc_hd__mux2_1
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19202_ rbzero.spi_registers.new_sky\[4\] rbzero.spi_registers.got_new_sky _02711_
+ _02741_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a31o_1
X_16414_ _09056_ _09058_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__xnor2_2
X_13626_ _06361_ _06362_ _06078_ _05982_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a211o_1
X_10838_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _03762_ vssd1 vssd1 vccd1 vccd1 _03764_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17394_ _09661_ _08356_ _09960_ vssd1 vssd1 vccd1 vccd1 _09961_ sky130_fd_sc_hd__or3_1
XFILLER_73_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _02701_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__clkbuf_1
X_16345_ _08987_ _08989_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__xnor2_2
X_13557_ _05995_ _06113_ _06045_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a21o_1
X_10769_ _03727_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19064_ _02664_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
X_12508_ rbzero.wall_tracer.trackDistX\[-4\] vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__inv_2
X_13488_ _06197_ _06198_ _06224_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o21ai_1
XFILLER_160_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16276_ _08869_ _08919_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__or2_1
XFILLER_200_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18015_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__nand2_1
X_15227_ rbzero.wall_tracer.rayAddendX\[9\] _00013_ _07831_ _07875_ _07877_ vssd1
+ vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_17_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12439_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__buf_4
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158_ _07800_ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__xor2_1
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _06763_ _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15089_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__nor2_1
X_19966_ rbzero.pov.ready_buffer\[39\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-3\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__a221o_1
XFILLER_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18917_ rbzero.spi_registers.spi_counter\[3\] _02580_ vssd1 vssd1 vccd1 vccd1 _02584_
+ sky130_fd_sc_hd__or2_1
XFILLER_122_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19897_ rbzero.pov.ready_buffer\[46\] _02823_ _03193_ _03201_ vssd1 vssd1 vccd1 vccd1
+ _03202_ sky130_fd_sc_hd__a211o_1
XFILLER_171_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18848_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__or2_1
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20182__208 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__inv_2
XFILLER_110_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18779_ _09812_ _09597_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__nand2_1
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20810_ clknet_leaf_28_i_clk _00579_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20741_ clknet_leaf_10_i_clk _00510_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.side
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20672_ clknet_leaf_12_i_clk _00456_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21224_ clknet_leaf_73_i_clk _00993_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
X_21155_ clknet_leaf_83_i_clk _00924_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21086_ net176 _00855_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20037_ _03277_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _04582_ _04584_ _04587_ _04208_ _04142_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a221o_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05532_ _05283_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__nor2_2
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _03478_ _04026_ _04047_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a21oi_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ clknet_leaf_67_i_clk _00708_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14460_ _07170_ _07182_ _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o21ai_1
X_11672_ _04004_ _04419_ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__and3b_1
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13411_ _06144_ _06091_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10623_ rbzero.tex_g1\[44\] rbzero.tex_g1\[45\] _03647_ vssd1 vssd1 vccd1 vccd1 _03651_
+ sky130_fd_sc_hd__mux2_1
X_14391_ _06675_ _06761_ _07108_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__o21ai_1
XFILLER_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20278__294 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__inv_2
X_13342_ _06053_ _06056_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and2_1
XFILLER_167_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16130_ _08773_ _08772_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__or2b_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10554_ _03614_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13273_ _05973_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nor2_1
X_16061_ _08594_ _08705_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__nor2_1
X_10485_ rbzero.tex_r0\[46\] rbzero.tex_r0\[45\] _03569_ vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ _04987_ _04988_ _04991_ _04993_ net16 _04960_ vssd1 vssd1 vccd1 vccd1 _04994_
+ sky130_fd_sc_hd__mux4_1
X_15012_ rbzero.wall_tracer.state\[14\] _04037_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__nand2_2
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19820_ _03140_ rbzero.pov.ready_buffer\[59\] _03141_ vssd1 vssd1 vccd1 vccd1 _03142_
+ sky130_fd_sc_hd__mux2_1
X_12155_ net51 _04904_ net47 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a21o_1
XFILLER_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11106_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _03898_ vssd1 vssd1 vccd1 vccd1 _03904_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03320_ clknet_0__03320_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03320_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19751_ rbzero.pov.spi_buffer\[49\] rbzero.pov.spi_buffer\[50\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
X_12086_ net43 _04857_ _04838_ net41 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a22o_1
X_16963_ _09085_ _09603_ vssd1 vssd1 vccd1 vccd1 _09604_ sky130_fd_sc_hd__nand2_1
X_18702_ _09808_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__nand2_1
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11037_ rbzero.tex_b0\[40\] rbzero.tex_b0\[39\] _03865_ vssd1 vssd1 vccd1 vccd1 _03868_
+ sky130_fd_sc_hd__mux2_1
X_15914_ _07923_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__or3_1
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19682_ _03067_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16894_ _09533_ _09534_ vssd1 vssd1 vccd1 vccd1 _09535_ sky130_fd_sc_hd__xor2_1
XFILLER_65_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18633_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__xnor2_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _07945_ rbzero.wall_tracer.stepDistX\[-11\] vssd1 vssd1 vccd1 vccd1 _08490_
+ sky130_fd_sc_hd__nand2_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ _01739_ _09027_ _02260_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__or3_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _08062_ _08158_ _08150_ _08054_ vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__o22a_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand2_2
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _09664_ _09665_ _09945_ vssd1 vssd1 vccd1 vccd1 _10081_ sky130_fd_sc_hd__a21oi_1
X_14727_ _05892_ _07395_ _07398_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__o21a_1
X_19583__39 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
X_11939_ _04712_ _04713_ _04714_ _04247_ _04306_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o221a_1
X_18495_ _02185_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__xor2_1
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17446_ _09680_ _09721_ _10012_ vssd1 vssd1 vccd1 vccd1 _10013_ sky130_fd_sc_hd__a21o_1
X_14658_ _07352_ _07362_ _05779_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13609_ _06281_ _06283_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17377_ _09245_ _08427_ vssd1 vssd1 vccd1 vccd1 _09944_ sky130_fd_sc_hd__nor2_1
X_14589_ _07131_ _07325_ _07206_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19116_ _02692_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16328_ _07981_ _07989_ _08189_ _08971_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__or4_1
XFILLER_158_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19047_ _02655_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16259_ _08892_ _08899_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19949_ rbzero.pov.ready _02707_ _02820_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__and3_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20724_ clknet_leaf_86_i_clk _00493_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_180_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20655_ clknet_leaf_93_i_clk _00439_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20586_ rbzero.wall_tracer.rayAddendX\[-7\] _03443_ _07756_ _03455_ vssd1 vssd1 vccd1
+ vccd1 _01426_ sky130_fd_sc_hd__a22o_1
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21207_ clknet_leaf_17_i_clk _00976_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21138_ clknet_leaf_61_i_clk _00907_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13960_ _06696_ _06671_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__nor2_1
X_21069_ net159 _00838_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12911_ _05646_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__xnor2_4
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13891_ _06572_ _06627_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ _07951_ rbzero.wall_tracer.stepDistY\[-1\] _08272_ _08274_ vssd1 vssd1 vccd1
+ vccd1 _08275_ sky130_fd_sc_hd__a22oi_4
X_12842_ _04030_ _05346_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a21o_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _08193_ _08205_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__xnor2_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _05518_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _09871_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _07247_ _07248_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__nor2_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18280_ _01882_ _01877_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__and2b_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ rbzero.debug_overlay.playerY\[0\] _04459_ _04460_ rbzero.debug_overlay.playerY\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a22o_1
XFILLER_202_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15492_ _08131_ _08136_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__xor2_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17231_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09809_ vssd1 vssd1 vccd1 vccd1 _09810_ sky130_fd_sc_hd__a21o_1
XFILLER_30_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14443_ _07176_ _07178_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__a21oi_1
X_11655_ gpout0.hpos\[6\] _04430_ _04431_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__and3_1
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17162_ _07706_ vssd1 vssd1 vccd1 vccd1 _09768_ sky130_fd_sc_hd__buf_2
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _03641_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__clkbuf_1
X_14374_ _06689_ _07072_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__nor2_1
X_11586_ rbzero.tex_r1\[25\] rbzero.tex_r1\[24\] _04342_ vssd1 vssd1 vccd1 vccd1 _04365_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16113_ _08737_ _08757_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__nor2_1
X_13325_ _06059_ _06060_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a21oi_1
X_10537_ _03605_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17093_ _09730_ _09732_ vssd1 vssd1 vccd1 vccd1 _09733_ sky130_fd_sc_hd__xor2_2
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16044_ _08683_ _08688_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__or2b_1
X_13256_ _05988_ _05989_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__and3_1
X_10468_ _03557_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12207_ net17 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__inv_2
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13187_ _05695_ _05724_ _05793_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__mux2_1
X_10399_ rbzero.tex_r1\[20\] rbzero.tex_r1\[21\] _03527_ vssd1 vssd1 vccd1 vccd1 _03531_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ net8 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__inv_2
X_19803_ _03130_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17995_ _01566_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03303_ clknet_0__03303_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03303_
+ sky130_fd_sc_hd__clkbuf_16
X_12069_ _04840_ net61 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__or2_1
X_19734_ rbzero.pov.spi_buffer\[41\] rbzero.pov.spi_buffer\[42\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
X_16946_ _09476_ _09586_ vssd1 vssd1 vccd1 vccd1 _09587_ sky130_fd_sc_hd__xnor2_1
X_19665_ _03058_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16877_ _09393_ _09402_ _09400_ vssd1 vssd1 vccd1 vccd1 _09518_ sky130_fd_sc_hd__a21o_1
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18616_ _02125_ _02128_ _02222_ _02223_ _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a311oi_2
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _07995_ _07981_ _07989_ _07931_ vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__o22ai_1
XFILLER_53_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18547_ _02151_ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__xnor2_1
X_15759_ _08396_ _08392_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__or2b_1
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18478_ _02174_ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nand2_1
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17429_ _08519_ _09699_ vssd1 vssd1 vccd1 vccd1 _09996_ sky130_fd_sc_hd__or2_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20440_ _03272_ _03346_ _03347_ _03327_ rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1
+ _01388_ sky130_fd_sc_hd__a32o_1
XFILLER_193_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__buf_1
XFILLER_147_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20707_ clknet_leaf_2_i_clk _00013_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11440_ _04215_ _04216_ _04219_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
X_20638_ clknet_leaf_27_i_clk _00422_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11371_ rbzero.row_render.size\[5\] rbzero.row_render.size\[4\] _04150_ vssd1 vssd1
+ vccd1 vccd1 _04151_ sky130_fd_sc_hd__or3_1
X_20569_ gpout0.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nor2_1
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ _05798_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__inv_2
X_10322_ _03490_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
X_14090_ _06805_ _06740_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__nor2_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13041_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16800_ _09415_ _09441_ vssd1 vssd1 vccd1 vccd1 _09442_ sky130_fd_sc_hd__xnor2_2
XFILLER_121_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17780_ _01482_ _01483_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__and2b_1
XFILLER_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14992_ _07666_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16731_ _09092_ _09095_ _09229_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__a21oi_1
X_13943_ _06161_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__clkbuf_4
XFILLER_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19450_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.debug_overlay.vplaneY\[-6\] _02930_
+ _02931_ _03913_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__o41a_1
XFILLER_207_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16662_ _09275_ _09303_ _09304_ vssd1 vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__nand3_1
X_13874_ _06607_ _06610_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and2b_1
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18401_ _02065_ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__xor2_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15613_ _08257_ _08238_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__nor2_1
X_19381_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__or2_1
X_12825_ _05561_ _05492_ _05493_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or3_4
XFILLER_188_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16593_ _09234_ _09235_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__nor2_1
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18332_ _02029_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__and2b_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15544_ _08147_ rbzero.wall_tracer.stepDistX\[2\] _08188_ vssd1 vssd1 vccd1 vccd1
+ _08189_ sky130_fd_sc_hd__a21boi_4
XFILLER_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _05496_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__inv_2
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18263_ _01960_ _01962_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__xor2_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11707_ rbzero.debug_overlay.facingY\[-8\] _04466_ _04483_ _04485_ vssd1 vssd1 vccd1
+ vccd1 _04486_ sky130_fd_sc_hd__a211o_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15475_ _08012_ _08026_ _08119_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__a21o_1
X_12687_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] _05434_
+ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__and3_1
XFILLER_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17214_ rbzero.wall_tracer.mapX\[9\] _09781_ _09779_ _09795_ vssd1 vssd1 vccd1 vccd1
+ _00574_ sky130_fd_sc_hd__a22o_1
X_14426_ _06724_ _06663_ _07138_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__o21a_1
XFILLER_128_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11638_ _04024_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or2_1
X_18194_ _01770_ _01771_ _01772_ _01775_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a31o_1
XFILLER_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17145_ _07552_ _09763_ rbzero.row_render.size\[7\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00535_ sky130_fd_sc_hd__a2bb2o_1
X_14357_ _07090_ _07092_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__and2_1
XFILLER_128_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _04136_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__clkbuf_4
X_13308_ _05899_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20137__168 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__inv_2
X_17076_ _09559_ _09570_ _09715_ vssd1 vssd1 vccd1 vccd1 _09716_ sky130_fd_sc_hd__a21oi_2
X_14288_ _06757_ _06797_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__a21boi_2
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16027_ _08619_ _08671_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__and2b_1
X_13239_ _05974_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nor2_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17978_ _01678_ _01679_ _01680_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19717_ rbzero.pov.spi_buffer\[33\] rbzero.pov.spi_buffer\[34\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
X_16929_ _09567_ _09569_ vssd1 vssd1 vccd1 vccd1 _09570_ sky130_fd_sc_hd__xor2_2
Xclkbuf_0__03317_ _03317_ vssd1 vssd1 vccd1 vccd1 clknet_0__03317_ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19648_ rbzero.pov.spi_buffer\[0\] rbzero.pov.spi_buffer\[1\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20302__316 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__inv_2
XFILLER_129_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21610_ net127 _01379_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21541_ net462 _01310_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21472_ net393 _01241_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20423_ _03329_ _03330_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__and2_1
XFILLER_179_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10940_ _03646_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__clkbuf_4
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ rbzero.tex_b1\[54\] rbzero.tex_b1\[55\] _03773_ vssd1 vssd1 vccd1 vccd1 _03781_
+ sky130_fd_sc_hd__mux2_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__and2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _06304_ _06323_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__nor2_1
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12541_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] _05290_
+ _05293_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a221o_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_i_clk clknet_1_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_197_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__or3_1
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ _05221_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__03306_ clknet_0__03306_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03306_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ _06932_ _06945_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__xnor2_1
X_11423_ rbzero.row_render.size\[10\] rbzero.row_render.size\[9\] _04153_ _04202_
+ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__or4_2
X_15191_ _07785_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _07844_
+ sky130_fd_sc_hd__or2_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14142_ _06857_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__xor2_1
X_11354_ rbzero.floor_leak\[4\] _04121_ _04116_ rbzero.floor_leak\[5\] vssd1 vssd1
+ vccd1 vccd1 _04134_ sky130_fd_sc_hd__o22a_1
XFILLER_180_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__buf_6
XFILLER_193_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14073_ _06776_ _06740_ _06804_ _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__o31a_1
XFILLER_141_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11285_ rbzero.texV\[6\] _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__xor2_1
X_18950_ _02604_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13024_ _05677_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__inv_2
X_17901_ _01602_ _01603_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__nor2_1
XFILLER_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18881_ _05532_ _02552_ _02399_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__o21a_1
XFILLER_79_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17832_ _10273_ _10275_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__or2b_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ _09249_ _09359_ _10206_ _10205_ _09391_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__o32a_1
X_14975_ _00008_ _07530_ _07657_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19502_ _02905_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02981_
+ sky130_fd_sc_hd__nand2_1
X_16714_ _09354_ _09355_ vssd1 vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__xnor2_1
X_13926_ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__clkbuf_4
XFILLER_130_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17694_ _09292_ _09695_ _08895_ vssd1 vssd1 vccd1 vccd1 _10259_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19433_ _03912_ _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nand2_1
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16645_ _09284_ _09287_ _05210_ vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__a21o_1
X_13857_ _06273_ _06593_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__xor2_1
XFILLER_35_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19364_ _02851_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__or2b_1
X_12808_ rbzero.wall_tracer.mapY\[9\] _05404_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__and2_1
X_16576_ _09214_ _09218_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__xnor2_2
X_13788_ _06507_ _06523_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__nand2_1
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315_ _02013_ _02014_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15527_ _07560_ _08171_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12739_ _05440_ _05465_ _05462_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a21boi_1
X_19295_ _02803_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18246_ _01943_ _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__or2_1
X_15458_ _05197_ rbzero.wall_tracer.stepDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _08103_
+ sky130_fd_sc_hd__nor2_2
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14409_ _06239_ _07111_ _07145_ _07131_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o31a_1
X_18177_ _08895_ _08767_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _07990_ _05496_ _08028_ _08033_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__o31a_2
X_17128_ _04446_ _09750_ _09758_ vssd1 vssd1 vccd1 vccd1 _09759_ sky130_fd_sc_hd__and3_1
XFILLER_171_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17059_ _09283_ rbzero.wall_tracer.stepDistY\[11\] _08235_ _09698_ vssd1 vssd1 vccd1
+ vccd1 _09699_ sky130_fd_sc_hd__a22oi_4
XFILLER_132_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20972_ clknet_leaf_53_i_clk _00741_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21524_ net445 _01293_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21455_ net376 _01224_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21386_ net307 _01155_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 o_gpout[4] sky130_fd_sc_hd__clkbuf_1
X_11070_ rbzero.tex_b0\[24\] rbzero.tex_b0\[23\] _03876_ vssd1 vssd1 vccd1 vccd1 _03885_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 o_tex_oeb0 sky130_fd_sc_hd__buf_2
XFILLER_153_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20056__94 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__inv_2
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _07102_ _05952_ _05844_ _07366_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__and4b_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _04342_ vssd1 vssd1 vccd1 vccd1 _04747_
+ sky130_fd_sc_hd__mux2_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _06442_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__xor2_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _03808_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14691_ _07378_ _07413_ _07414_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o31a_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16430_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerX\[-7\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__mux2_1
X_13642_ _06347_ _06373_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__xnor2_2
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10854_ rbzero.tex_b1\[62\] rbzero.tex_b1\[63\] _03691_ vssd1 vssd1 vccd1 vccd1 _03772_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _08823_ _08058_ _09005_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__or3_1
XFILLER_197_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13573_ _05823_ _05939_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__or2_1
XFILLER_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10785_ rbzero.tex_g0\[32\] rbzero.tex_g0\[31\] _03729_ vssd1 vssd1 vccd1 vccd1 _03736_
+ sky130_fd_sc_hd__mux2_1
X_18100_ _01667_ _01800_ _01787_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a21o_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ rbzero.wall_tracer.visualWallDist\[-4\] _07925_ _05207_ vssd1 vssd1 vccd1
+ vccd1 _07957_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19080_ _02672_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
X_12524_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__inv_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16292_ _08764_ _08807_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__xor2_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18031_ _01698_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__xor2_1
X_15243_ _07890_ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12455_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11406_ _04151_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__nand2_1
XFILLER_125_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15174_ _07785_ rbzero.wall_tracer.rayAddendX\[6\] vssd1 vssd1 vccd1 vccd1 _07828_
+ sky130_fd_sc_hd__xnor2_1
X_12386_ net35 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__inv_2
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14125_ _06846_ _06847_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__xor2_1
X_20331__342 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__inv_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ _04096_ _04075_ _04093_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__nor3_1
XFILLER_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19982_ rbzero.pov.ready_buffer\[31\] _03247_ _03249_ rbzero.debug_overlay.facingY\[0\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__a221o_1
XFILLER_158_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14056_ _06787_ _06791_ _06792_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__o21ai_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18933_ rbzero.pov.spi_buffer\[0\] rbzero.pov.ready_buffer\[0\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
X_11268_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _04048_
+ sky130_fd_sc_hd__nand2_1
XFILLER_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007_ _05622_ _05635_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__xnor2_2
XFILLER_140_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18864_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__nand2_1
X_11199_ rbzero.map_rom.f4 _03933_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17815_ _01514_ _01518_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__xnor2_1
X_18795_ _02478_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17746_ _01448_ _01449_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__nand2_1
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14958_ _04019_ _07647_ _07648_ _07642_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__o211a_1
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13909_ _05752_ _06201_ _06621_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17677_ _10094_ _08057_ vssd1 vssd1 vccd1 vccd1 _10242_ sky130_fd_sc_hd__nor2_1
X_14889_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.trackDistX\[-10\]
+ _07592_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19416_ _02899_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__nand2_1
X_16628_ _09119_ _09270_ vssd1 vssd1 vccd1 vccd1 _09271_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16559_ rbzero.wall_tracer.texu\[1\] _09085_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__or2_1
X_19347_ _02826_ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__xnor2_1
X_19278_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_leak\[1\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XFILLER_30_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18229_ _01838_ _01852_ _01850_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a21o_1
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21240_ clknet_leaf_81_i_clk _01009_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21171_ clknet_leaf_78_i_clk _00940_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20053_ _03285_ _03288_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__nor2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19589__45 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ clknet_leaf_41_i_clk _00724_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ clknet_leaf_82_i_clk _00655_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _03622_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21507_ net428 _01276_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ _04960_ _04961_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__nand2_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21438_ net359 _01207_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ net11 _04908_ _04937_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a31o_1
XFILLER_150_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21369_ net290 _01138_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11122_ _03911_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_8
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11053_ _03717_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__clkbuf_4
X_15930_ _08498_ _08574_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__xnor2_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15861_ _08489_ _08505_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__or2b_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_17600_ _10037_ _10038_ _10164_ vssd1 vssd1 vccd1 vccd1 _10166_ sky130_fd_sc_hd__a21o_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _07486_ _07455_ _07539_ _07527_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__a221o_4
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18580_ _02275_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__xor2_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _08435_ _08436_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__and2_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _08275_ _08356_ vssd1 vssd1 vccd1 vccd1 _10097_ sky130_fd_sc_hd__nor2_1
XFILLER_91_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14743_ _07475_ _07476_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__mux2_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_103 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_103/HI zeros[13]
+ sky130_fd_sc_hd__conb_1
X_11955_ _04729_ _04730_ _04329_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__mux2_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_114 vssd1 vssd1 vccd1 vccd1 ones[8] top_ew_algofoogle_114/LO sky130_fd_sc_hd__conb_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _03799_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17462_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _10029_ sky130_fd_sc_hd__nand2_1
X_14674_ _06239_ _07149_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__nor2_1
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11886_ _04628_ _04206_ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__or3b_4
XFILLER_189_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16413_ _08169_ _08469_ _09057_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__a21o_1
X_19201_ _02747_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__clkbuf_1
X_13625_ _06041_ _06031_ _06285_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__o21ai_1
X_10837_ _03763_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17393_ _09663_ _09959_ vssd1 vssd1 vccd1 vccd1 _09960_ sky130_fd_sc_hd__xnor2_1
X_19132_ rbzero.spi_registers.sclk_buffer\[1\] rbzero.spi_registers.sclk_buffer\[0\]
+ _05189_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XFILLER_160_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16344_ _08237_ _08239_ _08229_ _08988_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__o31a_1
XFILLER_197_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13556_ _06057_ _05940_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ rbzero.tex_g0\[40\] rbzero.tex_g0\[39\] _03718_ vssd1 vssd1 vccd1 vccd1 _03727_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19063_ rbzero.pov.spi_buffer\[62\] rbzero.pov.ready_buffer\[62\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_12507_ _05258_ rbzero.wall_tracer.trackDistX\[-1\] _05251_ rbzero.wall_tracer.trackDistX\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a22o_1
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16275_ _08869_ _08919_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__nand2_1
X_13487_ _06209_ _06223_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10699_ _03690_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18014_ _01474_ _08423_ _01596_ _01594_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__o31a_1
X_15226_ _07858_ _07862_ _07876_ _04034_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__a211o_1
XFILLER_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12438_ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__buf_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15157_ _07785_ _04462_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__xor2_1
X_12369_ _05115_ _05123_ _05130_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__or4_2
XFILLER_141_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _06704_ _06668_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__nor2_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15088_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__and2_1
X_19965_ _02695_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14039_ _05984_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__buf_2
X_18916_ rbzero.spi_registers.spi_counter\[3\] _02580_ vssd1 vssd1 vccd1 vccd1 _02583_
+ sky130_fd_sc_hd__and2_1
XFILLER_141_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19896_ _08004_ _03141_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__nor2_1
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18847_ _02523_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18778_ _02463_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17729_ _10292_ _10293_ vssd1 vssd1 vccd1 vccd1 _10294_ sky130_fd_sc_hd__nor2_2
XFILLER_208_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20740_ clknet_leaf_14_i_clk _00509_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20671_ clknet_leaf_12_i_clk _00455_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21223_ clknet_leaf_73_i_clk _00992_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_191_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21154_ clknet_leaf_83_i_clk _00923_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20105_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__buf_1
X_21085_ net175 _00854_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20036_ _03275_ _03276_ _05190_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__and3b_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04041_ _04497_ _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o21ai_2
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ clknet_leaf_67_i_clk _00707_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_187_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _04448_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__inv_2
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ clknet_leaf_66_i_clk _00638_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _06138_ _06141_ _06146_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__o21a_1
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10622_ _03650_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__clkbuf_1
X_14390_ _07120_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__xor2_1
X_13341_ _06045_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ rbzero.tex_r0\[14\] rbzero.tex_r0\[13\] _03613_ vssd1 vssd1 vccd1 vccd1 _03614_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16060_ _07929_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__clkbuf_4
X_13272_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__buf_2
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _03577_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15011_ _03912_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__clkbuf_4
X_12223_ _04891_ _04992_ _04890_ _04892_ _04969_ _04966_ vssd1 vssd1 vccd1 vccd1 _04993_
+ sky130_fd_sc_hd__mux4_1
XFILLER_154_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ _04907_ _04905_ _04921_ _04923_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a2111o_2
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _03903_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19750_ _03047_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12085_ net3 _04852_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__nor2_2
X_16962_ _09470_ _09602_ vssd1 vssd1 vccd1 vccd1 _09603_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18701_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _02395_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a21o_1
X_11036_ _03867_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__clkbuf_1
X_15913_ _08556_ _08552_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__xor2_1
X_19681_ rbzero.pov.spi_buffer\[16\] rbzero.pov.spi_buffer\[17\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
X_16893_ _09395_ _09396_ _09397_ _09398_ vssd1 vssd1 vccd1 vccd1 _09534_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15844_ _08487_ _08488_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__nand2_1
X_18632_ _08159_ _09138_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__nor2_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18563_ _08257_ _09162_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__or2_1
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15775_ _08054_ _08419_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__nor2_1
X_12987_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__inv_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _07462_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__clkbuf_1
X_17514_ _10070_ _10079_ vssd1 vssd1 vccd1 vccd1 _10080_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11938_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _04263_ vssd1 vssd1 vccd1 vccd1 _04714_
+ sky130_fd_sc_hd__mux2_1
X_18494_ _02186_ _02191_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__xor2_1
XFILLER_33_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _09718_ _09720_ vssd1 vssd1 vccd1 vccd1 _10012_ sky130_fd_sc_hd__nor2_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__buf_2
XFILLER_159_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11869_ rbzero.tex_g1\[19\] rbzero.tex_g1\[18\] _04336_ vssd1 vssd1 vccd1 vccd1 _04646_
+ sky130_fd_sc_hd__mux2_1
X_13608_ _05988_ _06337_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__o21ba_1
XFILLER_177_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ _09941_ _09942_ vssd1 vssd1 vccd1 vccd1 _09943_ sky130_fd_sc_hd__or2b_1
X_14588_ _07116_ _07324_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__or2_1
XFILLER_159_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19115_ rbzero.spi_registers.spi_cmd\[0\] rbzero.spi_registers.spi_cmd\[1\] _02690_
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
X_16327_ _08180_ _08189_ _08971_ _08170_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__o22a_1
X_13539_ _06232_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__xor2_1
XFILLER_201_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19046_ rbzero.pov.spi_buffer\[54\] rbzero.pov.ready_buffer\[54\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
X_16258_ _08889_ _08891_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__nor2_1
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15209_ _07850_ _07854_ _07860_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__and3_1
XFILLER_173_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16189_ _08820_ _08826_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19948_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__clkbuf_4
XFILLER_96_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19879_ _03184_ _03187_ _02714_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__o21a_1
XFILLER_114_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20723_ clknet_leaf_90_i_clk _00492_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20654_ clknet_leaf_93_i_clk _00438_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20585_ _07689_ _03454_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_78_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21206_ clknet_leaf_16_i_clk _00975_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21137_ clknet_leaf_61_i_clk _00906_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21068_ net158 _00837_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20019_ net59 _03263_ _03264_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__a21oi_1
X_12910_ _05615_ _05601_ _05566_ _05563_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__o211a_1
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13890_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__inv_2
XFILLER_150_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12841_ rbzero.wall_tracer.visualWallDist\[-4\] _05570_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05578_ sky130_fd_sc_hd__a21o_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15560_ _08194_ _08204_ vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__nor2_1
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ rbzero.map_rom.f1 _05517_ _05414_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__mux2_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14511_ _07234_ _07246_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__and2_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ gpout0.vpos\[3\] _04041_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__nand2_1
X_15491_ _08059_ _08135_ vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__nor2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09807_ vssd1 vssd1 vccd1 vccd1 _09809_ sky130_fd_sc_hd__o21ai_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14442_ _07108_ _07063_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__and2b_1
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _04422_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__nor2_1
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17161_ rbzero.traced_texa\[-8\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a22o_1
X_10605_ rbzero.tex_g1\[52\] rbzero.tex_g1\[53\] _03635_ vssd1 vssd1 vccd1 vccd1 _03641_
+ sky130_fd_sc_hd__mux2_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14373_ _07108_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__xnor2_2
XFILLER_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ rbzero.tex_r1\[27\] rbzero.tex_r1\[26\] _04262_ vssd1 vssd1 vccd1 vccd1 _04364_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _08725_ _08734_ _08736_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__and3_1
X_13324_ _05944_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10536_ rbzero.tex_r0\[22\] rbzero.tex_r0\[21\] _03602_ vssd1 vssd1 vccd1 vccd1 _03605_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17092_ _09476_ _09586_ _09731_ vssd1 vssd1 vccd1 vccd1 _09732_ sky130_fd_sc_hd__a21oi_2
XFILLER_127_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16043_ _08284_ _08128_ _08623_ _08687_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__o31ai_2
X_13255_ _05990_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nand2_1
XFILLER_143_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10467_ _03568_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ net17 _04968_ _04971_ _04975_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o211a_1
X_13186_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__clkbuf_4
X_10398_ _03530_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19802_ rbzero.pov.mosi rbzero.pov.mosi_buffer\[0\] _05189_ vssd1 vssd1 vccd1 vccd1
+ _03130_ sky130_fd_sc_hd__mux2_1
X_12137_ net10 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__inv_2
X_17994_ _01694_ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__nor2_1
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03302_ clknet_0__03302_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03302_
+ sky130_fd_sc_hd__clkbuf_16
X_19733_ _03094_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
X_12068_ net2 vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__clkbuf_4
XFILLER_81_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16945_ _09583_ _09585_ vssd1 vssd1 vccd1 vccd1 _09586_ sky130_fd_sc_hd__xor2_1
XFILLER_133_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _03858_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19664_ rbzero.pov.spi_buffer\[8\] rbzero.pov.spi_buffer\[9\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
XFILLER_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16876_ _09477_ _09516_ vssd1 vssd1 vccd1 vccd1 _09517_ sky130_fd_sc_hd__xnor2_1
X_18615_ _02310_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__or2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _08471_ _08023_ vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__xor2_1
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15758_ _08393_ _08395_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__or2_1
X_18546_ _10248_ _01524_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__nor2_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14709_ _05742_ _07400_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__nor2_1
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15689_ _08330_ _08333_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__nand2_1
X_18477_ _10239_ _09215_ _02173_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17428_ _05211_ _08215_ _09565_ vssd1 vssd1 vccd1 vccd1 _09995_ sky130_fd_sc_hd__or3_1
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17359_ _09924_ _09925_ vssd1 vssd1 vccd1 vccd1 _09926_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19029_ rbzero.pov.spi_buffer\[46\] rbzero.pov.ready_buffer\[46\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_161_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20114__147 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__inv_2
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20706_ clknet_leaf_4_i_clk _00490_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20195__219 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__inv_2
XFILLER_200_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20637_ clknet_leaf_27_i_clk _00421_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ rbzero.row_render.size\[3\] _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__or2_1
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20568_ rbzero.traced_texVinit\[11\] _03443_ _07756_ _01552_ vssd1 vssd1 vccd1 vccd1
+ _01419_ sky130_fd_sc_hd__a22o_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10321_ rbzero.tex_r1\[57\] rbzero.tex_r1\[58\] _03483_ vssd1 vssd1 vccd1 vccd1 _03490_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20499_ _03390_ _03394_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nand2_1
X_13040_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20089__124 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__inv_2
XFILLER_59_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14991_ rbzero.wall_tracer.stepDistX\[2\] _07562_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07666_ sky130_fd_sc_hd__mux2_1
XFILLER_208_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13942_ _06675_ _06678_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__nor2_1
X_16730_ _09363_ _09371_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16661_ _09299_ _09300_ _09302_ vssd1 vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__a21o_1
X_13873_ _06609_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18400_ _02083_ _02098_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__xnor2_1
X_15612_ _08214_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__buf_4
XFILLER_90_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12824_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__clkbuf_4
X_19380_ rbzero.wall_tracer.rayAddendY\[-2\] _00013_ _02867_ vssd1 vssd1 vccd1 vccd1
+ _00808_ sky130_fd_sc_hd__o21a_1
X_16592_ _09231_ _09233_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__and2_1
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18331_ _01646_ _01972_ _10271_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a21o_1
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15543_ _08148_ _08183_ _08185_ _08187_ vssd1 vssd1 vccd1 vccd1 _08188_ sky130_fd_sc_hd__a31o_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12755_ _05502_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18262_ _01839_ _01847_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ rbzero.debug_overlay.facingY\[-5\] _04454_ _04463_ rbzero.debug_overlay.facingY\[-3\]
+ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a221o_1
XFILLER_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15474_ _08064_ _08118_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__xnor2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__or2_1
XFILLER_203_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14425_ _07144_ _07161_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__nand2_1
XFILLER_147_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17213_ _09791_ _09794_ vssd1 vssd1 vccd1 vccd1 _09795_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11637_ gpout0.hpos\[3\] _04023_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_1
X_18193_ _01892_ _01893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17144_ _07549_ _09763_ rbzero.row_render.size\[6\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00534_ sky130_fd_sc_hd__a2bb2o_1
X_14356_ _07090_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__nor2_1
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11568_ _04135_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13307_ _06040_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10519_ rbzero.tex_r0\[30\] rbzero.tex_r0\[29\] _03591_ vssd1 vssd1 vccd1 vccd1 _03596_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17075_ _09567_ _09569_ vssd1 vssd1 vccd1 vccd1 _09715_ sky130_fd_sc_hd__nor2_1
X_14287_ _06784_ _06796_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__or2b_1
X_11499_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _04273_ vssd1 vssd1 vccd1 vccd1 _04279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_115_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16026_ _08620_ _08670_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__nor2_1
X_13238_ _05889_ _05899_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__xnor2_4
XFILLER_100_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _05863_ _05868_ _05811_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17977_ _01555_ _01557_ _01554_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a21boi_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19716_ _03085_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16928_ _09428_ _09435_ _09568_ vssd1 vssd1 vccd1 vccd1 _09569_ sky130_fd_sc_hd__a21oi_2
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03316_ _03316_ vssd1 vssd1 vccd1 vccd1 clknet_0__03316_ sky130_fd_sc_hd__clkbuf_16
X_19647_ _03049_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__clkbuf_1
X_16859_ _09387_ _09390_ vssd1 vssd1 vccd1 vccd1 _09500_ sky130_fd_sc_hd__nand2_1
XFILLER_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18529_ _02125_ _02128_ _02225_ _05203_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a31o_1
XFILLER_33_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21540_ net461 _01309_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21471_ net392 _01240_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20422_ _09750_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__clkbuf_4
XFILLER_105_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ _03780_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__and2_1
XFILLER_197_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _05223_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and2b_1
XFILLER_185_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03305_ clknet_0__03305_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03305_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14210_ _06664_ _06940_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nand2_1
XFILLER_123_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11422_ _04175_ _04177_ _04201_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _04202_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15190_ _07820_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _07843_
+ sky130_fd_sc_hd__nand2_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ _06858_ _06876_ _06877_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a21boi_1
XFILLER_125_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11353_ rbzero.floor_leak\[3\] _04119_ _04121_ rbzero.floor_leak\[4\] _04132_ vssd1
+ vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a221o_1
X_10304_ net45 net44 vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__xor2_4
XFILLER_125_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _06806_ _06808_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__nand2_1
XFILLER_153_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11284_ _04062_ _04061_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__nand2_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13023_ _05695_ _05702_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__or2_1
X_17900_ _01472_ _01484_ _01482_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18880_ _02550_ _02551_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17831_ _01513_ _01534_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__xnor2_2
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17762_ _01464_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14974_ rbzero.wall_tracer.stepDistX\[-6\] _07650_ vssd1 vssd1 vccd1 vccd1 _07657_
+ sky130_fd_sc_hd__nor2_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19501_ _02905_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02980_
+ sky130_fd_sc_hd__or2_1
X_16713_ _08054_ _09164_ vssd1 vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__nor2_1
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _06661_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__clkbuf_2
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17693_ _10137_ _10141_ _10140_ vssd1 vssd1 vccd1 vccd1 _10258_ sky130_fd_sc_hd__a21bo_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19432_ _02899_ _02915_ _02914_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a21o_1
X_13856_ _06567_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16644_ _05194_ _09285_ _09286_ _08224_ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__a31o_1
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12807_ _05533_ _05546_ _05547_ _05284_ rbzero.wall_tracer.mapY\[8\] vssd1 vssd1
+ vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19363_ _04471_ rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02852_
+ sky130_fd_sc_hd__nand2_1
X_13787_ _06507_ _06523_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__nor2_1
XFILLER_50_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16575_ _08162_ _09217_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__nor2_1
X_10999_ rbzero.tex_b0\[58\] rbzero.tex_b0\[57\] _03843_ vssd1 vssd1 vccd1 vccd1 _03848_
+ sky130_fd_sc_hd__mux2_1
X_20143__173 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__inv_2
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18314_ _01903_ _01906_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nor2_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12738_ _05434_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__nand2_1
X_15526_ _07549_ _07552_ _07555_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__a21oi_4
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ rbzero.spi_registers.new_other\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__mux2_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15457_ _07925_ _08100_ _08101_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__a21oi_4
X_18245_ _09661_ _09359_ _01829_ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__o31a_1
XFILLER_198_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12669_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or2_1
XFILLER_204_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14408_ _06680_ _06761_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__nor2_1
XFILLER_175_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18176_ _01758_ _01760_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__nand2_1
X_15388_ _07990_ _08032_ vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__nand2_1
XFILLER_190_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14339_ _07071_ _07074_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__or2_1
X_17127_ _04154_ _04442_ vssd1 vssd1 vccd1 vccd1 _09758_ sky130_fd_sc_hd__or2_1
XFILLER_116_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17058_ _07585_ _09697_ _09431_ _09085_ vssd1 vssd1 vccd1 vccd1 _09698_ sky130_fd_sc_hd__a31o_1
X_16009_ _08622_ _08653_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__xor2_2
XFILLER_125_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20971_ clknet_leaf_53_i_clk _00740_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20226__248 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__inv_2
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21523_ net444 _01292_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21454_ net375 _01223_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21385_ net306 _01154_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 o_gpout[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 o_tex_out0 sky130_fd_sc_hd__buf_2
XFILLER_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ rbzero.tex_b1\[27\] rbzero.tex_b1\[26\] _04262_ vssd1 vssd1 vccd1 vccd1 _04746_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _06078_ _06016_ _06445_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__o31a_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ rbzero.tex_b1\[30\] rbzero.tex_b1\[31\] _03806_ vssd1 vssd1 vccd1 vccd1 _03808_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14690_ _07343_ _07344_ _07346_ _07378_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__o211ai_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _06279_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__nand2_1
XFILLER_147_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10853_ _03771_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _09003_ _09004_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__nand2_1
XFILLER_198_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13572_ _06103_ _06104_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _03735_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _07951_ _07955_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__nand2_1
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12523_ _05213_ _05232_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__o21a_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16291_ _08911_ _08934_ _08935_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__o21ba_1
XFILLER_185_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18030_ _01700_ _01731_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__xor2_1
X_15242_ _04035_ _07889_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__and2_1
X_12454_ _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ rbzero.row_render.size\[4\] _04150_ rbzero.row_render.size\[5\] vssd1 vssd1
+ vccd1 vccd1 _04185_ sky130_fd_sc_hd__o21ai_1
XFILLER_126_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15173_ _07827_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__clkbuf_1
X_12385_ _05145_ _05146_ gpout5.clk_div\[1\] _05151_ net34 vssd1 vssd1 vccd1 vccd1
+ _05152_ sky130_fd_sc_hd__a311o_2
XFILLER_153_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14124_ _06825_ _06832_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11336_ _04114_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__or2_4
XFILLER_193_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19981_ rbzero.pov.ready_buffer\[30\] _03252_ _03253_ rbzero.debug_overlay.facingY\[-1\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__o221a_1
XFILLER_67_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20173__199 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__inv_2
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14055_ _06778_ _06790_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nand2_1
X_18932_ _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__clkbuf_4
X_11267_ gpout0.vpos\[6\] _04043_ _04044_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_
+ sky130_fd_sc_hd__a211o_2
XFILLER_141_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13006_ _05700_ _05732_ _05738_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__nor3b_4
X_18863_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__or2_1
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11198_ _03972_ _03980_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__or3b_2
XFILLER_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17814_ _09434_ _09988_ _08895_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a21oi_2
X_18794_ rbzero.wall_tracer.trackDistY\[-1\] _02477_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17745_ _01445_ _01447_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__or2_1
X_14957_ rbzero.wall_tracer.visualWallDist\[10\] _07594_ vssd1 vssd1 vccd1 vccd1 _07648_
+ sky130_fd_sc_hd__or2_1
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13908_ _06574_ _06585_ _06634_ _06635_ _06636_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__a32o_1
XFILLER_165_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17676_ _10237_ _10240_ vssd1 vssd1 vccd1 vccd1 _10241_ sky130_fd_sc_hd__nand2_1
X_14888_ _07591_ _07597_ _07599_ _04039_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__o211a_1
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19415_ _02887_ _02890_ _02898_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__nand3_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16627_ _08283_ _08189_ vssd1 vssd1 vccd1 vccd1 _09270_ sky130_fd_sc_hd__nor2_1
X_13839_ _06015_ _05991_ _05978_ _06055_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__or4_1
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ _02827_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a21boi_1
X_16558_ _09082_ _09201_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15509_ _08152_ _08153_ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__or2_1
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19277_ _02793_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16489_ _07602_ _08230_ _08147_ _08236_ vssd1 vssd1 vccd1 vccd1 _09133_ sky130_fd_sc_hd__or4_1
XFILLER_164_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18228_ _01811_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18159_ _08237_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__buf_2
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21170_ clknet_leaf_79_i_clk _00939_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _04890_ _04037_ _03287_ _03911_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a31o_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ clknet_3_3_0_i_clk _00723_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20885_ clknet_leaf_82_i_clk _00654_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21506_ net427 _01275_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21437_ net358 _01206_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12170_ net42 _04918_ _04905_ _04940_ net12 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a311o_1
X_21368_ net289 _01137_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11121_ _03555_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__buf_4
XFILLER_123_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21299_ net220 _01068_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _03875_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15860_ _08492_ _08494_ _08503_ _08504_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__a31o_1
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14811_ _07459_ _07404_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__nor2_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _08406_ _08414_ _08434_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__nand3_1
X_20209__232 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__inv_2
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _10093_ _10095_ vssd1 vssd1 vccd1 vccd1 _10096_ sky130_fd_sc_hd__nand2_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20361__369 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__inv_2
X_14742_ _05807_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__buf_2
X_11954_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _04356_ vssd1 vssd1 vccd1 vccd1 _04730_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_104 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_104/HI zeros[14]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_115 vssd1 vssd1 vccd1 vccd1 ones[9] top_ew_algofoogle_115/LO sky130_fd_sc_hd__conb_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ rbzero.tex_b1\[38\] rbzero.tex_b1\[39\] _03795_ vssd1 vssd1 vccd1 vccd1 _03799_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14673_ _07409_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__inv_2
X_17461_ _09889_ _10027_ vssd1 vssd1 vccd1 vccd1 _10028_ sky130_fd_sc_hd__or2_1
X_11885_ _04140_ _04645_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__or3_1
X_19200_ _09753_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__and2_1
X_13624_ _05846_ _05975_ _06285_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__or3_1
X_16412_ _08439_ _08468_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__nor2_1
X_10836_ rbzero.tex_g0\[8\] rbzero.tex_g0\[7\] _03762_ vssd1 vssd1 vccd1 vccd1 _03763_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17392_ _08445_ _08332_ vssd1 vssd1 vccd1 vccd1 _09959_ sky130_fd_sc_hd__nand2_1
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19131_ _02700_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13555_ _05995_ _06113_ _06061_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__a21o_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16343_ _08977_ _08243_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__or2_1
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10767_ _03726_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ _05255_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.trackDistX\[0\]
+ _05257_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a22o_1
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19062_ _02663_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__clkbuf_1
X_16274_ _08915_ _08918_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__xor2_1
X_13486_ _06183_ _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__xor2_1
XFILLER_160_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10698_ rbzero.tex_g1\[8\] rbzero.tex_g1\[9\] _03680_ vssd1 vssd1 vccd1 vccd1 _03690_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18013_ _01705_ _01714_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__xor2_1
X_15225_ _07742_ _07730_ _07862_ _07821_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__a211oi_1
XFILLER_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12437_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__inv_2
X_20255__274 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__inv_2
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15156_ _07811_ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__clkbuf_1
X_12368_ _05121_ _05135_ net31 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__and3b_1
XFILLER_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ _05825_ _06668_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__nor2_1
X_11319_ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__inv_2
XFILLER_141_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15087_ _07741_ _07745_ _07746_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__a21oi_1
X_19964_ rbzero.pov.ready_buffer\[38\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-4\]
+ _03250_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__a221o_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12299_ _05044_ _05047_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__nand2_1
XFILLER_113_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14038_ _06771_ _06772_ _06773_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__o21bai_1
X_18915_ _02582_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19895_ rbzero.debug_overlay.playerY\[-8\] _03198_ _03200_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00990_ sky130_fd_sc_hd__o211a_1
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18846_ rbzero.wall_tracer.trackDistY\[6\] _02522_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02523_ sky130_fd_sc_hd__mux2_1
XFILLER_110_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18777_ rbzero.wall_tracer.trackDistY\[-3\] _02462_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02463_ sky130_fd_sc_hd__mux2_1
X_15989_ _08630_ _08631_ _08632_ _08633_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17728_ _10289_ _10291_ vssd1 vssd1 vccd1 vccd1 _10293_ sky130_fd_sc_hd__and2_1
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _10222_ _10223_ vssd1 vssd1 vccd1 vccd1 _10224_ sky130_fd_sc_hd__and2b_1
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20670_ clknet_leaf_11_i_clk _00454_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19329_ _02728_ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__or2_1
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21222_ clknet_leaf_73_i_clk _00991_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21153_ clknet_leaf_83_i_clk _00922_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21084_ net174 _00853_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20035_ _04021_ _04026_ _02705_ _04989_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a31o_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ clknet_leaf_65_i_clk _00706_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11670_ _04427_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__nor2_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20868_ clknet_leaf_59_i_clk _00637_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ rbzero.tex_g1\[45\] rbzero.tex_g1\[46\] _03647_ vssd1 vssd1 vccd1 vccd1 _03650_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20799_ clknet_leaf_18_i_clk _00568_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13340_ _06040_ _06043_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10552_ _03557_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ _05946_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__or2_1
XFILLER_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10483_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _03569_ vssd1 vssd1 vccd1 vccd1 _03577_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15010_ _07675_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__clkbuf_1
X_12222_ gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__buf_2
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ clknet_1_1__leaf__04835_ _04918_ _04905_ vssd1 vssd1 vccd1 vccd1 _04924_
+ sky130_fd_sc_hd__and3_2
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ rbzero.tex_b0\[8\] rbzero.tex_b0\[7\] _03898_ vssd1 vssd1 vccd1 vccd1 _03903_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12084_ net46 _04853_ _04854_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__a22o_1
X_16961_ _09082_ _09601_ vssd1 vssd1 vccd1 vccd1 _09602_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18700_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _09807_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__o21ai_1
X_11035_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _03865_ vssd1 vssd1 vccd1 vccd1 _03867_
+ sky130_fd_sc_hd__mux2_1
X_15912_ _08552_ _08556_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__or2b_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19680_ _03066_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16892_ _09531_ _09532_ vssd1 vssd1 vccd1 vccd1 _09533_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ _02271_ _02280_ _02278_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a21oi_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _08478_ _08485_ _08486_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__nand3_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _02257_ _02258_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _05670_ _05671_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__nand2_1
XFILLER_92_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15774_ _08417_ _08418_ vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__nand2_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17513_ _10072_ _10078_ vssd1 vssd1 vccd1 vccd1 _10079_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ rbzero.wall_tracer.stepDistY\[-12\] _07460_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07462_ sky130_fd_sc_hd__mux2_1
X_11937_ rbzero.tex_b0\[55\] _04221_ _04222_ _04218_ vssd1 vssd1 vccd1 vccd1 _04713_
+ sky130_fd_sc_hd__a31o_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _02189_ _02190_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__xor2_1
XFILLER_75_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17444_ _09972_ _10010_ vssd1 vssd1 vccd1 vccd1 _10011_ sky130_fd_sc_hd__xnor2_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14656_ _05703_ _05928_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__or2_1
X_11868_ _04371_ _04632_ _04636_ _04644_ _04244_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__o311a_1
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13607_ _06338_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__and2b_1
X_10819_ rbzero.tex_g0\[16\] rbzero.tex_g0\[15\] _03751_ vssd1 vssd1 vccd1 vccd1 _03754_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17375_ _09522_ _08705_ _08419_ vssd1 vssd1 vccd1 vccd1 _09942_ sky130_fd_sc_hd__or3_1
X_14587_ _06696_ _07072_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__and2_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11799_ rbzero.tex_g0\[46\] _04336_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__and2_1
XFILLER_186_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19114_ _02691_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16326_ _05209_ rbzero.wall_tracer.stepDistX\[3\] _08214_ vssd1 vssd1 vccd1 vccd1
+ _08971_ sky130_fd_sc_hd__a21boi_2
X_13538_ _06273_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nor2_1
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19045_ _02654_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
X_13469_ _06154_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__xnor2_1
X_16257_ _08836_ _08842_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _07742_ _07847_ _07859_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__a21o_1
X_16188_ _08828_ _08832_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ rbzero.wall_tracer.rayAddendX\[3\] _07695_ _07795_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _07796_ sky130_fd_sc_hd__a22o_1
XFILLER_142_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19947_ rbzero.pov.ready _02708_ _02820_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__nand3_4
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ rbzero.pov.ready_buffer\[72\] _03164_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_
+ sky130_fd_sc_hd__o21a_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18829_ _09863_ _02506_ _02507_ _01677_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__o31ai_1
XFILLER_110_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20722_ clknet_leaf_87_i_clk _00491_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20653_ clknet_leaf_5_i_clk _00437_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20584_ _07684_ _07690_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__and2b_1
XFILLER_192_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21205_ clknet_leaf_17_i_clk _00974_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21136_ clknet_leaf_60_i_clk _00905_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21067_ net157 _00836_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20018_ _04006_ _04811_ _04813_ _03262_ _03911_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a41o_1
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12840_ _05561_ _05468_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__or2_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ rbzero.debug_overlay.playerX\[3\] _05516_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05517_ sky130_fd_sc_hd__mux2_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _07234_ _07246_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__nor2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ rbzero.debug_overlay.playerY\[2\] _04451_ _04466_ rbzero.debug_overlay.playerY\[-8\]
+ _04500_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a221o_1
X_19573__30 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
X_15490_ _07951_ _08133_ _08134_ _05197_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__o211ai_4
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14441_ _07109_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__xnor2_1
X_11653_ _04430_ _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2b_1
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ _03640_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__clkbuf_1
X_14372_ _06240_ _06658_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__or2_1
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17160_ rbzero.traced_texa\[-9\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__a22o_1
X_11584_ _04359_ _04362_ _04332_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ _05923_ _05989_ _05983_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a21bo_1
X_16111_ _08740_ _08755_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__nand2_1
X_10535_ _03604_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17091_ _09583_ _09585_ vssd1 vssd1 vccd1 vccd1 _09731_ sky130_fd_sc_hd__nor2_1
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13254_ _05920_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16042_ _08684_ _08686_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__or2b_1
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10466_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _03558_ vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ _04960_ net16 _04972_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__and4_1
X_13185_ _05889_ _05900_ _05910_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a31o_1
XFILLER_123_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10397_ rbzero.tex_r1\[21\] rbzero.tex_r1\[22\] _03527_ vssd1 vssd1 vccd1 vccd1 _03530_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19801_ _03129_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__clkbuf_1
X_12136_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__clkbuf_4
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ _01687_ _01609_ _01693_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__and3_1
XFILLER_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19732_ rbzero.pov.spi_buffer\[40\] rbzero.pov.spi_buffer\[41\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03094_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03301_ clknet_0__03301_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03301_
+ sky130_fd_sc_hd__clkbuf_16
X_12067_ _04837_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nand2_1
X_16944_ _09382_ _09447_ _09584_ vssd1 vssd1 vccd1 vccd1 _09585_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20367__375 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__inv_2
XFILLER_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _03854_ vssd1 vssd1 vccd1 vccd1 _03858_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19663_ _03057_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20066__103 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__inv_2
X_16875_ _09514_ _09515_ vssd1 vssd1 vccd1 vccd1 _09516_ sky130_fd_sc_hd__nand2_1
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18614_ _02307_ _02309_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__and2_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _08024_ _08014_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__nand2_1
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18545_ _10248_ _10266_ _02151_ _02045_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__o31a_1
X_15757_ _08064_ _08118_ _08401_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__a21o_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _05563_ _05566_ _05591_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__and3_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _05779_ _07428_ _07429_ _05742_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__o211a_1
X_18476_ _10239_ _09215_ _02173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__or3_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ _08129_ _08104_ _08331_ _08332_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17427_ _09987_ _09993_ vssd1 vssd1 vccd1 vccd1 _09994_ sky130_fd_sc_hd__xor2_2
X_14639_ _05742_ _05755_ _07105_ _07374_ _07375_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__a32o_1
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17358_ _08416_ _09704_ vssd1 vssd1 vccd1 vccd1 _09925_ sky130_fd_sc_hd__nor2_1
X_16309_ _08619_ _08950_ _08946_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__and3b_1
XFILLER_146_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ rbzero.wall_tracer.trackDistX\[-6\] _09861_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09862_ sky130_fd_sc_hd__mux2_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19028_ _02645_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20705_ clknet_leaf_0_i_clk _00489_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03321_ clknet_0__03321_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03321_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20636_ clknet_leaf_27_i_clk _00420_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20567_ rbzero.traced_texVinit\[10\] _03443_ _09771_ _10297_ vssd1 vssd1 vccd1 vccd1
+ _01418_ sky130_fd_sc_hd__a22o_1
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10320_ _03489_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20498_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03396_
+ sky130_fd_sc_hd__nand2_1
XFILLER_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21119_ net209 _00888_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[59\] sky130_fd_sc_hd__dfxtp_1
X_19625__78 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__inv_2
XFILLER_94_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14990_ _07665_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__clkbuf_1
X_13941_ _06677_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16660_ _09299_ _09300_ _09302_ vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__nand3_2
X_13872_ _06548_ _06608_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__or2_1
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ _08253_ _08255_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__xnor2_2
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12823_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__clkinv_2
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16591_ _09231_ _09233_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__nor2_1
XFILLER_55_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18330_ _01646_ _02028_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _07951_ _08186_ _05207_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__a21o_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ rbzero.map_rom.f3 _05501_ _05414_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__mux2_1
XFILLER_188_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18261_ _01846_ _01840_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__and2b_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ rbzero.debug_overlay.facingY\[0\] _04459_ _04460_ rbzero.debug_overlay.facingY\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a22o_1
X_15473_ _08108_ _08117_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__xor2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _05431_ _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and2_2
XFILLER_188_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17212_ _09792_ _09793_ vssd1 vssd1 vccd1 vccd1 _09794_ sky130_fd_sc_hd__or2_1
X_14424_ _07133_ _07143_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__nand2_1
X_11636_ gpout0.hpos\[9\] _04414_ _04046_ _04020_ vssd1 vssd1 vccd1 vccd1 _04415_
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18192_ _01890_ _01891_ _01855_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a21o_1
X_17143_ _09765_ _09763_ rbzero.row_render.size\[5\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00533_ sky130_fd_sc_hd__a2bb2o_1
X_14355_ _06735_ _07030_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__a21oi_1
X_11567_ _04343_ _04344_ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13306_ _05943_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__and2_1
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10518_ _03595_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
X_14286_ _07015_ _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__xnor2_2
XFILLER_155_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17074_ _09702_ _09713_ vssd1 vssd1 vccd1 vccd1 _09714_ sky130_fd_sc_hd__xnor2_2
X_11498_ rbzero.tex_r0\[15\] _04221_ _04222_ _04219_ vssd1 vssd1 vccd1 vccd1 _04278_
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__buf_2
X_16025_ _08666_ _08668_ _08669_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__o21a_1
X_10449_ _03559_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13168_ _05902_ _05874_ _05904_ _05755_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__o22a_1
XFILLER_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12119_ gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__buf_2
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13099_ _05640_ _05648_ _05791_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__mux2_1
X_17976_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__and2_1
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19715_ rbzero.pov.spi_buffer\[32\] rbzero.pov.spi_buffer\[33\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_62_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16927_ _08215_ _09294_ _09427_ vssd1 vssd1 vccd1 vccd1 _09568_ sky130_fd_sc_hd__nor3_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03315_ _03315_ vssd1 vssd1 vccd1 vccd1 clknet_0__03315_ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19646_ rbzero.pov.mosi rbzero.pov.spi_buffer\[0\] _03048_ vssd1 vssd1 vccd1 vccd1
+ _03049_ sky130_fd_sc_hd__mux2_1
X_16858_ _09366_ _09369_ _09365_ vssd1 vssd1 vccd1 vccd1 _09499_ sky130_fd_sc_hd__a21bo_1
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20395__20 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15809_ _08444_ _08450_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__nor2_1
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16789_ _07575_ _08983_ _09430_ vssd1 vssd1 vccd1 vccd1 _09431_ sky130_fd_sc_hd__nor3_2
XFILLER_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_77_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18528_ _02125_ _02128_ _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18459_ _02155_ _02156_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__nor2_1
XFILLER_166_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20120__152 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__inv_2
X_21470_ net391 _01239_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20421_ _03272_ _03330_ _03331_ _03327_ rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1
+ _01385_ sky130_fd_sc_hd__a32o_1
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_175_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20283_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__buf_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20203__227 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__inv_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ rbzero.wall_tracer.trackDistY\[5\] _05222_ _05224_ rbzero.wall_tracer.trackDistY\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__o22ai_1
XFILLER_71_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21668_ clknet_leaf_47_i_clk _01437_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03304_ clknet_0__03304_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03304_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _04154_ _04179_ _04180_ _04181_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__o221a_1
X_20619_ clknet_leaf_72_i_clk _00403_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.b6 sky130_fd_sc_hd__dfxtp_1
XFILLER_165_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21599_ net140 _01368_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14140_ _06859_ _06875_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__or2b_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11352_ rbzero.floor_leak\[2\] _04123_ _04119_ rbzero.floor_leak\[3\] _04131_ vssd1
+ vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__o221a_1
XFILLER_193_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10303_ _03476_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__and2_1
X_14071_ _06776_ _06739_ _06804_ _06807_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__o31a_1
X_11283_ rbzero.texV\[6\] _04061_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__a21boi_1
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022_ _05756_ _05758_ _05737_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17830_ _01532_ _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__and2b_1
XFILLER_126_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17761_ _09391_ _09359_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__nor2_1
XFILLER_94_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14973_ _00008_ _07524_ _07656_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19500_ _02952_ _02976_ _02977_ _02975_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a31o_1
XFILLER_208_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16712_ _08331_ _09353_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__nand2_1
X_13924_ _06613_ _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__or2_1
X_17692_ _09974_ _10255_ _10256_ _10117_ vssd1 vssd1 vccd1 vccd1 _10257_ sky130_fd_sc_hd__a22o_1
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19431_ _02890_ _02898_ _02885_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a21bo_1
X_16643_ _07575_ _07579_ _08983_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__or3_1
X_13855_ _06589_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__xor2_1
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19362_ _04471_ rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02851_
+ sky130_fd_sc_hd__nor2_1
X_12806_ _05539_ _05541_ _05545_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__o21ai_1
X_16574_ _09216_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13786_ _06509_ _06519_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__a21o_1
X_10998_ _03847_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18313_ _02011_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__or2b_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _07981_ vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__clkbuf_4
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__nand2_1
X_19293_ _02802_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__clkbuf_1
X_20178__204 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__inv_2
XFILLER_188_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _01827_ _01828_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__nand2_1
XFILLER_176_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15456_ _07904_ rbzero.wall_tracer.stepDistY\[-8\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _08101_ sky130_fd_sc_hd__a21o_1
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12668_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nand2_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14407_ _07133_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__or2_1
XFILLER_204_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11619_ rbzero.tex_r1\[47\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04398_
+ sky130_fd_sc_hd__a31o_1
X_18175_ _01857_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__xnor2_1
X_15387_ rbzero.wall_tracer.visualWallDist\[0\] _08031_ _07904_ vssd1 vssd1 vccd1
+ vccd1 _08032_ sky130_fd_sc_hd__mux2_1
X_12599_ _05352_ _05291_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__xnor2_2
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17126_ _09757_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__clkbuf_1
X_14338_ _07071_ _07074_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__nand2_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17057_ _07589_ vssd1 vssd1 vccd1 vccd1 _09697_ sky130_fd_sc_hd__inv_2
X_14269_ _07005_ _06732_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__xnor2_2
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16008_ _08638_ _08651_ _08652_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__a21oi_2
XFILLER_48_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _01454_ _01542_ _01661_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a21oi_1
XFILLER_211_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20970_ clknet_leaf_52_i_clk _00739_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.vinf
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21522_ net443 _01291_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21453_ net374 _01222_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21384_ net305 _01153_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 o_hsync sky130_fd_sc_hd__buf_2
XFILLER_0_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _04741_ _04744_ _04332_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__mux2_1
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10921_ _03807_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13640_ _06336_ _06375_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__nor3_1
X_10852_ rbzero.tex_b1\[63\] net48 _03691_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _06306_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _03729_ vssd1 vssd1 vccd1 vccd1 _03735_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _07954_ rbzero.debug_overlay.playerY\[-4\] _05374_ vssd1 vssd1 vccd1 vccd1
+ _07955_ sky130_fd_sc_hd__mux2_1
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12522_ _05235_ _05276_ _05228_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or3b_1
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _08849_ _08845_ _08847_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__and3_1
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ rbzero.wall_tracer.wall\[0\] _03999_ _05280_ _03987_ vssd1 vssd1 vccd1 vccd1
+ _07889_ sky130_fd_sc_hd__a22o_1
XFILLER_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12453_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__clkbuf_4
X_11404_ _04152_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__nor2_1
XFILLER_201_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12384_ net123 _05145_ _05146_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a21oi_2
XFILLER_153_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ rbzero.wall_tracer.rayAddendX\[5\] _07826_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07827_ sky130_fd_sc_hd__mux2_1
XFILLER_126_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14123_ _06851_ _06853_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11335_ _04101_ _04105_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19980_ rbzero.pov.ready_buffer\[29\] _03247_ _03249_ rbzero.debug_overlay.facingY\[-2\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__a221o_1
XFILLER_180_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18931_ _02593_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__clkbuf_4
XFILLER_107_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14054_ _06778_ _06790_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__xnor2_1
X_11266_ gpout0.hpos\[7\] gpout0.hpos\[8\] _04045_ gpout0.hpos\[9\] vssd1 vssd1 vccd1
+ vccd1 _04046_ sky130_fd_sc_hd__a31oi_2
X_13005_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__clkbuf_4
X_18862_ _02536_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
X_11197_ rbzero.map_rom.d6 _03942_ _03981_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_
+ sky130_fd_sc_hd__o31a_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17813_ _10130_ _10266_ _10265_ _10267_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18793_ _05204_ _02475_ _02476_ _09897_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a31o_1
XFILLER_208_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17744_ _01445_ _01447_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__nand2_1
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14956_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.trackDistX\[10\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13907_ _06637_ _06619_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__and2b_1
X_20062__99 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__inv_2
X_17675_ _09126_ _08493_ _10238_ _10239_ vssd1 vssd1 vccd1 vccd1 _10240_ sky130_fd_sc_hd__o22ai_1
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _07598_ _04019_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__nand2_1
XFILLER_165_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19414_ _02887_ _02890_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a21o_1
X_16626_ _09128_ _09130_ _09131_ _09127_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__a22o_1
X_13838_ _06258_ _06261_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__and2b_1
XFILLER_51_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19345_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nand2_1
X_16557_ _09199_ _09200_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13769_ _06486_ _06487_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__or2_1
XFILLER_188_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15508_ _08131_ _08136_ _08127_ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19276_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_leak\[0\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XFILLER_203_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16488_ _09127_ _09131_ vssd1 vssd1 vccd1 vccd1 _09132_ sky130_fd_sc_hd__xor2_2
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18227_ _01925_ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__nor2_1
XFILLER_176_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15439_ _05207_ _08079_ _08082_ _08083_ vssd1 vssd1 vccd1 vccd1 _08084_ sky130_fd_sc_hd__a22o_4
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18158_ _08237_ _08493_ _08044_ _09973_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or4_1
XFILLER_141_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17109_ _09747_ vssd1 vssd1 vccd1 vccd1 _09748_ sky130_fd_sc_hd__buf_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18089_ _01667_ _01676_ _01789_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a21oi_1
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20232__253 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__inv_2
XFILLER_113_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20051_ _04990_ _04989_ _04322_ _02705_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a41o_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ clknet_leaf_49_i_clk _00722_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ clknet_leaf_82_i_clk _00653_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21505_ net426 _01274_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21436_ net357 _01205_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[15\] sky130_fd_sc_hd__dfxtp_1
X_20315__328 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__inv_2
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21367_ net288 _01136_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11120_ rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkinv_8
XFILLER_123_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21298_ net219 _01067_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11051_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _03865_ vssd1 vssd1 vccd1 vccd1 _03875_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20249_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__buf_1
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _05884_ _05952_ _07469_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__a31o_1
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _08406_ _08414_ _08434_ vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__a21o_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _07107_ _07350_ _07379_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__a21boi_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _04356_ vssd1 vssd1 vccd1 vccd1 _04729_
+ sky130_fd_sc_hd__mux2_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_105 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_105/HI zeros[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_116 vssd1 vssd1 vccd1 vccd1 ones[10] top_ew_algofoogle_116/LO sky130_fd_sc_hd__conb_1
XFILLER_205_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _03798_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17460_ _09906_ _10026_ vssd1 vssd1 vccd1 vccd1 _10027_ sky130_fd_sc_hd__xor2_4
X_14672_ _07342_ _07408_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__nand2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ _04241_ _04652_ _04660_ _04143_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__o211a_1
XFILLER_205_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16411_ _09053_ _09055_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__xnor2_2
X_13623_ _06355_ _06359_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__xor2_1
XFILLER_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10835_ _03717_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17391_ _09682_ _09690_ _09689_ vssd1 vssd1 vccd1 vccd1 _09958_ sky130_fd_sc_hd__a21o_1
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19130_ net43 rbzero.spi_registers.sclk_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02700_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16342_ _08979_ _08986_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__xnor2_2
X_13554_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__xnor2_2
XFILLER_185_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _03718_ vssd1 vssd1 vccd1 vccd1 _03726_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19061_ rbzero.pov.spi_buffer\[61\] rbzero.pov.ready_buffer\[61\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
X_12505_ _05253_ _05256_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__nand3_1
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16273_ _08816_ _08335_ _08916_ _08917_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__o31ai_2
X_13485_ _06211_ _06221_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ _03689_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18012_ _01712_ _01713_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__nor2_1
XFILLER_173_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _07873_ _07874_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__and2_1
XFILLER_126_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12436_ rbzero.wall_tracer.state\[6\] vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15155_ rbzero.wall_tracer.rayAddendX\[4\] _07810_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07811_ sky130_fd_sc_hd__mux2_1
X_12367_ _05131_ _05132_ _05133_ _05134_ net28 _05082_ vssd1 vssd1 vccd1 vccd1 _05135_
+ sky130_fd_sc_hd__mux4_1
XFILLER_154_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14106_ _06704_ _06760_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__nor2_1
XFILLER_181_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _04060_ _04063_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12298_ clknet_1_0__leaf__04835_ _05046_ _05047_ vssd1 vssd1 vccd1 vccd1 _05067_
+ sky130_fd_sc_hd__and3_2
X_15086_ _07741_ _07745_ _04034_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__o21ai_1
X_19963_ rbzero.pov.ready_buffer\[37\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-5\]
+ _03250_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__a221o_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14037_ _06771_ _06772_ _06773_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__or3b_1
X_18914_ _02580_ _02581_ _02574_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__and3b_1
X_11249_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__buf_2
XFILLER_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19894_ _07982_ _02823_ _03198_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o211ai_1
XFILLER_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18845_ _02520_ _02521_ _01908_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a21bo_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18776_ _09863_ _02460_ _02461_ _09885_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__o31ai_1
X_15988_ _08008_ _08022_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__nor2_1
XFILLER_209_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17727_ _10289_ _10291_ vssd1 vssd1 vccd1 vccd1 _10292_ sky130_fd_sc_hd__nor2_1
X_14939_ _07621_ _07634_ _07635_ _07620_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__o211a_1
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ _10216_ _10221_ vssd1 vssd1 vccd1 vccd1 _10223_ sky130_fd_sc_hd__or2_1
XFILLER_36_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16609_ _08282_ _08383_ _08111_ _08570_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__or4_1
XFILLER_189_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17589_ _10152_ _10154_ vssd1 vssd1 vccd1 vccd1 _10155_ sky130_fd_sc_hd__xor2_1
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19328_ net39 net38 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__nor2_4
XFILLER_189_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19259_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21221_ clknet_leaf_17_i_clk _00990_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_144_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21152_ clknet_leaf_83_i_clk _00921_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21083_ net173 _00852_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20034_ _04989_ _04037_ _02705_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and3_1
XFILLER_113_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ clknet_leaf_65_i_clk _00705_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ clknet_leaf_59_i_clk _00636_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10620_ _03649_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20798_ clknet_leaf_18_i_clk _00567_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10551_ _03612_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20239__259 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__inv_2
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10482_ _03576_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
X_13270_ _05852_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and3_1
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ _04989_ _04990_ _04961_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__mux2_1
X_21419_ net340 _01188_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12152_ gpout1.clk_div\[1\] _04922_ _04905_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__and3_1
XFILLER_123_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11103_ _03902_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12083_ net3 net2 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and2_2
X_16960_ _09599_ _09600_ vssd1 vssd1 vccd1 vccd1 _09601_ sky130_fd_sc_hd__nor2_1
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11034_ _03866_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__clkbuf_1
X_15911_ _08475_ _08553_ _08554_ _08555_ vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__a2bb2o_1
X_16891_ _08383_ _09103_ vssd1 vssd1 vccd1 vccd1 _09532_ sky130_fd_sc_hd__or2_1
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18630_ _02268_ _02284_ _02282_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a21o_1
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _08478_ _08485_ _08486_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__a21o_1
XFILLER_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _08445_ _09704_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__nor2_1
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _05208_ _08149_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__nor2_4
X_12985_ _05705_ _05708_ _05719_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a211oi_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17512_ _10076_ _10077_ vssd1 vssd1 vccd1 vccd1 _10078_ sky130_fd_sc_hd__xor2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _05188_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__buf_4
X_11936_ rbzero.tex_b0\[54\] _04338_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__and2_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _01739_ _08423_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__nor2_1
XFILLER_73_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17443_ _10007_ _10009_ vssd1 vssd1 vccd1 vccd1 _10010_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14655_ _05742_ _05755_ _07377_ _07391_ _07375_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__a32o_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _04209_ _04639_ _04643_ _04142_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a211o_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _06295_ _06339_ _06340_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__a22o_1
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10818_ _03753_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17374_ _08705_ _08159_ _08151_ _09522_ vssd1 vssd1 vccd1 vccd1 _09941_ sky130_fd_sc_hd__o22a_1
X_14586_ _07284_ _07321_ _07322_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__a21o_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11798_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _04341_ vssd1 vssd1 vccd1 vccd1 _04576_
+ sky130_fd_sc_hd__mux2_1
X_19113_ net512 rbzero.spi_registers.spi_cmd\[0\] _02690_ vssd1 vssd1 vccd1 vccd1
+ _02691_ sky130_fd_sc_hd__mux2_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16325_ _08968_ _08969_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__and2_1
X_13537_ _06225_ _06233_ _06272_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__and3_1
XFILLER_186_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10749_ _03716_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19044_ rbzero.pov.spi_buffer\[53\] rbzero.pov.ready_buffer\[53\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XFILLER_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16256_ _08885_ _08888_ _08900_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__a21oi_1
X_13468_ _06201_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__xor2_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _07857_ _07858_ _07847_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12419_ net35 _05180_ _05182_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__o211a_1
XFILLER_145_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16187_ _08829_ _08831_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__and2b_1
X_13399_ _06132_ _06133_ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__o21ba_1
XFILLER_114_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15138_ _07775_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15069_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__clkbuf_4
X_19946_ _03236_ _03238_ _02714_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__o21a_1
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19877_ _02820_ _03185_ _03155_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__o21a_1
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18828_ _02503_ _02504_ _02505_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__o21a_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20344__354 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__inv_2
X_18759_ _02443_ _02444_ _02445_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a21oi_1
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20721_ clknet_leaf_22_i_clk _00014_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20652_ clknet_leaf_5_i_clk _00436_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20583_ rbzero.wall_tracer.rayAddendX\[-8\] _03443_ _03452_ _03453_ vssd1 vssd1 vccd1
+ vccd1 _01425_ sky130_fd_sc_hd__a22o_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21204_ clknet_leaf_53_i_clk _00973_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21135_ clknet_leaf_62_i_clk _00904_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21066_ net156 _00835_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20017_ _04006_ _04811_ _04813_ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__or4bb_1
XFILLER_150_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _05514_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ rbzero.debug_overlay.playerY\[1\] _04449_ _04499_ rbzero.debug_overlay.playerY\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__a22o_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ clknet_leaf_70_i_clk _00688_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _06680_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__and3b_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11652_ _04423_ _04426_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and2_1
XFILLER_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ rbzero.tex_g1\[53\] rbzero.tex_g1\[54\] _03635_ vssd1 vssd1 vccd1 vccd1 _03640_
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14371_ _06680_ _07072_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__or2_2
XFILLER_126_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11583_ _04360_ _04361_ _04345_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__mux2_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16110_ _08741_ _08753_ _08754_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__a21oi_1
X_13322_ _05923_ _06054_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nand2_1
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10534_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _03602_ vssd1 vssd1 vccd1 vccd1 _03604_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17090_ _09616_ _09729_ vssd1 vssd1 vccd1 vccd1 _09730_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16041_ _08623_ _08685_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__xnor2_1
X_10465_ _03567_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_1
X_13253_ _05909_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__buf_2
XFILLER_196_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12204_ _04966_ net66 _04973_ net18 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a211o_1
X_13184_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__clkinv_2
X_10396_ _03529_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19800_ _04867_ rbzero.pov.mosi_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1 _03129_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12135_ net9 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__inv_2
XFILLER_69_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17992_ _01687_ _01609_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03300_ clknet_0__03300_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03300_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19731_ _03093_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
X_16943_ _09445_ _09446_ vssd1 vssd1 vccd1 vccd1 _09584_ sky130_fd_sc_hd__nor2_1
X_12066_ net3 net2 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__nor2_2
X_11017_ _03857_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__clkbuf_1
X_19662_ rbzero.pov.spi_buffer\[7\] rbzero.pov.spi_buffer\[8\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
X_16874_ _09478_ _09479_ _09513_ vssd1 vssd1 vccd1 vccd1 _09515_ sky130_fd_sc_hd__nand3_1
XFILLER_133_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15825_ _08169_ _08469_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__xnor2_1
X_18613_ _02307_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__nor2_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__buf_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15756_ _08108_ _08117_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__nor2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _02239_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _05589_ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__xnor2_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _07375_ _07440_ _07441_ _07443_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__a31o_1
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11919_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _04271_ vssd1 vssd1 vccd1 vccd1 _04695_
+ sky130_fd_sc_hd__mux2_1
X_18475_ _02071_ _02172_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15687_ _05210_ _08044_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__nor2_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _05622_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__xor2_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17426_ _08266_ _09696_ _09989_ _09992_ vssd1 vssd1 vccd1 vccd1 _09993_ sky130_fd_sc_hd__a31oi_2
X_14638_ _05932_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__buf_2
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17357_ _09922_ _09923_ vssd1 vssd1 vccd1 vccd1 _09924_ sky130_fd_sc_hd__nand2_1
XFILLER_202_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14569_ _07305_ _07093_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__nand2_1
XFILLER_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _08619_ _08952_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__xnor2_4
XFILLER_140_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17288_ _09812_ _09857_ _09858_ _09860_ vssd1 vssd1 vccd1 vccd1 _09861_ sky130_fd_sc_hd__o31ai_1
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19027_ rbzero.pov.spi_buffer\[45\] rbzero.pov.ready_buffer\[45\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
X_16239_ _08879_ _08883_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19929_ _03223_ _03224_ _02822_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20704_ clknet_leaf_92_i_clk _00488_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__03320_ clknet_0__03320_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03320_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20635_ clknet_leaf_8_i_clk _00419_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20566_ rbzero.traced_texVinit\[9\] _09764_ _07831_ _10171_ vssd1 vssd1 vccd1 vccd1
+ _01417_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_164_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20497_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03395_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21118_ net208 _00887_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13940_ _06612_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__nor2_2
X_21049_ clknet_leaf_2_i_clk _00818_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _06547_ _06497_ _06498_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__and3_1
XFILLER_90_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15610_ _07601_ _04015_ _05198_ _08254_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__and4_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12822_ rbzero.wall_tracer.mapY\[11\] _05284_ _05533_ _05559_ vssd1 vssd1 vccd1 vccd1
+ _00418_ sky130_fd_sc_hd__a22o_1
XFILLER_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16590_ _09167_ _09174_ _09232_ vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__a21oi_1
XFILLER_131_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15541_ rbzero.wall_tracer.stepDistY\[2\] vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__inv_2
X_12753_ _05204_ _05498_ _05499_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a31o_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18260_ _01952_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__xnor2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11704_ rbzero.debug_overlay.facingY\[-4\] _04464_ _04465_ rbzero.debug_overlay.facingY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a22o_1
XFILLER_203_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15472_ _08115_ _08116_ _08110_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__o21a_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12684_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__or2_1
XFILLER_187_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ rbzero.wall_tracer.mapX\[9\] _05525_ vssd1 vssd1 vccd1 vccd1 _09793_ sky130_fd_sc_hd__nor2_1
X_14423_ _07158_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__or2_1
XFILLER_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ gpout0.hpos\[6\] _04008_ _04023_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__and3_1
X_18191_ _01855_ _01890_ _01891_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__nand3_1
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17142_ _07468_ _07544_ vssd1 vssd1 vccd1 vccd1 _09765_ sky130_fd_sc_hd__nor2_1
X_14354_ _07027_ _07029_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__nor2_1
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _04224_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__buf_6
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _06041_ _05940_ _05942_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__o21ai_1
X_20373__380 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__inv_2
XFILLER_171_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10517_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _03591_ vssd1 vssd1 vccd1 vccd1 _03595_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17073_ _09709_ _09712_ vssd1 vssd1 vccd1 vccd1 _09713_ sky130_fd_sc_hd__xor2_2
X_14285_ _07020_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__xor2_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11497_ rbzero.tex_r0\[14\] _04214_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__and2_1
XFILLER_137_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16024_ _08621_ _08665_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__or2_1
XFILLER_100_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _05969_ _05972_ _05871_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__mux2_2
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10448_ net46 rbzero.tex_r0\[63\] _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__mux2_1
XFILLER_136_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _05890_ _05903_ _05826_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__mux2_1
XFILLER_124_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10379_ _03520_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__buf_2
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13098_ _05740_ _05828_ _05832_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__o211a_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17975_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__nor2_1
X_19714_ _03084_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12049_ rbzero.row_render.texu\[2\] _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16926_ _09562_ _09566_ vssd1 vssd1 vccd1 vccd1 _09567_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_0__03314_ _03314_ vssd1 vssd1 vccd1 vccd1 clknet_0__03314_ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19645_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16857_ _09487_ _09497_ vssd1 vssd1 vccd1 vccd1 _09498_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _08452_ _08009_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__xnor2_2
X_16788_ _07579_ _07582_ vssd1 vssd1 vccd1 vccd1 _09430_ sky130_fd_sc_hd__or2_1
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18527_ _02222_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__nand2_1
X_15739_ _08383_ _07981_ _08180_ _08282_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__o22ai_1
XFILLER_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18458_ _02153_ _02154_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__and2_1
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ _09288_ _09695_ vssd1 vssd1 vccd1 vccd1 _09976_ sky130_fd_sc_hd__and2_1
XFILLER_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18389_ _01739_ _01475_ _01476_ _01860_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__o22ai_1
XFILLER_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20420_ _03328_ _03329_ _03325_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19630__82 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__inv_2
XFILLER_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21667_ clknet_leaf_47_i_clk _01436_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03303_ clknet_0__03303_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03303_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ _03475_ _04182_ _04179_ _04154_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__a221o_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20618_ clknet_leaf_72_i_clk _00402_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.c6 sky130_fd_sc_hd__dfxtp_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21598_ net139 _01367_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ rbzero.floor_leak\[2\] _04123_ _04126_ rbzero.floor_leak\[1\] _04130_ vssd1
+ vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a221o_1
XFILLER_180_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20549_ _03430_ _03435_ _03436_ _03437_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand4_1
XFILLER_152_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__buf_2
XFILLER_125_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14070_ _06769_ _06615_ _06738_ _06707_ _06776_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__o32ai_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11282_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _04062_ sky130_fd_sc_hd__nand2_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _05710_ _05713_ _05757_ _05687_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__or4_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14972_ rbzero.wall_tracer.stepDistX\[-7\] _00008_ vssd1 vssd1 vccd1 vccd1 _07656_
+ sky130_fd_sc_hd__nor2_1
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17760_ _01462_ _10205_ _01463_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__o21ba_1
XFILLER_102_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13923_ _06603_ _06612_ _06560_ _06601_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__o211a_1
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16711_ _09028_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__inv_2
X_17691_ _09980_ _10115_ vssd1 vssd1 vccd1 vccd1 _10256_ sky130_fd_sc_hd__or2_1
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19430_ _02912_ _02913_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__nand2_1
X_16642_ _07575_ _08983_ _07579_ vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__o21ai_1
X_13854_ _06255_ _06265_ _06590_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ _05539_ _05541_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__or3_1
X_19361_ rbzero.debug_overlay.vplaneY\[-7\] _02847_ vssd1 vssd1 vccd1 vccd1 _02850_
+ sky130_fd_sc_hd__nand2_1
X_16573_ _05210_ _09215_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__or2_1
X_13785_ _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__and2_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10997_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _03843_ vssd1 vssd1 vccd1 vccd1 _03847_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15524_ _08120_ _08146_ _08168_ vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__a21oi_2
XFILLER_31_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18312_ _01915_ _01916_ _02010_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a21o_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ rbzero.spi_registers.new_other\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__mux2_1
X_12736_ _05461_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nor2_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _01941_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__xnor2_1
X_15455_ _07933_ _07514_ _08099_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__o21ai_1
XFILLER_203_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12667_ _05415_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ _07134_ _07135_ _07142_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__a21oi_1
XFILLER_198_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ rbzero.tex_r1\[46\] _04272_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and2_1
X_18174_ _01858_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__xor2_1
X_15386_ _05374_ _08030_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__nor2_1
XFILLER_184_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12598_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17125_ _04443_ _09750_ vssd1 vssd1 vccd1 vccd1 _09757_ sky130_fd_sc_hd__and2_1
X_14337_ _06017_ _07073_ _06770_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11549_ _04136_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__buf_4
XFILLER_184_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ _09292_ _09695_ _08872_ vssd1 vssd1 vccd1 vccd1 _09696_ sky130_fd_sc_hd__a21oi_2
X_14268_ _07003_ _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__xnor2_2
X_16007_ _08639_ _08650_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__nor2_1
X_13219_ _05740_ _05828_ _05932_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14199_ _06776_ _06610_ _06671_ _06769_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__o22a_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20150__179 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__inv_2
XFILLER_111_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _01539_ _01541_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16909_ _09539_ _09549_ vssd1 vssd1 vccd1 vccd1 _09550_ sky130_fd_sc_hd__xor2_2
X_17889_ _01478_ _01480_ _01477_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a21bo_1
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19559_ rbzero.pov.spi_counter\[3\] _03028_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nand2_1
XFILLER_179_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21521_ net442 _01290_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21452_ net373 _01221_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21383_ net304 _01152_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ rbzero.tex_b1\[31\] rbzero.tex_b1\[32\] _03806_ vssd1 vssd1 vccd1 vccd1 _03807_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _03770_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13570_ _06107_ _06106_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__and2b_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _03734_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _05250_ _05260_ _05271_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o31a_1
XFILLER_73_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ rbzero.wall_tracer.rayAddendX\[11\] _07855_ _07679_ _07888_ _07880_ vssd1
+ vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a221o_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12452_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__buf_4
XFILLER_173_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ rbzero.row_render.size\[6\] _04151_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__nor2_1
XFILLER_123_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15171_ _07814_ _07815_ _04033_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__a2bb2o_1
X_12383_ net50 _05142_ _05148_ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a211o_1
XFILLER_201_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ _06822_ _06835_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11334_ rbzero.row_render.vinf _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__nor2_8
XFILLER_67_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14053_ _06776_ _06739_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__nor2_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18930_ rbzero.pov.spi_done _03480_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__nand2_1
X_11265_ _04008_ _04023_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_76_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _05740_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__buf_2
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18861_ rbzero.wall_tracer.trackDistY\[8\] _02535_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02536_ sky130_fd_sc_hd__mux2_1
XFILLER_79_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11196_ rbzero.map_rom.f3 _03942_ _03976_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_
+ sky130_fd_sc_hd__a211o_1
X_17812_ _10110_ _09973_ _10260_ _01515_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o31ai_2
X_18792_ _02474_ _02469_ _02472_ _02473_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a211o_1
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17743_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
X_14955_ _04019_ _07645_ _07646_ _07642_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__o211a_1
XFILLER_94_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ _06640_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__inv_2
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17674_ _08259_ vssd1 vssd1 vccd1 vccd1 _10239_ sky130_fd_sc_hd__clkbuf_4
X_14886_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1 vccd1 vccd1 _07598_
+ sky130_fd_sc_hd__inv_2
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19413_ _04471_ rbzero.debug_overlay.vplaneY\[-7\] vssd1 vssd1 vccd1 vccd1 _02898_
+ sky130_fd_sc_hd__xnor2_1
X_13837_ _06572_ _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__and2_1
X_16625_ _08963_ _09119_ _09267_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__a21bo_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_165_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _09065_ _09077_ _09078_ _09064_ vssd1 vssd1 vccd1 vccd1 _09200_ sky130_fd_sc_hd__a31o_1
X_19344_ _02828_ _02833_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13768_ _05825_ _06240_ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__or3_1
XFILLER_210_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12719_ _05430_ _05433_ _05431_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a21boi_1
X_15507_ _08135_ _08151_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__or2_2
XFILLER_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19275_ _02791_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__buf_2
X_16487_ _09128_ _09130_ vssd1 vssd1 vccd1 vccd1 _09131_ sky130_fd_sc_hd__xor2_2
XFILLER_188_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13699_ _06428_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__or2_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18226_ _01918_ _01919_ _01924_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__and3_1
X_15438_ rbzero.wall_tracer.visualWallDist\[-2\] _07925_ _05206_ vssd1 vssd1 vccd1
+ vccd1 _08083_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_29_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15369_ _07913_ _07941_ _07967_ _07924_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__o22ai_1
X_18157_ _01755_ _01763_ _01762_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a21bo_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17108_ _03555_ _04037_ vssd1 vssd1 vccd1 vccd1 _09747_ sky130_fd_sc_hd__or2_1
X_18088_ _01667_ _01676_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__and3_1
XFILLER_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17039_ _09660_ _09678_ vssd1 vssd1 vccd1 vccd1 _09679_ sky130_fd_sc_hd__xor2_2
XFILLER_131_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20050_ _03266_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__inv_2
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ clknet_leaf_59_i_clk _00721_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ clknet_leaf_61_i_clk _00652_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21504_ net425 _01273_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21435_ net356 _01204_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21366_ net287 _01135_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21297_ net218 _01066_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[4\] sky130_fd_sc_hd__dfxtp_1
X_11050_ _03874_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _07107_ _07356_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__a21oi_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11952_ _04218_ _04727_ _04253_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__o21a_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_106 vssd1 vssd1 vccd1 vccd1 ones[0] top_ew_algofoogle_106/LO sky130_fd_sc_hd__conb_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_117 vssd1 vssd1 vccd1 vccd1 ones[11] top_ew_algofoogle_117/LO sky130_fd_sc_hd__conb_1
XFILLER_205_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ rbzero.tex_b1\[39\] rbzero.tex_b1\[40\] _03795_ vssd1 vssd1 vccd1 vccd1 _03798_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14671_ _07213_ _07328_ _07332_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__a21o_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _04229_ _04655_ _04659_ _04119_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a211o_1
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _08413_ _09054_ _08435_ vssd1 vssd1 vccd1 vccd1 _09055_ sky130_fd_sc_hd__o21a_1
X_13622_ _06313_ _06356_ _06357_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__o22a_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10834_ _03761_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17390_ _09665_ _09666_ _09677_ _09956_ vssd1 vssd1 vccd1 vccd1 _09957_ sky130_fd_sc_hd__a31o_1
XFILLER_201_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16341_ _08239_ _08985_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__nor2_1
X_13553_ _06112_ _06118_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__xor2_2
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10765_ _03725_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19060_ _02662_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__clkbuf_1
X_12504_ rbzero.wall_tracer.trackDistX\[0\] _05257_ _05258_ rbzero.wall_tracer.trackDistX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o22a_1
XFILLER_201_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16272_ _08215_ _08226_ _08135_ _08160_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__or4_1
X_13484_ _06219_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and2_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10696_ rbzero.tex_g1\[9\] rbzero.tex_g1\[10\] _03680_ vssd1 vssd1 vccd1 vccd1 _03689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _01710_ _01711_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__and2_1
X_15223_ _07872_ _07868_ _07869_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__or3_1
XFILLER_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12435_ _05194_ _03914_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nor2_1
XFILLER_154_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15154_ _04034_ _07799_ _07807_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__a22o_1
X_12366_ _04891_ _04992_ _04890_ _04892_ _05091_ _05083_ vssd1 vssd1 vccd1 vccd1 _05134_
+ sky130_fd_sc_hd__mux4_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14105_ _06703_ _06841_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ _04075_ _04093_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__o21a_1
XFILLER_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19962_ _02695_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__buf_4
X_15085_ _07743_ _07744_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__nor2_1
X_12297_ _05062_ _05064_ _05065_ _05047_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a2bb2o_1
X_14036_ _06009_ _06658_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__nor2_1
XFILLER_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18913_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ _02558_ rbzero.spi_registers.spi_counter\[2\] vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a31o_1
X_11248_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__buf_2
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19893_ rbzero.pov.ready_buffer\[45\] _02823_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__nand2_1
XFILLER_122_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18844_ _02517_ _02518_ _02519_ _09807_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__o31a_1
XFILLER_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ _03957_ _03965_ _03966_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__and4b_1
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18775_ _02457_ _02458_ _02459_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15987_ _08630_ _08631_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__xor2_1
XFILLER_48_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17726_ _10039_ _10163_ _10290_ vssd1 vssd1 vccd1 vccd1 _10291_ sky130_fd_sc_hd__a21oi_1
X_14938_ rbzero.wall_tracer.visualWallDist\[4\] _07618_ vssd1 vssd1 vccd1 vccd1 _07635_
+ sky130_fd_sc_hd__or2_1
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17657_ _10216_ _10221_ vssd1 vssd1 vccd1 vccd1 _10222_ sky130_fd_sc_hd__and2_1
X_14869_ _07394_ _07440_ _07441_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__and3_1
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16608_ _09248_ _09250_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__and2_1
X_17588_ _09972_ _10010_ _10153_ vssd1 vssd1 vccd1 vccd1 _10154_ sky130_fd_sc_hd__a21boi_1
XFILLER_189_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19327_ rbzero.spi_registers.got_new_vshift _02730_ _02728_ _02813_ vssd1 vssd1 vccd1
+ vccd1 _00803_ sky130_fd_sc_hd__a31o_1
XFILLER_182_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16539_ _09156_ _09182_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19258_ _02772_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or3b_2
XFILLER_191_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__and2_1
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19189_ rbzero.floor_leak\[5\] _02732_ _02739_ _02722_ vssd1 vssd1 vccd1 vccd1 _00745_
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21220_ clknet_leaf_73_i_clk _00989_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_89_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20156__185 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__inv_2
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21151_ clknet_leaf_83_i_clk _00920_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21082_ net172 _00851_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20033_ _09753_ _03267_ _03274_ _03272_ _04884_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__a32o_1
XFILLER_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ clknet_leaf_64_i_clk _00704_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20321__333 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__inv_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20866_ clknet_leaf_66_i_clk _00635_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20797_ clknet_leaf_18_i_clk _00566_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10550_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _03602_ vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10481_ rbzero.tex_r0\[48\] rbzero.tex_r0\[47\] _03569_ vssd1 vssd1 vccd1 vccd1 _03576_
+ sky130_fd_sc_hd__mux2_1
X_12220_ gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__buf_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21418_ net339 _01187_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ _04906_ _04909_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nor2_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21349_ net270 _01118_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11102_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _03898_ vssd1 vssd1 vccd1 vccd1 _03902_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ net51 _04837_ net47 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a21o_1
XFILLER_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11033_ rbzero.tex_b0\[42\] rbzero.tex_b0\[41\] _03865_ vssd1 vssd1 vccd1 vccd1 _03866_
+ sky130_fd_sc_hd__mux2_1
X_15910_ _08008_ _07967_ vssd1 vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__nor2_1
XFILLER_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16890_ _09529_ _09530_ vssd1 vssd1 vccd1 vccd1 _09531_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _08137_ _08143_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _02167_ _02255_ _02256_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a21o_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _05596_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__xor2_4
X_15772_ _05208_ _08157_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__nor2_2
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17511_ _09526_ _08427_ vssd1 vssd1 vccd1 vccd1 _10077_ sky130_fd_sc_hd__nor2_1
X_11935_ _04709_ _04710_ _04247_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__mux2_1
X_14723_ _07456_ _07458_ _07459_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__mux2_1
XFILLER_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18491_ _02187_ _02188_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__nand2_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _05741_ _07383_ _07390_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a21oi_1
X_17442_ _09692_ _09717_ _10008_ vssd1 vssd1 vccd1 vccd1 _10009_ sky130_fd_sc_hd__a21o_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _04640_ _04641_ _04642_ _04139_ _04253_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__o221a_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20296__310 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__inv_2
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ _06292_ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__xnor2_1
X_10817_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _03751_ vssd1 vssd1 vccd1 vccd1 _03753_
+ sky130_fd_sc_hd__mux2_1
X_14585_ _07279_ _07282_ _07281_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__o21bai_1
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17373_ _09664_ _09665_ vssd1 vssd1 vccd1 vccd1 _09940_ sky130_fd_sc_hd__nand2_1
XFILLER_198_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ _04573_ _04574_ _04217_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19112_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ _02567_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__or4_2
X_13536_ _06225_ _06233_ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16324_ _08959_ _08967_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__or2_1
X_10748_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _03706_ vssd1 vssd1 vccd1 vccd1 _03716_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19043_ _02653_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
X_16255_ _08892_ _08899_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__xnor2_1
X_13467_ _06160_ _06202_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a21o_1
XFILLER_174_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10679_ _03646_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__clkbuf_4
X_15206_ _07821_ _07742_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__or2_1
XFILLER_103_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12418_ net37 _05184_ _05145_ net34 vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__and4bb_1
X_16186_ _08788_ _08830_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__nand2_1
X_13398_ _06065_ _06058_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__nor3_1
XFILLER_86_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15137_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__xnor2_1
X_12349_ net29 net28 _05116_ net30 vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a31o_1
XFILLER_141_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15068_ rbzero.debug_overlay.vplaneX\[-1\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__or2_1
X_19945_ rbzero.pov.ready_buffer\[58\] _03164_ _03197_ _03237_ vssd1 vssd1 vccd1 vccd1
+ _03238_ sky130_fd_sc_hd__o211a_1
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14019_ _06752_ _06754_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__and2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19876_ rbzero.debug_overlay.playerX\[4\] _03180_ vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__and2b_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18827_ _02503_ _02504_ _02505_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__nor3_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18758_ _02443_ _02444_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__and3_1
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17709_ _10123_ _10148_ _10145_ vssd1 vssd1 vccd1 vccd1 _10274_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18689_ _02252_ _02286_ _02384_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20720_ clknet_leaf_9_i_clk _00010_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20651_ clknet_leaf_5_i_clk _00435_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20582_ _07688_ _07831_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__nor2_1
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21203_ clknet_leaf_52_i_clk _00972_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21134_ clknet_leaf_60_i_clk _00903_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21065_ net155 _00834_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20016_ _03474_ _04809_ _03554_ _04815_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nor4_1
XFILLER_48_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11720_ _04022_ _04444_ _04440_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__and3_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ clknet_leaf_74_i_clk _00687_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _04008_ _04023_ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a21oi_2
XFILLER_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ clknet_leaf_93_i_clk _00618_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10602_ _03639_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14370_ _05893_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__buf_2
XFILLER_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11582_ rbzero.tex_r1\[23\] rbzero.tex_r1\[22\] _04290_ vssd1 vssd1 vccd1 vccd1 _04361_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _06053_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a21o_1
X_10533_ _03603_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16040_ _07923_ _08125_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__nor2_1
X_13252_ _05939_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__clkinv_2
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10464_ rbzero.tex_r0\[56\] rbzero.tex_r0\[55\] _03558_ vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12203_ _04966_ _04325_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__nor2_1
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _05834_ _05913_ _05914_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a31o_4
X_10395_ rbzero.tex_r1\[22\] rbzero.tex_r1\[23\] _03527_ vssd1 vssd1 vccd1 vccd1 _03529_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12134_ net11 net10 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__nor2_2
XFILLER_151_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17991_ _01691_ _01692_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__nand2_1
XFILLER_81_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19730_ rbzero.pov.spi_buffer\[39\] rbzero.pov.spi_buffer\[40\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
X_12065_ net7 net6 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nor2_1
XFILLER_78_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16942_ _09517_ _09582_ vssd1 vssd1 vccd1 vccd1 _09583_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11016_ rbzero.tex_b0\[50\] rbzero.tex_b0\[49\] _03854_ vssd1 vssd1 vccd1 vccd1 _03857_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20328__339 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__inv_2
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19661_ _03056_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16873_ _09478_ _09479_ _09513_ vssd1 vssd1 vccd1 vccd1 _09514_ sky130_fd_sc_hd__a21o_1
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18612_ _02218_ _02220_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__o21a_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _08439_ _08468_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__xor2_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _01620_ _09292_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__nor2_1
X_15755_ _08372_ _08399_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__xor2_1
X_12967_ _05591_ _05593_ _05628_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__o21a_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _07375_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__nor2_1
X_11918_ _04345_ _04693_ _04253_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o21a_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18474_ _08257_ _09027_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__nor2_1
XFILLER_166_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12898_ _05609_ _05619_ _05562_ _05566_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__o211a_1
XFILLER_61_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15686_ _08039_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__clkbuf_4
XFILLER_206_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17425_ _08873_ _09977_ _09991_ _08872_ vssd1 vssd1 vccd1 vccd1 _09992_ sky130_fd_sc_hd__o22a_1
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14637_ _05741_ _07348_ _07353_ _07373_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__a31o_1
XFILLER_53_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11849_ _04620_ _04622_ _04625_ _04306_ _04241_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a221o_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14568_ _07297_ _07299_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__xor2_1
XFILLER_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17356_ _08335_ _09483_ _09910_ vssd1 vssd1 vccd1 vccd1 _09923_ sky130_fd_sc_hd__o21ai_1
XFILLER_147_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16307_ _08950_ _08946_ _08671_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__a21o_1
X_13519_ _05921_ _06176_ _06215_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
X_14499_ _07188_ _07189_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__xor2_1
X_17287_ _09807_ _09859_ vssd1 vssd1 vccd1 vccd1 _09860_ sky130_fd_sc_hd__or2_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20073__109 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__inv_2
XFILLER_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19026_ _02644_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__clkbuf_1
X_16238_ _08881_ _08882_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__xor2_1
XFILLER_115_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _08791_ _08787_ _08790_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19928_ rbzero.debug_overlay.playerY\[1\] _03216_ rbzero.debug_overlay.playerY\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__o21ai_1
XFILLER_141_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19859_ rbzero.debug_overlay.playerX\[1\] _03167_ vssd1 vssd1 vccd1 vccd1 _03171_
+ sky130_fd_sc_hd__nor2_1
X_20268__286 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__inv_2
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_opt_3_0_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20703_ clknet_leaf_93_i_clk _00487_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20634_ clknet_leaf_76_i_clk _00418_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20565_ rbzero.traced_texVinit\[8\] _09764_ _07831_ _10027_ vssd1 vssd1 vccd1 vccd1
+ _01416_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_149_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20496_ _09750_ _03392_ _03394_ _03250_ rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1
+ _01397_ sky130_fd_sc_hd__a32o_1
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21117_ net207 _00886_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21048_ clknet_leaf_2_i_clk _00817_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13870_ _06552_ _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and2_2
XFILLER_47_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _07894_ _05456_ _08184_ _05193_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__a211o_1
X_12752_ _03926_ _05394_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nor2_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ rbzero.debug_overlay.facingY\[-6\] _04475_ _04458_ rbzero.debug_overlay.facingY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a22o_1
XFILLER_203_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15471_ _08097_ _08042_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__or2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__nand2_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14422_ _07114_ _07127_ _07157_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__a21oi_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ rbzero.wall_tracer.mapX\[9\] _05525_ vssd1 vssd1 vccd1 vccd1 _09792_ sky130_fd_sc_hd__and2_1
X_11634_ _04206_ _04412_ _04314_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a21o_1
X_18190_ _01887_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a21o_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14353_ _07044_ _07089_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17141_ rbzero.row_render.size\[4\] _09762_ _07541_ _07756_ vssd1 vssd1 vccd1 vccd1
+ _00532_ sky130_fd_sc_hd__a22o_1
X_11565_ rbzero.tex_r1\[7\] rbzero.tex_r1\[6\] _04342_ vssd1 vssd1 vccd1 vccd1 _04344_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13304_ _05846_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__buf_2
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10516_ _03594_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
X_17072_ _09710_ _09566_ _09711_ vssd1 vssd1 vccd1 vccd1 _09712_ sky130_fd_sc_hd__a21oi_2
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14284_ _06766_ _06767_ _06782_ _06781_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__a31o_1
X_11496_ _04274_ _04275_ _04226_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XFILLER_171_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13235_ _05800_ _05864_ _05970_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__o211a_1
XFILLER_143_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16023_ _08658_ _08662_ _08667_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__o21a_2
XFILLER_109_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10447_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ _05783_ _05757_ _05791_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10378_ rbzero.tex_r1\[30\] rbzero.tex_r1\[31\] _03516_ vssd1 vssd1 vccd1 vccd1 _03520_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ gpout0.vpos\[4\] gpout0.vpos\[5\] _04840_ vssd1 vssd1 vccd1 vccd1 _04889_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13097_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__clkbuf_4
X_17974_ _05203_ _01674_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or3b_1
XFILLER_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19616__69 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
X_19713_ rbzero.pov.spi_buffer\[31\] rbzero.pov.spi_buffer\[32\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03084_ sky130_fd_sc_hd__mux2_1
XFILLER_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12048_ rbzero.row_render.texu\[3\] _03473_ _04163_ vssd1 vssd1 vccd1 vccd1 _04822_
+ sky130_fd_sc_hd__or3b_1
X_16925_ _08816_ _09565_ vssd1 vssd1 vccd1 vccd1 _09566_ sky130_fd_sc_hd__nor2_1
XFILLER_172_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03313_ _03313_ vssd1 vssd1 vccd1 vccd1 clknet_0__03313_ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19644_ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16856_ _09495_ _09496_ vssd1 vssd1 vccd1 vccd1 _09497_ sky130_fd_sc_hd__nor2_1
XFILLER_168_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15807_ _08010_ _07997_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__nand2_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16787_ _08230_ rbzero.wall_tracer.stepDistY\[9\] vssd1 vssd1 vccd1 vccd1 _09429_
+ sky130_fd_sc_hd__nand2_1
X_13999_ _06719_ _06723_ _06734_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__and3_1
XFILLER_209_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18526_ _02223_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__inv_2
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _08276_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _02153_ _02154_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__nor2_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15669_ _07913_ _07996_ _07932_ _07924_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__o22ai_1
XFILLER_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17408_ _09553_ _09974_ _09687_ _09684_ vssd1 vssd1 vccd1 vccd1 _09975_ sky130_fd_sc_hd__a22o_1
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18388_ _01739_ _01860_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__or4_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17339_ _09594_ _09596_ _09737_ _09905_ vssd1 vssd1 vccd1 vccd1 _09906_ sky130_fd_sc_hd__a31oi_4
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20274__290 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__inv_2
XFILLER_134_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19009_ _02635_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21666_ clknet_leaf_43_i_clk _01435_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__03302_ clknet_0__03302_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03302_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20617_ clknet_leaf_71_i_clk _00401_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.d6 sky130_fd_sc_hd__dfxtp_2
X_21597_ net138 _01366_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11350_ rbzero.floor_leak\[1\] _04125_ _04129_ rbzero.floor_leak\[0\] vssd1 vssd1
+ vccd1 vccd1 _04130_ sky130_fd_sc_hd__o211a_1
XFILLER_193_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20548_ _03435_ _03436_ _03437_ _03430_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a22o_1
XFILLER_153_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10301_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__inv_2
XFILLER_152_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11281_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _04061_ sky130_fd_sc_hd__or2_1
XFILLER_134_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20479_ _03373_ _03377_ _03378_ _03379_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o211a_1
X_13020_ _05584_ _05714_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14971_ _00008_ _07514_ _07655_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__a21oi_1
X_16710_ _08162_ _09351_ vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__or2_1
X_13922_ _05825_ _06658_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__nor2_2
X_17690_ _08767_ _09693_ vssd1 vssd1 vccd1 vccd1 _10255_ sky130_fd_sc_hd__nor2_1
XFILLER_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _09283_ rbzero.wall_tracer.stepDistY\[8\] vssd1 vssd1 vccd1 vccd1 _09284_
+ sky130_fd_sc_hd__nand2_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13853_ _06219_ _06266_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__nor2_1
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19360_ rbzero.debug_overlay.vplaneY\[-7\] _02847_ vssd1 vssd1 vccd1 vccd1 _02849_
+ sky130_fd_sc_hd__or2_1
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ rbzero.wall_tracer.mapY\[8\] _05404_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__xor2_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16572_ rbzero.wall_tracer.visualWallDist\[8\] _04015_ vssd1 vssd1 vccd1 vccd1 _09215_
+ sky130_fd_sc_hd__nand2_4
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13784_ _06509_ _06519_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__xor2_1
X_10996_ _03846_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18311_ _01915_ _01916_ _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__and3_1
X_15523_ _08154_ _08167_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__xor2_1
XFILLER_31_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19291_ _02800_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__clkbuf_4
X_12735_ _05466_ _05468_ _05469_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__or4_1
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20104__138 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__inv_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _08275_ _09217_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__or2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ rbzero.map_rom.f4 _05410_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_1
X_15454_ _07971_ _05481_ _08098_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__o21ai_1
XFILLER_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14405_ _07140_ _07141_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__and2b_1
X_11617_ rbzero.tex_r1\[45\] rbzero.tex_r1\[44\] _04392_ vssd1 vssd1 vccd1 vccd1 _04396_
+ sky130_fd_sc_hd__mux2_1
X_18173_ _01865_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12597_ _05350_ _05293_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__xor2_2
X_15385_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerY\[-2\] _08029_
+ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__or3_1
X_17124_ _04422_ _09748_ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__nor2_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14336_ _06776_ _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__or2_1
XFILLER_156_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11548_ _04135_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__buf_4
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14267_ _06744_ _06751_ _06755_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__a21oi_2
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _05210_ rbzero.wall_tracer.stepDistX\[8\] vssd1 vssd1 vccd1 vccd1 _09695_
+ sky130_fd_sc_hd__nand2_4
X_11479_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _04213_ vssd1 vssd1 vccd1 vccd1 _04259_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13218_ _05952_ _05916_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a21oi_1
X_16006_ _08639_ _08650_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__xor2_1
X_14198_ _06769_ _06610_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__nor2_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _05884_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__nor2_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _01572_ _01659_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16908_ _09547_ _09548_ vssd1 vssd1 vccd1 vccd1 _09549_ sky130_fd_sc_hd__and2b_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17888_ _01580_ _01590_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__xor2_1
XFILLER_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16839_ _09351_ vssd1 vssd1 vccd1 vccd1 _09480_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19558_ _03028_ _03029_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18509_ _02067_ _02069_ _02066_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__o21ba_1
XFILLER_55_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ _02948_ _02954_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nand2_1
XFILLER_146_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21520_ net441 _01289_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20079__115 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__inv_2
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21451_ net372 _01220_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21382_ net303 _01151_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10850_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _03762_ vssd1 vssd1 vccd1 vccd1 _03770_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10781_ rbzero.tex_g0\[34\] rbzero.tex_g0\[33\] _03729_ vssd1 vssd1 vccd1 vccd1 _03734_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12520_ rbzero.wall_tracer.trackDistY\[3\] _05264_ _05269_ _05274_ vssd1 vssd1 vccd1
+ vccd1 _05275_ sky130_fd_sc_hd__a22o_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _05195_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__buf_4
X_21649_ clknet_leaf_18_i_clk _01418_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20290__305 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__inv_2
XFILLER_138_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11402_ rbzero.row_render.size\[7\] _04152_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15170_ _07823_ _07824_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__and2b_1
X_12382_ net34 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__inv_2
XFILLER_193_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14121_ _06699_ _06855_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ _04110_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__xnor2_4
XFILLER_158_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14052_ _06787_ _06788_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__xnor2_1
X_11264_ gpout0.vpos\[9\] gpout0.vpos\[8\] gpout0.vpos\[7\] net1 vssd1 vssd1 vccd1
+ vccd1 _04044_ sky130_fd_sc_hd__or4b_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13003_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__clkbuf_2
XFILLER_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18860_ _02128_ _02130_ _02533_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
X_11195_ _03919_ _03925_ rbzero.map_rom.a6 _03983_ rbzero.map_rom.f1 vssd1 vssd1 vccd1
+ vccd1 _03984_ sky130_fd_sc_hd__a2111o_1
X_17811_ _10115_ _01514_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__nand2_1
XFILLER_97_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18791_ _02472_ _02473_ _02474_ _02469_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__o211ai_1
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _08331_ _09610_ _10201_ _10200_ _09368_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__o32a_1
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14954_ rbzero.wall_tracer.visualWallDist\[9\] _07594_ vssd1 vssd1 vccd1 vccd1 _07646_
+ sky130_fd_sc_hd__or2_1
XFILLER_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13905_ _06595_ _06598_ _06640_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a21o_2
XFILLER_208_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17673_ _08044_ vssd1 vssd1 vccd1 vccd1 _10238_ sky130_fd_sc_hd__buf_2
X_14885_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.trackDistX\[-11\]
+ _07592_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__mux2_1
XFILLER_36_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19412_ _02893_ _02894_ _02895_ _02879_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a22o_1
X_16624_ _08383_ _09114_ _09121_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__or3_1
X_13836_ _06242_ _06244_ _06571_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__nand3_1
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand2_1
X_16555_ _09197_ _09198_ vssd1 vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__or2b_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13767_ _06501_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__and2_1
X_10979_ _03837_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15506_ _08150_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__buf_4
X_12718_ _05463_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__xnor2_2
X_19274_ rbzero.spi_registers.spi_cmd\[0\] _02772_ rbzero.spi_registers.spi_cmd\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__or3b_1
XFILLER_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16486_ _08242_ _09129_ _08170_ vssd1 vssd1 vccd1 vccd1 _09130_ sky130_fd_sc_hd__a21oi_2
X_13698_ _06431_ _06433_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__o21a_1
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18225_ _01918_ _01919_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a21oi_2
XFILLER_175_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15437_ _07951_ _08081_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__nand2_1
X_12649_ _05388_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nand2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _01743_ _01750_ _01856_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a21o_1
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15368_ _08011_ _07969_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__xor2_1
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17107_ rbzero.wall_tracer.texu\[5\] _09085_ _04035_ _09746_ vssd1 vssd1 vccd1 vccd1
+ _00516_ sky130_fd_sc_hd__o211a_1
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _07007_ _07012_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nand2_1
X_18087_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
X_15299_ _07942_ _07943_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__nand2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17038_ _09667_ _09677_ vssd1 vssd1 vccd1 vccd1 _09678_ sky130_fd_sc_hd__xor2_2
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ rbzero.pov.spi_buffer\[27\] rbzero.pov.ready_buffer\[27\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20951_ clknet_leaf_59_i_clk _00720_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20882_ clknet_leaf_60_i_clk _00651_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21503_ net424 _01272_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21434_ net355 _01203_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21365_ net286 _01134_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20316_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__buf_1
XFILLER_135_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21296_ net217 _01065_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20133__164 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__inv_2
XFILLER_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _04262_ vssd1 vssd1 vccd1 vccd1 _04727_
+ sky130_fd_sc_hd__mux2_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_107 vssd1 vssd1 vccd1 vccd1 ones[1] top_ew_algofoogle_107/LO sky130_fd_sc_hd__conb_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _03797_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14670_ _07218_ _07323_ _07345_ _07334_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__and4_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_118 vssd1 vssd1 vccd1 vccd1 ones[12] top_ew_algofoogle_118/LO sky130_fd_sc_hd__conb_1
X_11882_ _04139_ _04656_ _04657_ _04658_ _04208_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__o221a_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13621_ _05920_ _06009_ _06310_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__o21a_1
X_10833_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _03751_ vssd1 vssd1 vccd1 vccd1 _03761_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _08980_ _08984_ _08147_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__a21o_1
XFILLER_201_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13552_ _06286_ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__or2_1
X_10764_ rbzero.tex_g0\[42\] rbzero.tex_g0\[41\] _03718_ vssd1 vssd1 vccd1 vccd1 _03725_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__inv_2
X_13483_ _06212_ _06213_ _06218_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__or3_1
XFILLER_160_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16271_ _08215_ _08162_ _08160_ _08226_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__o22a_1
XFILLER_201_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10695_ _03688_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18010_ _01710_ _01711_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__nor2_1
XFILLER_200_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15222_ _07868_ _07869_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__o21ai_1
X_12434_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__buf_4
XFILLER_199_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ _04989_ _04990_ _05083_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__mux2_1
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ _04033_ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__nor2_1
XFILLER_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14104_ _06818_ _06840_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__xor2_1
X_11316_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__inv_2
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15084_ _07742_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _07744_
+ sky130_fd_sc_hd__and2_1
X_19961_ _03248_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__buf_2
X_12296_ net45 _05043_ _05049_ gpout3.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _05065_
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ _05984_ _06769_ _06658_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__a21o_1
X_18912_ rbzero.spi_registers.spi_counter\[2\] rbzero.spi_registers.spi_counter\[1\]
+ rbzero.spi_registers.spi_counter\[0\] _02558_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__and4_1
XFILLER_171_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11247_ _04003_ _03913_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__nor2_1
X_19892_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__buf_2
XFILLER_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18843_ _02517_ _02518_ _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11178_ rbzero.othery\[1\] _03942_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18774_ _02457_ _02458_ _02459_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__and3_1
XFILLER_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15986_ _07988_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__or3_1
XFILLER_208_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17725_ _10160_ _10162_ vssd1 vssd1 vccd1 vccd1 _10290_ sky130_fd_sc_hd__nor2_1
XFILLER_76_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.trackDistX\[4\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__mux2_1
XFILLER_209_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _10219_ _10220_ vssd1 vssd1 vccd1 vccd1 _10221_ sky130_fd_sc_hd__and2_1
X_14868_ _07583_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16607_ _09249_ _08356_ _09247_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__o21ai_1
X_13819_ _06333_ _06377_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__nor2_1
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ _10007_ _10009_ vssd1 vssd1 vccd1 vccd1 _10153_ sky130_fd_sc_hd__or2b_1
X_14799_ _07487_ _07456_ _07529_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__a21oi_4
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19326_ _02819_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__clkbuf_1
X_16538_ _09158_ _09181_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19257_ rbzero.spi_registers.got_new_sky _02730_ _02728_ _02781_ vssd1 vssd1 vccd1
+ vccd1 _00771_ sky130_fd_sc_hd__a31o_1
X_16469_ _09090_ _09112_ vssd1 vssd1 vccd1 vccd1 _09113_ sky130_fd_sc_hd__xor2_1
XFILLER_192_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18208_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nor2_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19188_ rbzero.spi_registers.new_leak\[5\] _02733_ vssd1 vssd1 vccd1 vccd1 _02739_
+ sky130_fd_sc_hd__or2_1
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ _01740_ _01742_ _01738_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a21bo_1
XFILLER_117_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21150_ clknet_leaf_83_i_clk _00919_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21081_ net171 _00850_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20032_ _02705_ _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nor2_1
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20934_ clknet_leaf_64_i_clk _00703_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19585__41 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20865_ clknet_leaf_65_i_clk _00634_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20796_ clknet_leaf_18_i_clk _00565_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10480_ _03575_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21417_ net338 _01186_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12150_ net11 net10 _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__and3b_1
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21348_ net269 _01117_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11101_ _03901_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12081_ net3 _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__and2_1
XFILLER_155_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21279_ clknet_leaf_59_i_clk _01048_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11032_ _03717_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_131_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _08479_ _08484_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__or2b_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15771_ _08124_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__clkinv_2
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _05563_ _05566_ _05594_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__and3_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _10073_ _10075_ vssd1 vssd1 vccd1 vccd1 _10076_ sky130_fd_sc_hd__nand2_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _05871_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__clkbuf_4
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11934_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _04263_ vssd1 vssd1 vccd1 vccd1 _04710_
+ sky130_fd_sc_hd__mux2_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ _01860_ _01475_ _01476_ _09141_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__o22ai_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _09714_ _09716_ vssd1 vssd1 vccd1 vccd1 _10008_ sky130_fd_sc_hd__nor2_1
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ _05741_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ rbzero.tex_g1\[1\] rbzero.tex_g1\[0\] _04336_ vssd1 vssd1 vccd1 vccd1 _04642_
+ sky130_fd_sc_hd__mux2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _05877_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__and3_1
X_10816_ _03752_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
X_17372_ _09641_ _09644_ _09643_ vssd1 vssd1 vccd1 vccd1 _09939_ sky130_fd_sc_hd__a21bo_1
X_14584_ _07304_ _07308_ _07315_ _07318_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__a41o_1
XFILLER_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11796_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _04341_ vssd1 vssd1 vccd1 vccd1 _04574_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19111_ _02557_ _02558_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__nand2_1
X_16323_ _08959_ _08967_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__nand2_1
X_13535_ _06269_ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__xor2_1
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _03715_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19042_ rbzero.pov.spi_buffer\[52\] rbzero.pov.ready_buffer\[52\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16254_ _08897_ _08898_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__nor2_1
X_13466_ _05974_ _06159_ _06161_ _05983_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__o22a_1
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _03679_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15205_ _07821_ _07742_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__nand2_1
X_12417_ _05146_ _04738_ _05183_ net35 net36 vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__o2111a_1
XFILLER_173_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ _07981_ _08128_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__nor2_1
X_13397_ _06084_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15136_ _07777_ _07792_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__or2_1
XFILLER_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12348_ _03473_ _04814_ _04317_ _04809_ _05083_ _05082_ vssd1 vssd1 vccd1 vccd1 _05116_
+ sky130_fd_sc_hd__mux4_1
XFILLER_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12279_ net42 _05046_ _05047_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and3_1
X_19944_ _03235_ _03920_ _03227_ _02822_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a31o_1
X_15067_ _07679_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__buf_4
XFILLER_141_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _06752_ _06754_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nor2_1
XFILLER_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19875_ _03138_ _03183_ rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1 vccd1
+ _03184_ sky130_fd_sc_hd__o21a_1
XFILLER_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18826_ _02498_ _02500_ _02497_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a21boi_1
XFILLER_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18757_ _02435_ _02437_ _02436_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__o21bai_1
XFILLER_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15969_ _08585_ _08613_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__nand2_1
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17708_ _10264_ _10272_ vssd1 vssd1 vccd1 vccd1 _10273_ sky130_fd_sc_hd__xnor2_2
XFILLER_110_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18688_ _02254_ _02285_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__and2_1
XFILLER_93_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ _10202_ _10203_ vssd1 vssd1 vccd1 vccd1 _10204_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20650_ clknet_leaf_5_i_clk _00434_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19309_ _02810_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20581_ _07687_ _07686_ _07685_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a21bo_1
XFILLER_177_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21202_ clknet_leaf_38_i_clk _00971_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21133_ clknet_leaf_62_i_clk _00902_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21064_ net154 _00833_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20015_ _03257_ _03258_ _03261_ _03209_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__o211a_1
XFILLER_189_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20245__265 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__inv_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20917_ clknet_leaf_74_i_clk _00686_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11650_ _04005_ _04023_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a21oi_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20848_ clknet_leaf_4_i_clk _00617_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ rbzero.tex_g1\[54\] rbzero.tex_g1\[55\] _03635_ vssd1 vssd1 vccd1 vccd1 _03639_
+ sky130_fd_sc_hd__mux2_1
X_11581_ rbzero.tex_r1\[21\] rbzero.tex_r1\[20\] _04290_ vssd1 vssd1 vccd1 vccd1 _04360_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20779_ clknet_leaf_22_i_clk _00548_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532_ rbzero.tex_r0\[24\] rbzero.tex_r0\[23\] _03602_ vssd1 vssd1 vccd1 vccd1 _03603_
+ sky130_fd_sc_hd__mux2_1
X_13320_ _05947_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _05941_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__clkbuf_4
X_10463_ _03566_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12202_ net19 vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__inv_2
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13182_ _05814_ _05915_ _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a21oi_1
X_10394_ _03528_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12133_ net12 net13 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__nor2_2
XFILLER_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17990_ _01688_ _01690_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__or2_1
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12064_ net5 net4 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__or2_1
X_16941_ _09579_ _09581_ vssd1 vssd1 vccd1 vccd1 _09582_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _03856_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19660_ rbzero.pov.spi_buffer\[6\] rbzero.pov.spi_buffer\[7\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16872_ _09498_ _09512_ vssd1 vssd1 vccd1 vccd1 _09513_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18611_ _02215_ _02217_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__or2_1
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _08464_ _08466_ _08467_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _02237_ _02238_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__xnor2_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _08391_ _08397_ _08398_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__a21oi_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _05701_ _05702_ _05683_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor3_4
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14705_ _05894_ _07041_ _07389_ _05741_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__a22o_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11917_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _04290_ vssd1 vssd1 vccd1 vccd1 _04693_
+ sky130_fd_sc_hd__mux2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _02169_ _02170_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__xnor2_1
X_15685_ _08035_ _08046_ _08329_ _08104_ vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__or4_1
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _05626_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__xor2_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _09990_ vssd1 vssd1 vccd1 vccd1 _09991_ sky130_fd_sc_hd__clkbuf_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _05779_ _07362_ _07372_ _05892_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__o211a_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11848_ _04623_ _04624_ _04304_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__mux2_1
XFILLER_92_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17355_ _08335_ _09483_ _09910_ vssd1 vssd1 vccd1 vccd1 _09922_ sky130_fd_sc_hd__or3_1
X_14567_ _07302_ _07303_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__nor2_1
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11779_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _04262_ vssd1 vssd1 vccd1 vccd1 _04557_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16306_ _08944_ _08948_ _08949_ _08950_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_140_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13518_ _06154_ _06205_ _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a21bo_1
XFILLER_174_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17286_ _09061_ _09062_ vssd1 vssd1 vccd1 vccd1 _09859_ sky130_fd_sc_hd__nand2_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14498_ _07227_ _07231_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__xor2_1
XFILLER_118_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19025_ rbzero.pov.spi_buffer\[44\] rbzero.pov.ready_buffer\[44\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16237_ _08857_ _08859_ _08855_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__a21boi_1
X_13449_ _06175_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16168_ _08791_ _08787_ _08790_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__and3_1
XFILLER_142_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15119_ _04462_ rbzero.debug_overlay.vplaneX\[-7\] _07774_ _07775_ vssd1 vssd1 vccd1
+ vccd1 _07777_ sky130_fd_sc_hd__nor4_1
XFILLER_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16099_ _08704_ _08706_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19927_ rbzero.debug_overlay.playerY\[2\] rbzero.debug_overlay.playerY\[1\] _03216_
+ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__or3_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19858_ rbzero.debug_overlay.playerX\[0\] _03139_ _03170_ net60 vssd1 vssd1 vccd1
+ vccd1 _00983_ sky130_fd_sc_hd__a211o_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18809_ rbzero.wall_tracer.trackDistY\[1\] _02490_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19642__92 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__inv_2
XFILLER_55_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19789_ _03123_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03289_ clknet_0__03289_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03289_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20702_ clknet_leaf_93_i_clk _00486_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20633_ clknet_leaf_76_i_clk _00417_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20564_ rbzero.traced_texVinit\[7\] _03443_ _09771_ _09739_ vssd1 vssd1 vccd1 vccd1
+ _01415_ sky130_fd_sc_hd__a22o_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20495_ _03393_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__inv_2
XFILLER_192_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21116_ net206 _00885_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21047_ clknet_leaf_87_i_clk _00816_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20169__196 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__inv_2
XFILLER_75_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ rbzero.wall_tracer.mapY\[11\] _05404_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__xnor2_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ rbzero.map_rom.f4 _05497_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__nand2_1
XFILLER_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _04040_ _04315_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__or2_1
X_15470_ _08110_ _08114_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__nand2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05422_ _05423_ _05428_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__o31ai_4
XFILLER_91_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ _07114_ _07127_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__and3_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ rbzero.color_sky\[1\] rbzero.color_floor\[1\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04412_ sky130_fd_sc_hd__mux2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _07536_ _09763_ rbzero.row_render.size\[3\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00531_ sky130_fd_sc_hd__a2bb2o_1
X_14352_ _07086_ _07088_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__xor2_1
XFILLER_196_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11564_ rbzero.tex_r1\[5\] rbzero.tex_r1\[4\] _04342_ vssd1 vssd1 vccd1 vccd1 _04343_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13303_ _06033_ _06036_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nand2_1
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10515_ rbzero.tex_r0\[32\] rbzero.tex_r0\[31\] _03591_ vssd1 vssd1 vccd1 vccd1 _03594_
+ sky130_fd_sc_hd__mux2_1
X_17071_ _09560_ _09561_ vssd1 vssd1 vccd1 vccd1 _09711_ sky130_fd_sc_hd__nor2_1
X_11495_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _04273_ vssd1 vssd1 vccd1 vccd1 _04275_
+ sky130_fd_sc_hd__mux2_1
X_14283_ _07017_ _07019_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__xor2_2
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16022_ _08657_ _08656_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__or2b_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13234_ _05725_ _05764_ _05793_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__mux2_1
X_10446_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__buf_4
XFILLER_171_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10377_ _03519_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13165_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__inv_2
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12116_ _04886_ _04887_ _04840_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__mux2_1
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13096_ _05700_ _05703_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__or2_1
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17973_ _01669_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__or2_1
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12047_ _04814_ _03473_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19712_ _03083_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__clkbuf_1
X_16924_ _09283_ rbzero.wall_tracer.stepDistY\[10\] _08235_ _09564_ vssd1 vssd1 vccd1
+ vccd1 _09565_ sky130_fd_sc_hd__a22oi_4
XFILLER_211_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03312_ _03312_ vssd1 vssd1 vccd1 vccd1 clknet_0__03312_ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19643_ _03020_ _03019_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__nand2_1
X_16855_ _09492_ _09494_ vssd1 vssd1 vccd1 vccd1 _09496_ sky130_fd_sc_hd__and2_1
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15806_ _08444_ _08450_ vssd1 vssd1 vccd1 vccd1 _08451_ sky130_fd_sc_hd__xor2_4
XFILLER_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16786_ _09426_ _09427_ vssd1 vssd1 vccd1 vccd1 _09428_ sky130_fd_sc_hd__xnor2_2
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ _06719_ _06723_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__a21oi_2
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18525_ _02138_ _02120_ _02221_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__and3_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _08375_ _08381_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__xor2_2
XFILLER_209_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _05582_ _05600_ _05628_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__o21a_1
XFILLER_179_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _10248_ _09991_ _02046_ _02045_ _10266_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__o32a_1
XFILLER_209_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15668_ _08298_ _08312_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__xor2_1
XFILLER_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17407_ _08895_ _09973_ vssd1 vssd1 vccd1 vccd1 _09974_ sky130_fd_sc_hd__nor2_1
X_14619_ _07354_ _07355_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__nor2_1
XFILLER_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18387_ _02085_ _01985_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__nand2_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15599_ _08183_ _08185_ _07602_ _08230_ _05208_ vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__a2111o_1
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17338_ _09592_ _09904_ _09736_ vssd1 vssd1 vccd1 vccd1 _09905_ sky130_fd_sc_hd__a21o_1
XFILLER_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _09812_ _09841_ _09842_ _09843_ vssd1 vssd1 vccd1 vccd1 _09844_ sky130_fd_sc_hd__o31ai_1
XFILLER_105_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19008_ rbzero.pov.spi_buffer\[36\] rbzero.pov.ready_buffer\[36\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20386__12 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
XFILLER_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03301_ clknet_0__03301_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03301_
+ sky130_fd_sc_hd__clkbuf_16
X_21665_ clknet_leaf_43_i_clk _01434_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20357__366 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__inv_2
XFILLER_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20616_ clknet_leaf_10_i_clk _00012_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_21596_ net137 _01365_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20547_ rbzero.traced_texa\[9\] rbzero.texV\[9\] _03432_ vssd1 vssd1 vccd1 vccd1
+ _03437_ sky130_fd_sc_hd__a21o_1
XFILLER_119_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__buf_2
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ rbzero.texV\[7\] _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__xor2_1
X_20478_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03379_
+ sky130_fd_sc_hd__nand2_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14970_ rbzero.wall_tracer.stepDistX\[-8\] _00008_ vssd1 vssd1 vccd1 vccd1 _07655_
+ sky130_fd_sc_hd__nor2_1
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13921_ _06615_ _06641_ _06642_ _06657_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a31o_4
XFILLER_207_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16640_ _08230_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__buf_4
X_13852_ _06568_ _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _05533_ _05542_ _05544_ _05284_ rbzero.wall_tracer.mapY\[7\] vssd1 vssd1
+ vccd1 vccd1 _00414_ sky130_fd_sc_hd__a32o_1
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16571_ _09212_ _09213_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__nand2_1
X_13783_ _06432_ _06504_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10995_ rbzero.tex_b0\[60\] rbzero.tex_b0\[59\] _03843_ vssd1 vssd1 vccd1 vccd1 _03846_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18310_ _01917_ _02009_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__xor2_1
X_15522_ _08165_ _08166_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__nor2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19290_ rbzero.spi_registers.spi_done _03480_ _02569_ vssd1 vssd1 vccd1 vccd1 _02800_
+ sky130_fd_sc_hd__and3_1
X_12734_ _05472_ _05475_ _05478_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__or4_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _01939_ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__xnor2_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _07893_ _05353_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _08098_
+ sky130_fd_sc_hd__o21a_1
XFILLER_128_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12665_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__buf_6
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14404_ _07122_ _07124_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__xnor2_1
X_11616_ _04393_ _04394_ _04304_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18172_ _01870_ _01872_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__xor2_1
XFILLER_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15384_ rbzero.debug_overlay.playerY\[-3\] _07952_ vssd1 vssd1 vccd1 vccd1 _08029_
+ sky130_fd_sc_hd__or2_1
X_12596_ _05294_ _05290_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__and2b_1
XFILLER_156_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17123_ _09756_ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__clkbuf_1
X_14335_ _06658_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__buf_2
X_11547_ rbzero.tex_r1\[14\] _04213_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__and2_1
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17054_ _08873_ _09693_ vssd1 vssd1 vccd1 vccd1 _09694_ sky130_fd_sc_hd__nor2_1
X_14266_ _07001_ _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__or2_2
XFILLER_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11478_ _04226_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or2_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16005_ _08640_ _08648_ _08649_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__a21oi_1
X_13217_ _05952_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__nor2_1
X_10429_ _03546_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14197_ _06929_ _06933_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13148_ _05713_ _05718_ _05721_ _05715_ _05778_ _05801_ vssd1 vssd1 vccd1 vccd1 _05885_
+ sky130_fd_sc_hd__mux4_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13079_ _05642_ _05636_ _05791_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__mux2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _01656_ _01658_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16907_ _09418_ _09422_ _09546_ _09542_ vssd1 vssd1 vccd1 vccd1 _09548_ sky130_fd_sc_hd__a211o_1
X_17887_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nor2_1
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19626_ clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__buf_1
X_16838_ _09404_ _09383_ vssd1 vssd1 vccd1 vccd1 _09479_ sky130_fd_sc_hd__or2b_1
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19557_ rbzero.pov.spi_counter\[2\] _03022_ _03020_ vssd1 vssd1 vccd1 vccd1 _03029_
+ sky130_fd_sc_hd__o21ai_1
X_16769_ _09270_ _09409_ _09410_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__a21o_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18508_ _02100_ _02062_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or2b_1
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19488_ _02904_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _02968_
+ sky130_fd_sc_hd__xor2_1
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18439_ _02131_ _02137_ rbzero.wall_tracer.trackDistX\[8\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00597_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_210_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21450_ net371 _01219_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21381_ net302 _01150_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20194_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__buf_1
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _03733_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ rbzero.debug_overlay.playerY\[0\] _03925_ _05204_ vssd1 vssd1 vccd1 vccd1
+ _05205_ sky130_fd_sc_hd__mux2_1
X_21648_ clknet_leaf_19_i_clk _01417_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ rbzero.row_render.size\[9\] _04153_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and2_1
X_12381_ net52 _05144_ _05139_ net49 _05147_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a221o_1
X_21579_ net500 _01348_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14120_ _06820_ _06838_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11332_ _04049_ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__xnor2_2
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14051_ _06777_ _06778_ _06779_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__a21bo_1
X_11263_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] _04042_ vssd1 vssd1 vccd1
+ vccd1 _04043_ sky130_fd_sc_hd__or4_1
XFILLER_141_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13002_ _05700_ _05732_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__or3b_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11194_ rbzero.map_rom.f4 rbzero.map_rom.d6 _03982_ _03924_ vssd1 vssd1 vccd1 vccd1
+ _03983_ sky130_fd_sc_hd__a22o_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17810_ _09292_ _09695_ _08767_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a21oi_2
X_18790_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__nand2_1
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20110__143 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__inv_2
X_17741_ _10204_ _10213_ _10211_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a21o_1
X_14953_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.trackDistX\[9\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13904_ _06595_ _06598_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__nand3_4
XFILLER_169_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17672_ _08259_ _09126_ _08493_ _08044_ vssd1 vssd1 vccd1 vccd1 _10237_ sky130_fd_sc_hd__or4_1
XFILLER_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14884_ _07591_ _07593_ _07596_ _04039_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__o211a_1
XFILLER_208_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19411_ _02879_ _02893_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nand4_2
X_16623_ _09240_ _09265_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__xnor2_1
X_13835_ _06242_ _06244_ _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__a21o_1
XFILLER_63_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16554_ _09194_ _09196_ vssd1 vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__nand2_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ _02829_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__and2_1
X_13766_ _05855_ _06153_ _06501_ _06502_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__nand4_1
XFILLER_204_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10978_ rbzero.tex_b1\[3\] rbzero.tex_b1\[4\] _03828_ vssd1 vssd1 vccd1 vccd1 _03837_
+ sky130_fd_sc_hd__mux2_1
XFILLER_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15505_ _08147_ _08149_ vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__or2_2
XFILLER_189_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19273_ rbzero.spi_registers.got_new_floor _02730_ _02728_ _02790_ vssd1 vssd1 vccd1
+ vccd1 _00778_ sky130_fd_sc_hd__a31o_1
X_12717_ _05421_ _05430_ _05433_ _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a31o_1
X_16485_ _05209_ rbzero.wall_tracer.stepDistX\[4\] vssd1 vssd1 vccd1 vccd1 _09129_
+ sky130_fd_sc_hd__nand2_2
XFILLER_189_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13697_ _06429_ _06430_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__or2b_1
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18224_ _01922_ _01923_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__nand2_1
X_15436_ _08080_ rbzero.debug_overlay.playerY\[-2\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _08081_ sky130_fd_sc_hd__mux2_1
X_12648_ _05389_ _05392_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__or2_1
XFILLER_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18155_ _01748_ _01749_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15367_ _07969_ _08011_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__or2b_1
XFILLER_102_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ _05320_ _05322_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17106_ _05194_ _09744_ _09745_ vssd1 vssd1 vccd1 vccd1 _09746_ sky130_fd_sc_hd__or3b_1
XFILLER_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14318_ _07053_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__or2_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18086_ _01786_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__nor2_1
XFILLER_102_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15298_ _07913_ _07932_ _07941_ _07924_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__o22ai_1
XFILLER_85_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17037_ _09673_ _09676_ vssd1 vssd1 vccd1 vccd1 _09677_ sky130_fd_sc_hd__xor2_2
X_14249_ _06909_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__nand2_1
XFILLER_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _02624_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__clkbuf_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17939_ _01639_ _01640_ _01635_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a21o_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20085__120 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__inv_2
XFILLER_113_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20950_ clknet_leaf_58_i_clk _00719_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20881_ clknet_leaf_61_i_clk _00650_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21502_ net423 _01271_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21433_ net354 _01202_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21364_ net285 _01133_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21295_ net216 _01064_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _04345_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__or2_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ rbzero.tex_b1\[40\] rbzero.tex_b1\[41\] _03795_ vssd1 vssd1 vccd1 vccd1 _03797_
+ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_108 vssd1 vssd1 vccd1 vccd1 ones[2] top_ew_algofoogle_108/LO sky130_fd_sc_hd__conb_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_119 vssd1 vssd1 vccd1 vccd1 ones[13] top_ew_algofoogle_119/LO sky130_fd_sc_hd__conb_1
X_11881_ rbzero.tex_g1\[30\] _04342_ _04126_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a21o_1
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13620_ _05990_ _06016_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__or2_1
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ _03760_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13551_ _05988_ _06287_ _06286_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__nor3_1
XFILLER_73_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10763_ _03724_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__inv_2
XFILLER_185_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16270_ _08863_ _08914_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__or2_1
X_13482_ _06212_ _06213_ _06218_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o21ai_1
XFILLER_200_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10694_ rbzero.tex_g1\[10\] rbzero.tex_g1\[11\] _03680_ vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15221_ _07870_ _07871_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__and2_1
X_12433_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__clkinv_4
XFILLER_200_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15152_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and2_1
X_12364_ _04886_ _04887_ _05083_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__mux2_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _06820_ _06838_ _06839_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _04069_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__or2_1
XFILLER_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15083_ _07742_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _07743_
+ sky130_fd_sc_hd__nor2_1
X_19960_ _02708_ _03137_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__nand2_4
X_12295_ net50 _05043_ _05063_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ _06002_ _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__and2_1
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18911_ _02579_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__clkbuf_1
X_11246_ _04029_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__buf_4
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19891_ net39 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__o21a_1
XFILLER_136_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18842_ _02510_ _02512_ _02511_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a21boi_1
X_11177_ rbzero.othery\[0\] rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15985_ _07980_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__or3_1
XFILLER_121_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18773_ _02450_ _02453_ _02451_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17724_ _10186_ _10288_ vssd1 vssd1 vccd1 vccd1 _10289_ sky130_fd_sc_hd__xnor2_1
X_14936_ _07621_ _07632_ _07633_ _07620_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__o211a_1
XFILLER_208_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17655_ _09522_ _08427_ _10218_ vssd1 vssd1 vccd1 vccd1 _10220_ sky130_fd_sc_hd__o21ai_1
X_14867_ rbzero.wall_tracer.stepDistY\[9\] _07582_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07583_ sky130_fd_sc_hd__mux2_1
XFILLER_91_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ _06464_ _06552_ _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a21bo_1
XFILLER_23_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ _09243_ vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17586_ _10109_ _10151_ vssd1 vssd1 vccd1 vccd1 _10152_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ _07486_ _07433_ _07442_ _07528_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__a31o_1
XFILLER_51_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ _09160_ _09180_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__xnor2_1
X_19325_ rbzero.spi_registers.new_vshift\[5\] rbzero.spi_registers.spi_buffer\[5\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
X_13749_ _06483_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__xor2_1
XFILLER_149_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16468_ _09110_ _09111_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__nor2_1
X_19256_ _02774_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__inv_2
XFILLER_176_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15419_ _08056_ _08063_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__xor2_1
X_18207_ _01906_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__or2_1
X_19187_ rbzero.floor_leak\[4\] _02732_ _02738_ _02722_ vssd1 vssd1 vccd1 vccd1 _00744_
+ sky130_fd_sc_hd__o211a_1
X_16399_ _09030_ _09043_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18138_ _01719_ _01721_ _01718_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a21bo_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20117__149 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__inv_2
X_18069_ _01768_ _01769_ _01753_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a21o_1
XFILLER_208_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21080_ net170 _00849_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20031_ _04884_ _02704_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__nor2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20933_ clknet_leaf_74_i_clk _00702_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20864_ clknet_leaf_59_i_clk _00633_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20795_ clknet_leaf_21_i_clk _00564_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21416_ net337 _01185_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21347_ net268 _01116_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ rbzero.tex_b0\[10\] rbzero.tex_b0\[9\] _03898_ vssd1 vssd1 vccd1 vccd1 _03901_
+ sky130_fd_sc_hd__mux2_1
X_12080_ net2 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__inv_2
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21278_ clknet_leaf_64_i_clk _01047_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_11031_ _03864_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15770_ _08059_ _08334_ _08335_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__or3_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _05716_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _07403_ _07457_ _07433_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__mux2_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _04263_ vssd1 vssd1 vccd1 vccd1 _04709_
+ sky130_fd_sc_hd__mux2_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17440_ _09986_ _10006_ vssd1 vssd1 vccd1 vccd1 _10007_ sky130_fd_sc_hd__xnor2_2
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _07386_ _07388_ _05931_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__mux2_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ rbzero.tex_g1\[2\] _04356_ _04126_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a21o_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20222__244 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__inv_2
X_13603_ _06065_ _05940_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nor2_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ rbzero.tex_g0\[18\] rbzero.tex_g0\[17\] _03751_ vssd1 vssd1 vccd1 vccd1 _03752_
+ sky130_fd_sc_hd__mux2_1
X_17371_ _09936_ _09937_ vssd1 vssd1 vccd1 vccd1 _09938_ sky130_fd_sc_hd__and2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14583_ _07316_ _07319_ _07317_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__a21oi_1
XFILLER_198_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11795_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _04211_ vssd1 vssd1 vccd1 vccd1 _04573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19110_ _02688_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__clkbuf_1
X_16322_ _08961_ _08966_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__xor2_1
X_13534_ _06211_ _06221_ _06270_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ rbzero.tex_g0\[50\] rbzero.tex_g0\[49\] _03706_ vssd1 vssd1 vccd1 vccd1 _03715_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19041_ _02652_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16253_ _08896_ _08893_ _08894_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__and3_1
X_13465_ _05974_ _06161_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__nor2_1
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10677_ rbzero.tex_g1\[18\] rbzero.tex_g1\[19\] _03669_ vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15204_ _07756_ _07845_ _07846_ _07856_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a31o_1
X_12416_ _05146_ net64 vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__nand2_1
XFILLER_173_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16184_ _08170_ _08042_ _08128_ _08180_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__o22a_1
X_13396_ _06065_ _06080_ _06084_ _06057_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__o22a_1
XFILLER_127_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15135_ _07778_ _07779_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__nor2_1
X_12347_ _05090_ _05102_ _05110_ _05114_ net30 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__a221oi_2
XFILLER_181_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15066_ _07727_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__clkbuf_1
X_19943_ _03235_ _03233_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__nor2_1
X_12278_ net23 net22 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__nor2_1
XFILLER_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14017_ _06753_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__inv_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__clkbuf_4
X_19874_ _02820_ _03180_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__nor2_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18825_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__and2_1
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18756_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__nand2_1
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15968_ _08609_ _08611_ _08612_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17707_ _10126_ _10269_ _10271_ vssd1 vssd1 vccd1 vccd1 _10272_ sky130_fd_sc_hd__a21oi_2
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14919_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.trackDistX\[-2\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__mux2_1
XFILLER_209_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15899_ _08511_ _08543_ vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__xor2_4
X_18687_ _02305_ _02306_ _02303_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__o21ba_1
XFILLER_91_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17638_ _08037_ _09704_ vssd1 vssd1 vccd1 vccd1 _10203_ sky130_fd_sc_hd__nor2_1
XFILLER_90_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _10134_ _10130_ _10131_ _10132_ vssd1 vssd1 vccd1 vccd1 _10135_ sky130_fd_sc_hd__a31o_1
XFILLER_210_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20197__221 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__inv_2
XFILLER_108_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19308_ rbzero.spi_registers.new_other\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
XFILLER_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20580_ _07685_ _07679_ _03451_ _03443_ rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__a32o_1
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19239_ rbzero.spi_registers.spi_done _02557_ _02558_ _02572_ vssd1 vssd1 vccd1 vccd1
+ _02771_ sky130_fd_sc_hd__and4b_1
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21201_ clknet_leaf_53_i_clk _00970_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21132_ clknet_leaf_60_i_clk _00901_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21063_ net153 _00832_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20014_ _03259_ _03260_ net71 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o21ai_1
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ clknet_leaf_74_i_clk _00685_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20847_ clknet_leaf_3_i_clk _00616_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10600_ _03638_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__clkbuf_1
X_11580_ _04357_ _04358_ _04329_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__mux2_1
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20778_ clknet_leaf_22_i_clk _00547_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10531_ _03557_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13250_ _05978_ _05982_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__or3_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _03558_ vssd1 vssd1 vccd1 vccd1 _03566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ _04966_ net64 _04969_ _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__a211o_1
XFILLER_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181_ _05844_ _05917_ _05834_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a21o_1
XFILLER_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10393_ rbzero.tex_r1\[23\] rbzero.tex_r1\[24\] _03527_ vssd1 vssd1 vccd1 vccd1 _03528_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12132_ net9 net8 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__nor2_2
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _09405_ _09444_ _09580_ vssd1 vssd1 vccd1 vccd1 _09581_ sky130_fd_sc_hd__a21o_1
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11014_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _03854_ vssd1 vssd1 vccd1 vccd1 _03856_
+ sky130_fd_sc_hd__mux2_1
XFILLER_133_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16871_ _09510_ _09511_ vssd1 vssd1 vccd1 vccd1 _09512_ sky130_fd_sc_hd__nor2_1
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18610_ _02305_ _02306_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _08440_ _08463_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__nor2_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _08373_ _08390_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__and2b_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18541_ _10238_ _09434_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__nor2_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _05673_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__buf_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11916_ _04329_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__or2_1
X_14704_ _05741_ _07383_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__or2_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _09661_ _09611_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__and2_1
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15684_ _08328_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__clkbuf_4
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _05609_ _05619_ _05622_ _05566_ _05562_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__o311a_1
XFILLER_79_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _05931_ _07371_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__or2_1
X_17423_ _09434_ _09988_ vssd1 vssd1 vccd1 vccd1 _09990_ sky130_fd_sc_hd__and2_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ rbzero.tex_g1\[37\] rbzero.tex_g1\[36\] _04392_ vssd1 vssd1 vccd1 vccd1 _04624_
+ sky130_fd_sc_hd__mux2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14566_ _07294_ _07301_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__nor2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _09679_ _09659_ vssd1 vssd1 vccd1 vccd1 _09921_ sky130_fd_sc_hd__or2b_1
XFILLER_198_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11778_ _04140_ _04539_ _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or3_1
XFILLER_158_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13517_ _06206_ _06200_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__or2b_1
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16305_ _08945_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__inv_2
XFILLER_53_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17285_ _09854_ _09855_ _09856_ vssd1 vssd1 vccd1 vccd1 _09858_ sky130_fd_sc_hd__o21a_1
X_10729_ _03557_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__clkbuf_4
X_14497_ _07184_ _07193_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19024_ _02643_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__clkbuf_1
X_16236_ _08825_ _08880_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__xor2_1
X_13448_ _06183_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__and2_1
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16167_ _08794_ _08796_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__xnor2_1
X_13379_ _05979_ _05909_ _05920_ _05900_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__or4b_2
XFILLER_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _04462_ rbzero.debug_overlay.vplaneX\[-7\] _07774_ _07775_ vssd1 vssd1 vccd1
+ vccd1 _07776_ sky130_fd_sc_hd__o22a_1
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16098_ _08722_ _08721_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__xor2_1
XFILLER_138_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ _07710_ _07711_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__or2b_1
X_19926_ rbzero.debug_overlay.playerY\[1\] _03193_ _03222_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00999_ sky130_fd_sc_hd__a211o_1
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19857_ rbzero.pov.ready_buffer\[68\] _03164_ _03155_ _03169_ vssd1 vssd1 vccd1 vccd1
+ _03170_ sky130_fd_sc_hd__o211a_1
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18808_ _05204_ _02488_ _02489_ _10173_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__a31o_1
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19788_ rbzero.pov.spi_buffer\[67\] rbzero.pov.spi_buffer\[68\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
XFILLER_49_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_89_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18739_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__nand2_1
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20701_ clknet_leaf_5_i_clk _00485_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20632_ clknet_leaf_75_i_clk _00416_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20563_ rbzero.traced_texVinit\[6\] _03443_ _09771_ _09597_ vssd1 vssd1 vccd1 vccd1
+ _01414_ sky130_fd_sc_hd__a22o_1
XFILLER_177_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20494_ _03389_ _03390_ _03391_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and3_1
XFILLER_121_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20251__270 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__inv_2
XFILLER_161_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21115_ net205 _00884_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21046_ clknet_leaf_88_i_clk _00815_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ rbzero.map_rom.f4 _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__or2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _04470_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__and2_1
XFILLER_203_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__nand2_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14420_ _07144_ _07156_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__xor2_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _04206_ _04374_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__and3b_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _07006_ _07026_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a21oi_1
XFILLER_168_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__clkbuf_8
XFILLER_156_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13302_ _06022_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10514_ _03593_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
X_17070_ _09560_ _09561_ vssd1 vssd1 vccd1 vccd1 _09710_ sky130_fd_sc_hd__nand2_1
X_14282_ _06774_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__nand2_1
XFILLER_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11494_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _04273_ vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20334__345 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__inv_2
X_16021_ _08621_ _08665_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__xnor2_4
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13233_ _05951_ _05924_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__nand2_1
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _03474_ _03554_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__or3_1
XFILLER_143_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _05743_ _05754_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__and2_1
X_10376_ rbzero.tex_r1\[31\] rbzero.tex_r1\[32\] _03516_ vssd1 vssd1 vccd1 vccd1 _03519_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__buf_2
XFILLER_151_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13095_ _05740_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_1
X_17972_ _01670_ _01673_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__and2_1
XFILLER_97_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19711_ rbzero.pov.spi_buffer\[30\] rbzero.pov.spi_buffer\[31\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03083_ sky130_fd_sc_hd__mux2_1
X_12046_ _04318_ _04810_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nor2_1
XFILLER_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16923_ _07585_ _09431_ _09563_ _09085_ vssd1 vssd1 vccd1 vccd1 _09564_ sky130_fd_sc_hd__a211o_1
XFILLER_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03311_ _03311_ vssd1 vssd1 vccd1 vccd1 clknet_0__03311_ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16854_ _09492_ _09494_ vssd1 vssd1 vccd1 vccd1 _09495_ sky130_fd_sc_hd__nor2_1
XFILLER_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _07976_ _08215_ _08446_ _08449_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__o31a_2
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13997_ _06732_ _06733_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__or2_1
X_16785_ _07598_ _09283_ _05209_ _09287_ vssd1 vssd1 vccd1 vccd1 _09427_ sky130_fd_sc_hd__or4_2
X_20405__6 clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
X_20380__387 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__inv_2
XFILLER_207_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18524_ _02138_ _02120_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a21o_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ _05577_ _05579_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__nand2_2
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15736_ _08259_ _08238_ _08379_ _08380_ vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__o31a_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18455_ _02151_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__xor2_1
X_12879_ _04030_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__and3_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15667_ _08306_ _08310_ _08311_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__a21oi_2
XFILLER_209_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17406_ _09540_ vssd1 vssd1 vccd1 vccd1 _09973_ sky130_fd_sc_hd__clkbuf_4
X_14618_ _07308_ _07315_ _07304_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__a21oi_1
X_18386_ _01982_ _01983_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__nand2_1
X_15598_ _08210_ _08213_ _07598_ _08002_ _05208_ vssd1 vssd1 vccd1 vccd1 _08243_ sky130_fd_sc_hd__a2111o_1
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14549_ _07270_ _07268_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__xor2_1
X_17337_ _09605_ _09606_ _09734_ vssd1 vssd1 vccd1 vccd1 _09904_ sky130_fd_sc_hd__or3_1
XFILLER_187_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17268_ _05531_ _09068_ vssd1 vssd1 vccd1 vccd1 _09843_ sky130_fd_sc_hd__nand2_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19007_ _02634_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16219_ _08854_ _08861_ _08863_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__a21oi_1
X_17199_ rbzero.wall_tracer.mapX\[7\] _05512_ vssd1 vssd1 vccd1 vccd1 _09783_ sky130_fd_sc_hd__and2_1
XFILLER_128_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19909_ _08070_ _03141_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__nor2_1
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21664_ clknet_leaf_47_i_clk _01433_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__03300_ clknet_0__03300_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03300_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20615_ clknet_leaf_10_i_clk _00011_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21595_ net136 _01364_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20546_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03436_
+ sky130_fd_sc_hd__nand2_1
XFILLER_192_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20477_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03378_
+ sky130_fd_sc_hd__or2_1
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20059__97 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__inv_2
XFILLER_43_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19606__60 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13920_ _06598_ _06643_ _06653_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__o211a_1
XFILLER_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21029_ clknet_leaf_51_i_clk _00798_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _06586_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__nand2_1
X_19621__74 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _05539_ _05543_ _05540_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o21bai_1
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13782_ _06515_ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__or2_1
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16570_ rbzero.wall_tracer.visualWallDist\[7\] _04015_ _08416_ _09211_ vssd1 vssd1
+ vccd1 vccd1 _09213_ sky130_fd_sc_hd__a31o_1
X_10994_ _03845_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15521_ _08155_ _08156_ _08164_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__nor3_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12733_ _05424_ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__xnor2_4
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15452_ _08096_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__buf_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ _10094_ _09162_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nor2_1
XFILLER_128_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05411_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__nor2_8
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _07136_ _07137_ _07139_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ rbzero.tex_r1\[41\] rbzero.tex_r1\[40\] _04392_ vssd1 vssd1 vccd1 vccd1 _04394_
+ sky130_fd_sc_hd__mux2_1
XFILLER_169_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18171_ _10248_ _09973_ _01746_ _01871_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__o31a_1
X_15383_ rbzero.debug_overlay.playerX\[-1\] rbzero.debug_overlay.playerX\[-2\] _08027_
+ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__or3_2
XFILLER_50_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12595_ _05347_ _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__and2_1
XFILLER_196_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14334_ _06705_ _07060_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__xor2_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17122_ _04430_ _09750_ vssd1 vssd1 vccd1 vccd1 _09756_ sky130_fd_sc_hd__and2_1
X_11546_ _04325_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkinv_2
XFILLER_129_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17053_ _09555_ vssd1 vssd1 vccd1 vccd1 _09693_ sky130_fd_sc_hd__clkbuf_4
X_14265_ _06999_ _07000_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__and2_1
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _04213_ vssd1 vssd1 vccd1 vccd1 _04257_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16004_ _08641_ _08647_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__nor2_1
X_13216_ _05725_ _05723_ _05893_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__mux2_1
X_10428_ rbzero.tex_r1\[6\] rbzero.tex_r1\[7\] _03538_ vssd1 vssd1 vccd1 vccd1 _03546_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14196_ _06805_ _06668_ _06928_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__o21bai_1
XFILLER_48_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13147_ _05820_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__buf_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ rbzero.tex_r1\[39\] net54 _03505_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _05640_ _05645_ _05648_ _05687_ _05795_ _05801_ vssd1 vssd1 vccd1 vccd1 _05815_
+ sky130_fd_sc_hd__mux4_1
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _01492_ _01538_ _01657_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12029_ _04244_ _04795_ _04803_ _04116_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a31o_1
X_16906_ _09542_ _09423_ _09546_ vssd1 vssd1 vccd1 vccd1 _09547_ sky130_fd_sc_hd__o21a_1
XFILLER_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17886_ _01586_ _01587_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__and2_1
XFILLER_211_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16837_ _09403_ _09386_ vssd1 vssd1 vccd1 vccd1 _09478_ sky130_fd_sc_hd__or2b_1
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19556_ rbzero.pov.spi_counter\[2\] _03022_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__and2_1
XFILLER_80_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16768_ _08284_ _09126_ _09276_ _08283_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__o22a_1
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18507_ _02099_ _02065_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__or2b_1
XFILLER_94_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719_ _08338_ _08339_ _08343_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__o21ba_1
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19487_ _02965_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__xnor2_1
X_16699_ _09207_ _09330_ _09328_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__a21bo_1
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18438_ _02135_ _02136_ _09780_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18369_ _02066_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__nor2_1
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21380_ net301 _01149_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20363__371 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__inv_2
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21647_ clknet_leaf_18_i_clk _01416_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11400_ rbzero.row_render.size\[9\] _04153_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nor2_1
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12380_ _04867_ _05145_ _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and3_1
XFILLER_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21578_ net499 _01347_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ rbzero.traced_texVinit\[11\] rbzero.texV\[11\] vssd1 vssd1 vccd1 vccd1 _04111_
+ sky130_fd_sc_hd__xor2_1
XFILLER_181_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20529_ _03416_ _03419_ _03417_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _06773_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__inv_2
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _04040_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_2
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13001_ _05733_ _05735_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__a211o_1
XFILLER_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11193_ _03942_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__inv_2
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17740_ _10232_ _10197_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__or2b_1
X_14952_ _04019_ _07643_ _07644_ _07642_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__o211a_1
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ _06616_ _06639_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__xnor2_2
X_17671_ _10112_ _10120_ _10119_ vssd1 vssd1 vccd1 vccd1 _10236_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14883_ rbzero.wall_tracer.visualWallDist\[-12\] _07595_ vssd1 vssd1 vccd1 vccd1
+ _07596_ sky130_fd_sc_hd__or2_1
XFILLER_75_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19410_ _02878_ _02880_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__or2b_1
X_16622_ _09263_ _09264_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__nand2_1
X_13834_ _06569_ _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__nand2_1
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19341_ _02830_ _02831_ _02829_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__nand3b_1
X_13765_ _06065_ _06031_ _06002_ _05877_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__a2bb2o_1
X_16553_ _09194_ _09196_ vssd1 vssd1 vccd1 vccd1 _09197_ sky130_fd_sc_hd__nor2_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _03836_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ rbzero.wall_tracer.visualWallDist\[3\] _08148_ vssd1 vssd1 vccd1 vccd1 _08149_
+ sky130_fd_sc_hd__nand2_4
XFILLER_206_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19272_ _02783_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__inv_2
X_12716_ _05437_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__inv_2
XFILLER_188_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13696_ _06383_ _06432_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__nand2_1
X_16484_ _08180_ _08971_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__nor2_1
XFILLER_189_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18223_ _01833_ _01836_ _01921_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__nand3_1
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12647_ _03935_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__xnor2_1
X_15435_ rbzero.debug_overlay.playerY\[-2\] _08029_ vssd1 vssd1 vccd1 vccd1 _08080_
+ sky130_fd_sc_hd__xor2_1
XFILLER_188_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15366_ _07997_ _08009_ _08010_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__a21bo_1
XFILLER_129_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18154_ _01819_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12578_ _05288_ _05319_ _05323_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__o21ai_1
XFILLER_106_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20191__216 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__inv_2
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _09470_ _09743_ _09600_ _09742_ vssd1 vssd1 vccd1 vccd1 _09745_ sky130_fd_sc_hd__a211o_1
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11529_ _04242_ _04298_ _04207_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o211a_1
X_14317_ _07050_ _07052_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and2_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15297_ _07913_ _07924_ _07932_ _07941_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__or4_1
X_18085_ _01684_ _01685_ _01785_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__and3_1
XFILLER_89_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ _06907_ _06908_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__or2_1
X_17036_ _08383_ _09674_ _09531_ _09675_ vssd1 vssd1 vccd1 vccd1 _09676_ sky130_fd_sc_hd__o31a_1
XFILLER_171_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14179_ _06905_ _06913_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__or2_1
XFILLER_124_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18987_ rbzero.pov.spi_buffer\[26\] rbzero.pov.ready_buffer\[26\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17938_ _01635_ _01639_ _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__nand3_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17869_ _01448_ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20880_ clknet_leaf_60_i_clk _00649_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19600__55 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_207_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19539_ rbzero.wall_tracer.rayAddendY\[10\] rbzero.wall_tracer.rayAddendY\[9\] _03001_
+ _02906_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__or4bb_1
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03039_ clknet_0__03039_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03039_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_210_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21501_ net422 _01270_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21432_ net353 _01201_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21363_ net284 _01132_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21294_ net215 _01063_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ _03796_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__clkbuf_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11880_ rbzero.tex_g1\[31\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__and3_1
Xtop_ew_algofoogle_109 vssd1 vssd1 vccd1 vccd1 ones[3] top_ew_algofoogle_109/LO sky130_fd_sc_hd__conb_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ rbzero.tex_g0\[10\] rbzero.tex_g0\[9\] _03751_ vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13550_ _05990_ _05975_ _05984_ _05991_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__o22a_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _03718_ vssd1 vssd1 vccd1 vccd1 _03724_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ _05254_ rbzero.wall_tracer.trackDistX\[2\] _05255_ rbzero.wall_tracer.trackDistX\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__o22a_1
XFILLER_198_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13481_ _06214_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__xnor2_1
X_10693_ _03687_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15220_ _07820_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _07871_
+ sky130_fd_sc_hd__or2_1
XFILLER_157_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12432_ _04002_ _03914_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nor2_1
XFILLER_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__or2_1
X_12363_ _04883_ _04884_ _05083_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__mux2_1
XFILLER_138_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _06821_ _06837_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__nor2_1
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11314_ _04065_ _04068_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__and2_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15082_ rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__buf_2
X_12294_ net49 _05044_ _05046_ net52 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a22o_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _06615_ _06641_ _06642_ _06657_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__a311oi_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18910_ _02557_ _02573_ _02578_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__and3_1
XFILLER_136_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11245_ _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__inv_2
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19890_ _03193_ _03195_ _03196_ _03157_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__o211a_1
XFILLER_107_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18841_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__and2_1
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _03960_ _03961_ _03962_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and4_1
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18772_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__nand2_1
X_15984_ _08559_ _08623_ _08624_ _08628_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17723_ _10285_ _10287_ vssd1 vssd1 vccd1 vccd1 _10288_ sky130_fd_sc_hd__xor2_1
XFILLER_76_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14935_ rbzero.wall_tracer.visualWallDist\[3\] _07618_ vssd1 vssd1 vccd1 vccd1 _07633_
+ sky130_fd_sc_hd__or2_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17654_ _09522_ _08425_ _10218_ vssd1 vssd1 vccd1 vccd1 _10219_ sky130_fd_sc_hd__or3_1
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _05929_ _07456_ _07581_ _07487_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__o31a_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16605_ _09243_ _08059_ _09247_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__or3_1
X_13817_ _06376_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__xor2_1
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17585_ _10147_ _10150_ vssd1 vssd1 vccd1 vccd1 _10151_ sky130_fd_sc_hd__xnor2_1
X_14797_ _07473_ _07471_ _07526_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__o211a_1
XFILLER_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19324_ _02818_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16536_ _09178_ _09179_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__and2_1
X_13748_ _06383_ _06432_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19255_ _02780_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16467_ _09091_ _08968_ _09109_ vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__and3_1
XFILLER_188_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13679_ _06395_ _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18206_ _01905_ _01799_ _01801_ _05203_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a31o_1
X_15418_ _08059_ _08062_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__nor2_1
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19186_ rbzero.spi_registers.new_leak\[4\] _02733_ vssd1 vssd1 vccd1 vccd1 _02738_
+ sky130_fd_sc_hd__or2_1
X_16398_ _09040_ _09042_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18137_ _01836_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__and2_1
X_15349_ _07925_ _07992_ _07993_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__a21oi_4
XFILLER_89_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18068_ _01753_ _01768_ _01769_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__nand3_1
XFILLER_208_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17019_ _09528_ _09535_ _09658_ vssd1 vssd1 vccd1 vccd1 _09659_ sky130_fd_sc_hd__a21o_1
X_20030_ _09753_ _03267_ _03271_ _03272_ _04883_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__a32o_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20932_ clknet_leaf_74_i_clk _00701_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ clknet_leaf_55_i_clk _00632_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20794_ clknet_leaf_20_i_clk _00563_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20174__200 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__inv_2
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21415_ net336 _01184_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21346_ net267 _01115_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21277_ clknet_leaf_63_i_clk _01046_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[0\]
+ sky130_fd_sc_hd__dfxtp_4
X_11030_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _03854_ vssd1 vssd1 vccd1 vccd1 _03864_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _05598_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__xor2_2
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _07431_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__clkinv_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _04210_ _04703_ _04707_ _04232_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a211o_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14651_ _07107_ _07356_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__a21bo_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11863_ rbzero.tex_g1\[3\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__and3_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _05995_ _06113_ _06057_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__a21oi_2
X_10814_ _03717_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _09926_ _09935_ vssd1 vssd1 vccd1 vccd1 _09937_ sky130_fd_sc_hd__or2_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14582_ _07294_ _07301_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__nand2_1
X_11794_ _04254_ _04567_ _04571_ _04241_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a211o_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16321_ _08964_ _08965_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__xnor2_1
X_13533_ _06183_ _06222_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__nor2_1
XFILLER_159_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10745_ _03714_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19040_ rbzero.pov.spi_buffer\[51\] rbzero.pov.ready_buffer\[51\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
X_13464_ _05923_ _05989_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__nand2_2
X_16252_ _08893_ _08894_ _08896_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__a21oi_1
X_10676_ _03678_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12415_ _05146_ net66 _05181_ net36 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a211o_1
X_15203_ _03913_ _07853_ _07854_ _07855_ rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__a32o_1
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _05824_ _06066_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__or2_1
X_16183_ _08194_ _08491_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__or2_1
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ _05101_ _05111_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__o21ba_1
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15134_ _07730_ rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 _07791_
+ sky130_fd_sc_hd__xor2_1
XFILLER_142_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ rbzero.wall_tracer.rayAddendX\[-2\] _07726_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07727_ sky130_fd_sc_hd__mux2_1
X_19942_ rbzero.debug_overlay.playerY\[5\] vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__inv_2
X_12277_ _05032_ net20 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__nor2_2
XFILLER_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _06680_ _06668_ _06714_ _06716_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__o31ai_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__buf_6
XFILLER_141_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19873_ rbzero.debug_overlay.playerX\[3\] _03143_ _03182_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00986_ sky130_fd_sc_hd__a211o_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18824_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nor2_1
X_11159_ rbzero.debug_overlay.playerX\[2\] _03929_ _03936_ rbzero.debug_overlay.playerX\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__o22a_1
XFILLER_68_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18755_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__or2_1
XFILLER_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15967_ _08586_ _08608_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__nor2_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17706_ _10270_ vssd1 vssd1 vccd1 vccd1 _10271_ sky130_fd_sc_hd__buf_4
XFILLER_208_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14918_ _04019_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__buf_2
X_18686_ _02325_ _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__xnor2_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _08539_ _08541_ _08542_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__a21oi_2
XFILLER_110_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17637_ _09368_ _10200_ _10201_ vssd1 vssd1 vccd1 vccd1 _10202_ sky130_fd_sc_hd__o21bai_1
XFILLER_64_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14849_ rbzero.wall_tracer.stepDistY\[5\] _07568_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07569_ sky130_fd_sc_hd__mux2_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17568_ _05211_ _09699_ _10128_ vssd1 vssd1 vccd1 vccd1 _10134_ sky130_fd_sc_hd__o21ai_4
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19307_ _02809_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16519_ _05209_ _09162_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__or2_1
XFILLER_32_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ _10062_ _10063_ vssd1 vssd1 vccd1 vccd1 _10065_ sky130_fd_sc_hd__nand2_1
XFILLER_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19238_ rbzero.spi_registers.vshift\[5\] _02762_ _02770_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00763_ sky130_fd_sc_hd__o211a_1
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19169_ rbzero.spi_registers.got_new_vinf vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__inv_2
XFILLER_129_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21200_ clknet_leaf_53_i_clk _00969_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21131_ clknet_leaf_59_i_clk _00900_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21062_ net152 _00831_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20013_ _04883_ _04992_ _03257_ _04884_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or4b_1
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20206__229 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__inv_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915_ clknet_leaf_75_i_clk _00684_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ clknet_leaf_4_i_clk _00615_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20777_ clknet_leaf_21_i_clk _00546_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10530_ _03601_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10461_ _03565_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12200_ _04966_ _04738_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nor2_1
XFILLER_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _05842_ _05916_ _05807_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__mux2_1
XFILLER_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10392_ _03482_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ net61 _04836_ _04839_ _04902_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__o31a_2
XFILLER_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21329_ net250 _01098_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12062_ clknet_leaf_46_i_clk vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__buf_1
XFILLER_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11013_ _03855_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16870_ _09507_ _09509_ vssd1 vssd1 vccd1 vccd1 _09511_ sky130_fd_sc_hd__and2_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _08169_ _08465_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__nor2_2
XFILLER_93_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _01737_ _10266_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__nor2_1
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _08392_ _08396_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__xnor2_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _05638_ _05649_ _05687_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__or3_2
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14703_ _07106_ _07415_ _07416_ _07417_ _05742_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__o311ai_2
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11915_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _04290_ vssd1 vssd1 vccd1 vccd1 _04691_
+ sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20146__176 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__inv_2
X_18471_ _02167_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _08148_ _08037_ _08038_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__a21oi_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _05623_ _05626_ _05628_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__o211a_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _09434_ _09988_ vssd1 vssd1 vccd1 vccd1 _09989_ sky130_fd_sc_hd__nand2_1
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14634_ _07366_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11846_ rbzero.tex_g1\[39\] rbzero.tex_g1\[38\] _04392_ vssd1 vssd1 vccd1 vccd1 _04623_
+ sky130_fd_sc_hd__mux2_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _09678_ _09660_ vssd1 vssd1 vccd1 vccd1 _09920_ sky130_fd_sc_hd__or2b_1
X_14565_ _07294_ _07301_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and2_1
X_11777_ _04142_ _04546_ _04554_ _04143_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__o211a_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _08941_ _08811_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__and2_1
X_13516_ _06251_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__and2_1
XFILLER_158_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10728_ _03705_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17284_ _09854_ _09855_ _09856_ vssd1 vssd1 vccd1 vccd1 _09857_ sky130_fd_sc_hd__nor3_1
X_14496_ _07227_ _07231_ _07232_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__a21o_1
XFILLER_159_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19023_ rbzero.pov.spi_buffer\[43\] rbzero.pov.ready_buffer\[43\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
X_16235_ _08816_ _08821_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__nor2_1
X_13447_ _06177_ _06178_ _06182_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__or3_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10659_ rbzero.tex_g1\[27\] rbzero.tex_g1\[28\] _03669_ vssd1 vssd1 vccd1 vccd1 _03670_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13378_ _06045_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__inv_2
XFILLER_154_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16166_ _08808_ _08810_ vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__xor2_4
XFILLER_127_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15117_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ _05090_ _05093_ _05094_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__and4_1
X_20311__324 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__inv_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _08700_ _08709_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15048_ _04462_ rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _07711_
+ sky130_fd_sc_hd__nand2_1
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19925_ rbzero.pov.ready_buffer\[54\] _03164_ _03197_ _03221_ vssd1 vssd1 vccd1 vccd1
+ _03222_ sky130_fd_sc_hd__o211a_1
XFILLER_170_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19856_ rbzero.debug_overlay.playerX\[0\] _08028_ _03168_ vssd1 vssd1 vccd1 vccd1
+ _03169_ sky130_fd_sc_hd__a21o_1
XFILLER_68_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18807_ _02481_ _02483_ _02486_ _02487_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__o211ai_2
XFILLER_96_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19787_ _03122_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16999_ _09501_ _09504_ _09503_ vssd1 vssd1 vccd1 vccd1 _09639_ sky130_fd_sc_hd__a21bo_1
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18738_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__or2_1
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401__26 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
XFILLER_83_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18669_ _02167_ _02255_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__nand2_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20700_ clknet_leaf_5_i_clk _00484_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20631_ clknet_leaf_76_i_clk _00415_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20562_ _07831_ _09458_ rbzero.traced_texVinit\[5\] _09762_ vssd1 vssd1 vccd1 vccd1
+ _01413_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20493_ _03389_ _03390_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a21o_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21114_ net204 _00883_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20286__301 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__inv_2
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21045_ clknet_leaf_88_i_clk _00814_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _04473_ _04478_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1
+ _04479_ sky130_fd_sc_hd__o211a_1
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05424_ _05425_ _05426_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__o211a_1
XFILLER_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11631_ _04207_ _04383_ _04391_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a31o_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ clknet_leaf_92_i_clk _00598_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14350_ _07023_ _07025_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__nor2_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11562_ _04128_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__buf_4
XFILLER_126_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13301_ _06024_ _06029_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o21ai_1
X_10513_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _03591_ vssd1 vssd1 vccd1 vccd1 _03593_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14281_ _06805_ _06761_ _06772_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__o21ai_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11493_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__buf_4
XFILLER_155_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13232_ _05901_ _05904_ _05964_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__a211o_1
X_16020_ _08654_ _08663_ _08664_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__a21oi_2
XFILLER_100_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10444_ _03479_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__clkinv_8
XFILLER_155_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13163_ _05846_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nor2_1
X_10375_ _03518_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__buf_2
XFILLER_152_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13094_ _05829_ _05830_ _05778_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__mux2_1
X_17971_ _01669_ _01670_ _01673_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__and3_1
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19710_ _03082_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
X_12045_ _04809_ _04810_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__xnor2_1
X_16922_ _07575_ _08983_ _09430_ _07586_ vssd1 vssd1 vccd1 vccd1 _09563_ sky130_fd_sc_hd__o31a_1
XFILLER_172_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03310_ _03310_ vssd1 vssd1 vccd1 vccd1 clknet_0__03310_ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16853_ _08335_ _09165_ _09354_ _09493_ vssd1 vssd1 vccd1 vccd1 _09494_ sky130_fd_sc_hd__o31a_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15804_ _08202_ _08238_ _08448_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__or3_1
X_16784_ _08377_ _09138_ vssd1 vssd1 vccd1 vccd1 _09426_ sky130_fd_sc_hd__nor2_1
XFILLER_207_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13996_ _06731_ _06700_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__and2_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18523_ _02218_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__xnor2_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15735_ _08303_ _08378_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__nand2_1
XFILLER_206_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12947_ _05673_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or2_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18454_ _10248_ _10266_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__nor2_1
XFILLER_179_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _08299_ _08305_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__nor2_1
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _05561_ _05466_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o21a_2
XFILLER_178_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17405_ _09957_ _09971_ vssd1 vssd1 vccd1 vccd1 _09972_ sky130_fd_sc_hd__xnor2_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _07304_ _07308_ _07315_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__and3_1
X_18385_ _01955_ _01957_ _01954_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a21bo_1
X_11829_ rbzero.tex_g1\[56\] _04272_ _04139_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a21o_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _08217_ _08225_ _05198_ vssd1 vssd1 vccd1 vccd1 _08242_ sky130_fd_sc_hd__o21ai_4
XFILLER_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17336_ rbzero.wall_tracer.trackDistX\[-1\] _09817_ _09897_ _09903_ vssd1 vssd1 vccd1
+ vccd1 _00588_ sky130_fd_sc_hd__o22a_1
XFILLER_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14548_ _07250_ _07272_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__xor2_1
XFILLER_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17267_ _09838_ _09839_ _09840_ vssd1 vssd1 vccd1 vccd1 _09842_ sky130_fd_sc_hd__o21a_1
X_14479_ _07200_ _07215_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__and2_1
XFILLER_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19006_ rbzero.pov.spi_buffer\[35\] rbzero.pov.ready_buffer\[35\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
X_16218_ _08250_ _08331_ _08862_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__and3_1
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ rbzero.wall_tracer.mapX\[6\] _05512_ _09778_ vssd1 vssd1 vccd1 vccd1 _09782_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16149_ _08776_ _08793_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19908_ rbzero.debug_overlay.playerY\[-4\] _03198_ _03208_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00994_ sky130_fd_sc_hd__o211a_1
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19839_ _05190_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20129__160 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__inv_2
XFILLER_45_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20281__297 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__inv_2
XFILLER_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21663_ clknet_leaf_47_i_clk _01432_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20614_ _03472_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21594_ net135 _01363_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20545_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03435_
+ sky130_fd_sc_hd__or2_1
XFILLER_71_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20476_ _03374_ _03375_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nor2_1
XFILLER_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21028_ clknet_leaf_50_i_clk _00797_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13850_ _06574_ _06585_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__or2_1
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12801_ rbzero.wall_tracer.mapY\[7\] _05404_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__nor2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13781_ _06503_ _06516_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__and3_1
X_10993_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _03843_ vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15520_ _08155_ _08156_ _08164_ vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__o21a_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20340__350 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__inv_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12732_ _05479_ _05425_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nor2_2
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _07945_ _08091_ _08095_ vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__o21ai_2
XFILLER_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12663_ rbzero.wall_tracer.state\[1\] _05211_ _04017_ _05278_ _05281_ vssd1 vssd1
+ vccd1 vccd1 _05412_ sky130_fd_sc_hd__o221ai_4
XFILLER_203_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14402_ _06724_ _06663_ _07138_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__nor3_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11614_ rbzero.tex_r1\[43\] rbzero.tex_r1\[42\] _04392_ vssd1 vssd1 vccd1 vccd1 _04393_
+ sky130_fd_sc_hd__mux2_1
X_18170_ _01744_ _01745_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__nand2_1
X_15382_ rbzero.debug_overlay.playerX\[-3\] _07946_ vssd1 vssd1 vccd1 vccd1 _08027_
+ sky130_fd_sc_hd__or2_1
XFILLER_168_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12594_ _05289_ _05295_ _05303_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a21o_1
XFILLER_168_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _04426_ _09748_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__nor2_1
XFILLER_129_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14333_ _07067_ _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__xor2_1
XFILLER_128_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20258__277 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__inv_2
X_11545_ _04047_ _04311_ _04313_ _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a31o_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17052_ _09682_ _09691_ vssd1 vssd1 vccd1 vccd1 _09692_ sky130_fd_sc_hd__xnor2_2
X_11476_ _04210_ _04248_ _04255_ _04232_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__a211o_1
X_14264_ _06999_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__nor2_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_88_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16003_ _08641_ _08647_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__xor2_1
X_10427_ _03545_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_1
X_13215_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14195_ _06923_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10358_ _03509_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
X_13146_ _05844_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nor2_1
XFILLER_151_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13077_ _05813_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__buf_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _01535_ _01537_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_1
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12028_ _04797_ _04799_ _04802_ _04306_ _04241_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a221o_1
X_16905_ _09544_ _09545_ vssd1 vssd1 vccd1 vccd1 _09546_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17885_ _01586_ _01587_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__nor2_1
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16836_ _09362_ _09377_ _09375_ vssd1 vssd1 vccd1 vccd1 _09477_ sky130_fd_sc_hd__a21o_1
XFILLER_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_207_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19555_ _03027_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16767_ _08284_ _09276_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__nor2_1
X_13979_ _06245_ _06678_ _06715_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__or3b_1
XFILLER_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ _02202_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__nor2_1
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15718_ _08361_ _08362_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19486_ _02938_ _02956_ _02958_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a21o_1
XFILLER_146_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16698_ _05194_ _09339_ _09340_ _07642_ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__o211a_1
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18437_ _02132_ _02133_ _02134_ _05204_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__o31a_1
X_15649_ _08292_ _08293_ vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__xnor2_1
XFILLER_210_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18368_ _01474_ _09350_ _01934_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__o21a_1
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17319_ _05532_ _09597_ vssd1 vssd1 vccd1 vccd1 _09888_ sky130_fd_sc_hd__and2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18299_ _01885_ _01887_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__and2_1
XFILLER_175_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21646_ clknet_leaf_18_i_clk _01415_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21577_ net498 _01346_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11330_ _04048_ _04051_ _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__o21ai_2
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20528_ rbzero.traced_texa\[7\] rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _03421_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11261_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nor2_1
X_20459_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03363_
+ sky130_fd_sc_hd__and2_1
X_13000_ _05649_ _05695_ _05673_ _05696_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__or4_4
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ _03933_ rbzero.map_rom.a6 rbzero.map_rom.i_row\[4\] _03974_ _03924_ vssd1
+ vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o32a_1
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14951_ rbzero.wall_tracer.visualWallDist\[8\] _07594_ vssd1 vssd1 vccd1 vccd1 _07644_
+ sky130_fd_sc_hd__or2_1
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13902_ _06617_ _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__xor2_2
XFILLER_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17670_ _10098_ _10106_ _10234_ vssd1 vssd1 vccd1 vccd1 _10235_ sky130_fd_sc_hd__a21o_1
X_14882_ _07594_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16621_ _09241_ _09242_ _09262_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__nand3_1
X_13833_ _05974_ _06245_ _06161_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__o21ai_1
XFILLER_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19340_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__or2_1
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16552_ rbzero.debug_overlay.playerX\[-5\] _07971_ _09195_ vssd1 vssd1 vccd1 vccd1
+ _09196_ sky130_fd_sc_hd__o21ai_2
X_13764_ _06065_ _05947_ _05975_ _05984_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__or4_1
XFILLER_204_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10976_ rbzero.tex_b1\[4\] rbzero.tex_b1\[5\] _03828_ vssd1 vssd1 vccd1 vccd1 _03836_
+ sky130_fd_sc_hd__mux2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15503_ _04014_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__buf_4
X_19271_ _02789_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ _05462_ _05440_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__nand2_1
X_16483_ _09126_ _08194_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__nor2_1
XFILLER_206_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13695_ _05824_ _06240_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__nor2_1
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18222_ _01833_ _01836_ _01921_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a21o_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15434_ _08077_ _08078_ _05496_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__mux2_1
X_12646_ _05374_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18153_ _01821_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ _07977_ _07995_ _07981_ _07989_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__or4_1
XFILLER_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ _05329_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _09461_ _09465_ _09600_ _09742_ _09743_ vssd1 vssd1 vccd1 vccd1 _09744_ sky130_fd_sc_hd__o311a_1
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14316_ _07050_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__nor2_1
XFILLER_117_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ _04230_ _04301_ _04232_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a211o_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18084_ _01684_ _01685_ _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15296_ _07940_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17035_ _09396_ _09669_ vssd1 vssd1 vccd1 vccd1 _09675_ sky130_fd_sc_hd__nand2_1
X_14247_ _06981_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__and2_1
X_11459_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _04214_ vssd1 vssd1 vccd1 vccd1 _04239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _06885_ _06911_ _06914_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__and3_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _05715_ _05721_ _05734_ _05718_ _05777_ _05801_ vssd1 vssd1 vccd1 vccd1 _05866_
+ sky130_fd_sc_hd__mux4_1
XFILLER_124_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _02623_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17937_ _01636_ _01637_ _01638_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a21o_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17868_ _01569_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__nor2_1
X_19597__52 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ _09458_ _09460_ vssd1 vssd1 vccd1 vccd1 _09461_ sky130_fd_sc_hd__nor2_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17799_ _09668_ _09973_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__nor2_1
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19538_ _03009_ _03013_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__nand2_1
XFILLER_185_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03038_ clknet_0__03038_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03038_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19469_ _02948_ _02949_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__nand2_1
X_21500_ net421 _01269_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21431_ net352 _01200_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21362_ net283 _01131_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21293_ net214 _01062_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10830_ _03759_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10761_ _03723_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12500_ rbzero.wall_tracer.trackDistY\[1\] vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__inv_2
XFILLER_197_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ _05921_ _06176_ _06215_ _06216_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__a31oi_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10692_ rbzero.tex_g1\[11\] rbzero.tex_g1\[12\] _03680_ vssd1 vssd1 vccd1 vccd1 _03687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12431_ _05192_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__clkbuf_1
X_21629_ clknet_leaf_19_i_clk _01398_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15150_ _07792_ _07791_ _07805_ _07775_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__o22a_1
XFILLER_194_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12362_ _05124_ _05129_ _05081_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__o21a_2
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14101_ _06821_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__xor2_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11313_ _04081_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o21a_1
XFILLER_126_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12293_ _05055_ net22 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nand2_1
X_15081_ _07729_ _07733_ _07731_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__a21bo_1
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14032_ _06016_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11244_ _03912_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nor2_1
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18840_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__nor2_1
XFILLER_84_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11175_ rbzero.otherx\[3\] _03936_ _03921_ rbzero.othery\[3\] _03963_ vssd1 vssd1
+ vccd1 vccd1 _03964_ sky130_fd_sc_hd__o221a_1
XFILLER_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20069__106 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__inv_2
XFILLER_122_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18771_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__or2_1
X_15983_ _08625_ _08627_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17722_ _10048_ _10159_ _10286_ vssd1 vssd1 vccd1 vccd1 _10287_ sky130_fd_sc_hd__a21oi_1
X_14934_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.trackDistX\[3\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__mux2_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _10074_ _10217_ vssd1 vssd1 vccd1 vccd1 _10218_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14865_ _07435_ _07436_ _07433_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__a21oi_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16604_ _09244_ _09246_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__nand2_1
X_13816_ _06336_ _06375_ _06424_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__o21ba_1
X_17584_ _10148_ _10149_ _10005_ _10006_ _09986_ vssd1 vssd1 vccd1 vccd1 _10150_ sky130_fd_sc_hd__a32o_1
X_14796_ _05834_ _05800_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__nor2_2
XFILLER_95_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ rbzero.spi_registers.new_vshift\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16535_ _09161_ _09166_ _09177_ vssd1 vssd1 vccd1 vccd1 _09179_ sky130_fd_sc_hd__o21bai_1
X_13747_ _06065_ _06240_ _06161_ _05824_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__o22a_1
X_10959_ rbzero.tex_b1\[12\] rbzero.tex_b1\[13\] _03817_ vssd1 vssd1 vccd1 vccd1 _03827_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19254_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_sky\[5\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16466_ _09091_ _08968_ _09109_ vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__a21oi_1
X_13678_ _06396_ _06413_ _06414_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18205_ _01799_ _01801_ _01905_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a21oi_1
X_15417_ _05193_ _07465_ _08061_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__a21oi_4
XFILLER_129_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19185_ rbzero.floor_leak\[3\] _02732_ _02737_ _02722_ vssd1 vssd1 vccd1 vccd1 _00743_
+ sky130_fd_sc_hd__o211a_1
X_12629_ _03933_ _05374_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__nor2_1
X_16397_ _08430_ _09041_ vssd1 vssd1 vccd1 vccd1 _09042_ sky130_fd_sc_hd__nor2_1
XFILLER_145_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18136_ _01826_ _01835_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__or2_1
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15348_ _07904_ rbzero.wall_tracer.stepDistY\[-3\] _05206_ vssd1 vssd1 vccd1 vccd1
+ _07993_ sky130_fd_sc_hd__a21o_1
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18067_ _01766_ _01767_ _01754_ _01647_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__o211ai_2
XFILLER_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15279_ _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__buf_2
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17018_ _09533_ _09534_ vssd1 vssd1 vccd1 vccd1 _09658_ sky130_fd_sc_hd__nor2_1
XFILLER_160_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _02614_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20931_ clknet_leaf_75_i_clk _00700_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20862_ clknet_leaf_55_i_clk _00631_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20793_ clknet_leaf_16_i_clk _00562_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21414_ net335 _01183_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21345_ net266 _01114_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21276_ clknet_leaf_65_i_clk _01045_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_104_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20227_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__buf_1
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ _05594_ _05596_ _05628_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__o21a_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _04704_ _04705_ _04706_ _04219_ _04254_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__o221a_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19576__33 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _05793_ _07369_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__nand2_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _04637_ _04638_ _04224_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__mux2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _05988_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _03750_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14581_ _07316_ _07317_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__nand2_1
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _04568_ _04569_ _04570_ _04225_ _04209_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o221a_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19591__47 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
X_16320_ _08282_ _07959_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__nor2_1
X_13532_ _06235_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10744_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _03706_ vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _08895_ _08579_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__or2_1
X_13463_ _06160_ _06162_ _06163_ _06164_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a22o_1
XFILLER_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ rbzero.tex_g1\[19\] rbzero.tex_g1\[20\] _03669_ vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15202_ _04028_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__clkbuf_4
X_12414_ _05146_ _04325_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__nor2_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16182_ _08820_ _08826_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__xor2_1
XFILLER_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13394_ _06129_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _07786_ _07787_ _07783_ _07784_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__a211o_1
X_12345_ net42 _05103_ _05085_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a31o_1
XFILLER_86_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15064_ _07720_ _07725_ _04033_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__mux2_1
X_19941_ _03231_ _03234_ _02714_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__o21a_1
X_12276_ net68 _05043_ _05044_ _04323_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a22o_1
XFILLER_135_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ _06744_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__xnor2_1
X_11227_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__clkinv_2
X_19872_ rbzero.pov.ready_buffer\[71\] _03146_ _03180_ _03181_ _03155_ vssd1 vssd1
+ vccd1 vccd1 _03182_ sky130_fd_sc_hd__o221a_1
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18823_ _02502_ _01553_ rbzero.wall_tracer.trackDistY\[3\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00616_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11158_ rbzero.wall_tracer.mapX\[7\] rbzero.wall_tracer.mapX\[6\] rbzero.wall_tracer.mapX\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or3_1
XFILLER_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15966_ _08584_ _08610_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__nor2_1
X_11089_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _03887_ vssd1 vssd1 vccd1 vccd1 _03895_
+ sky130_fd_sc_hd__mux2_1
X_18754_ _02442_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ _10125_ _10133_ _10135_ vssd1 vssd1 vccd1 vccd1 _10270_ sky130_fd_sc_hd__and3_1
X_14917_ _07591_ _07617_ _07619_ _07620_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__o211a_1
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ _08512_ _08538_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__nor2_1
X_18685_ _02375_ _02380_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ _07394_ _07464_ _07468_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__a21o_2
X_17636_ _09096_ _09480_ _09484_ _09368_ vssd1 vssd1 vccd1 vccd1 _10201_ sky130_fd_sc_hd__o22a_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _10130_ _10131_ _10132_ vssd1 vssd1 vccd1 vccd1 _10133_ sky130_fd_sc_hd__nand3_1
X_14779_ _07511_ _07447_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__nor2_1
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20123__155 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__inv_2
X_19306_ rbzero.spi_registers.new_other\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
X_16518_ rbzero.wall_tracer.visualWallDist\[7\] _04015_ vssd1 vssd1 vccd1 vccd1 _09162_
+ sky130_fd_sc_hd__nand2_2
XFILLER_143_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17498_ _10062_ _10063_ vssd1 vssd1 vccd1 vccd1 _10064_ sky130_fd_sc_hd__or2_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19237_ rbzero.spi_registers.new_vshift\[5\] _02763_ vssd1 vssd1 vccd1 vccd1 _02770_
+ sky130_fd_sc_hd__or2_1
X_16449_ _07941_ _08035_ _08046_ _08075_ vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__o22ai_1
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19168_ rbzero.othery\[4\] _02710_ _02725_ _02722_ vssd1 vssd1 vccd1 vccd1 _00738_
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18119_ _01751_ _01736_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__and2b_1
XFILLER_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19099_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.spi_buffer\[4\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
X_21130_ clknet_leaf_59_i_clk _00899_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21061_ net151 _00830_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20012_ _04892_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__inv_2
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ clknet_leaf_75_i_clk _00683_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20845_ clknet_leaf_3_i_clk _00614_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20776_ clknet_leaf_21_i_clk _00545_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20098__132 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__inv_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ rbzero.tex_r0\[58\] rbzero.tex_r0\[57\] _03558_ vssd1 vssd1 vccd1 vccd1 _03565_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10391_ _03526_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12130_ _04843_ _04845_ _04849_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__a31o_2
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21328_ net249 _01097_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ _04832_ _04834_ net68 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__a21oi_4
X_21259_ clknet_leaf_61_i_clk _01028_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_81_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11012_ rbzero.tex_b0\[52\] rbzero.tex_b0\[51\] _03854_ vssd1 vssd1 vccd1 vccd1 _03855_
+ sky130_fd_sc_hd__mux2_1
XFILLER_132_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15820_ _08120_ _08146_ _08168_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__and3_1
XFILLER_93_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _08393_ _08395_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__xnor2_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _05684_ _05689_ _05694_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__o211ai_4
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _07375_ _07435_ _07436_ _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__a31o_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11914_ _04686_ _04689_ _04209_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux2_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _08275_ _09484_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__nor2_1
X_15682_ _08297_ _08326_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__xor2_1
XFILLER_61_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12894_ _05454_ _05630_ _05561_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__mux2_1
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _05210_ rbzero.wall_tracer.stepDistX\[9\] vssd1 vssd1 vccd1 vccd1 _09988_
+ sky130_fd_sc_hd__nand2_2
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _05893_ _07369_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__nand2_1
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _04266_ _04621_ _04229_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__o21a_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _09638_ _09652_ _09650_ vssd1 vssd1 vccd1 vccd1 _09919_ sky130_fd_sc_hd__a21o_1
X_14564_ _07295_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__and2b_1
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _04253_ _04549_ _04553_ _04119_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a211o_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16303_ _08945_ _08947_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__xnor2_1
X_13515_ _06236_ _06250_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or2_1
X_17283_ _09846_ _09848_ _09847_ vssd1 vssd1 vccd1 vccd1 _09856_ sky130_fd_sc_hd__a21boi_1
X_10727_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _03624_ vssd1 vssd1 vccd1 vccd1 _03705_
+ sky130_fd_sc_hd__mux2_1
X_14495_ _07220_ _07226_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__nor2_1
XFILLER_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19022_ _02642_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16234_ _08877_ _08878_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__xnor2_1
X_13446_ _06177_ _06178_ _06182_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__o21ai_1
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10658_ _03646_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16165_ _08692_ _08718_ _08809_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__a21oi_2
XFILLER_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13377_ _05995_ _06113_ _05846_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a21o_1
XFILLER_170_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10589_ _03632_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15116_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__and2_1
X_12328_ _05087_ net66 _05095_ net30 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a211o_1
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16096_ _08733_ _08726_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ _04462_ rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _07710_
+ sky130_fd_sc_hd__nor2_1
X_19924_ rbzero.debug_overlay.playerY\[1\] _03216_ _03220_ vssd1 vssd1 vccd1 vccd1
+ _03221_ sky130_fd_sc_hd__a21o_1
X_12259_ _05021_ _04325_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__nor2_1
XFILLER_130_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19855_ _03145_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nand2_1
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18806_ _02486_ _02487_ _02481_ _02483_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a211o_1
X_20398__23 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
X_19786_ rbzero.pov.spi_buffer\[66\] rbzero.pov.spi_buffer\[67\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
XFILLER_110_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16998_ _09636_ _09637_ vssd1 vssd1 vccd1 vccd1 _09638_ sky130_fd_sc_hd__and2_1
XFILLER_96_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18737_ _02427_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15949_ _07990_ _08515_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__nand2_2
XFILLER_114_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18668_ _02350_ _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17619_ _09906_ _10183_ vssd1 vssd1 vccd1 vccd1 _10184_ sky130_fd_sc_hd__nor2_1
XFILLER_184_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18599_ _02179_ _02182_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20630_ clknet_leaf_76_i_clk _00414_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20561_ rbzero.traced_texVinit\[4\] _03443_ _09771_ _03444_ vssd1 vssd1 vccd1 vccd1
+ _01412_ sky130_fd_sc_hd__a22o_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20492_ _03384_ _03388_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__nand2_1
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21113_ net203 _00882_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21044_ clknet_leaf_77_i_clk _00813_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _04244_ _04400_ _04408_ _04116_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a31o_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20828_ clknet_leaf_92_i_clk _00597_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _04247_ _04334_ _04335_ _04339_ _04254_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__o221a_1
X_20759_ clknet_leaf_32_i_clk _00528_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13300_ _06030_ _06035_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nand3b_1
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10512_ _03592_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _06705_ _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__xnor2_2
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11492_ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__buf_4
XFILLER_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13231_ _05929_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__or2_1
X_10443_ _03475_ _03478_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nand2_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ _05834_ _05895_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a21oi_4
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10374_ rbzero.tex_r1\[32\] rbzero.tex_r1\[33\] _03516_ vssd1 vssd1 vccd1 vccd1 _03518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12113_ _04883_ _04884_ _04840_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__mux2_1
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ _05733_ _05705_ _05792_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__mux2_1
XFILLER_123_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17970_ _10294_ _10185_ _01550_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a31oi_4
X_20152__181 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__inv_2
XFILLER_78_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ rbzero.row_render.wall\[0\] rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1
+ vccd1 _04818_ sky130_fd_sc_hd__xnor2_2
X_16921_ _09560_ _09561_ vssd1 vssd1 vccd1 vccd1 _09562_ sky130_fd_sc_hd__xor2_1
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16852_ _09356_ _09357_ vssd1 vssd1 vccd1 vccd1 _09493_ sky130_fd_sc_hd__nand2_1
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _08446_ _08447_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__xnor2_4
X_19571_ clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__buf_1
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16783_ _09423_ _09424_ vssd1 vssd1 vccd1 vccd1 _09425_ sky130_fd_sc_hd__nor2_1
X_13995_ _06731_ _06700_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__nor2_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18522_ _01922_ _02219_ _02112_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__o21a_1
X_15734_ _08303_ _08378_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__xnor2_4
X_12946_ _05674_ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__or2_2
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _02045_ _02150_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__nand2_1
X_15665_ _08308_ _08309_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _04030_ _05337_ _05344_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a31o_1
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _05931_ _07352_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__or2_1
X_17404_ _09958_ _09970_ vssd1 vssd1 vccd1 vccd1 _09971_ sky130_fd_sc_hd__xnor2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _02081_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__and2_1
X_11828_ rbzero.tex_g1\[57\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__and3_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15596_ _08229_ _08240_ vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__xor2_2
XFILLER_92_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _09889_ _09901_ _09902_ _09780_ vssd1 vssd1 vccd1 vccd1 _09903_ sky130_fd_sc_hd__a31o_1
X_14547_ _07279_ _07283_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__xnor2_1
X_11759_ _04534_ _04535_ _04536_ _04224_ _04123_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__o221a_1
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17266_ _09838_ _09839_ _09840_ vssd1 vssd1 vccd1 vccd1 _09841_ sky130_fd_sc_hd__nor3_1
XFILLER_201_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14478_ _07213_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__nor2_1
XFILLER_128_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19005_ _02633_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__clkbuf_1
X_16217_ _08854_ _08861_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__xor2_1
X_13429_ _06158_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17197_ _09777_ _09778_ _09779_ _09781_ rbzero.wall_tracer.mapX\[6\] vssd1 vssd1
+ vccd1 vccd1 _00571_ sky130_fd_sc_hd__a32o_1
XFILLER_128_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20235__256 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__inv_2
XFILLER_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16148_ _08284_ _08579_ _08727_ vssd1 vssd1 vccd1 vccd1 _08793_ sky130_fd_sc_hd__nor3_1
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _08684_ _08686_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19907_ _05190_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__buf_4
XFILLER_116_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19838_ rbzero.debug_overlay.playerX\[-5\] _03155_ vssd1 vssd1 vccd1 vccd1 _03156_
+ sky130_fd_sc_hd__or2_1
XFILLER_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput1 i_debug_vec_overlay vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19769_ rbzero.pov.spi_buffer\[58\] rbzero.pov.spi_buffer\[59\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
XFILLER_209_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21662_ clknet_leaf_78_i_clk _01431_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20613_ _02721_ _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__and3_1
XFILLER_177_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21593_ net134 _01362_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20544_ _09750_ _03433_ _03434_ _03250_ rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1
+ _01405_ sky130_fd_sc_hd__a32o_1
XFILLER_193_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20475_ rbzero.texV\[-2\] _03175_ _03332_ _03376_ vssd1 vssd1 vccd1 vccd1 _01394_
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21027_ clknet_leaf_69_i_clk _00796_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_other
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12800_ _05539_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__or2b_1
XFILLER_210_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13780_ _06514_ _06513_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__xnor2_1
X_10992_ _03844_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__and2_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20392__18 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15450_ _05197_ _08094_ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__or2_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _03999_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__inv_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _07136_ _07137_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__xnor2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _04211_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__clkbuf_8
X_15381_ _08013_ _08025_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__or2b_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12593_ _05289_ _05295_ _05303_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__nand3_1
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _04417_ _09748_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__nor2_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14332_ _06675_ _06708_ _07064_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__o31a_1
X_11544_ _04314_ _04321_ _04323_ _04020_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a211o_1
XFILLER_168_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17051_ _09689_ _09690_ vssd1 vssd1 vccd1 vccd1 _09691_ sky130_fd_sc_hd__or2b_1
X_14263_ _06698_ _06726_ _06672_ _06729_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__o31a_1
XFILLER_52_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ _04219_ _04249_ _04252_ _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__o211a_1
XFILLER_183_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03289_ clknet_0__03289_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03289_
+ sky130_fd_sc_hd__clkbuf_16
X_16002_ _08644_ _08645_ _08646_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__a21oi_1
X_13214_ _05826_ _05893_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10426_ rbzero.tex_r1\[7\] rbzero.tex_r1\[8\] _03538_ vssd1 vssd1 vccd1 vccd1 _03545_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14194_ _06924_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13145_ _05710_ _05640_ _05648_ _05687_ _05778_ _05792_ vssd1 vssd1 vccd1 vccd1 _05882_
+ sky130_fd_sc_hd__mux4_1
XFILLER_87_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10357_ rbzero.tex_r1\[40\] rbzero.tex_r1\[41\] _03505_ vssd1 vssd1 vccd1 vccd1 _03509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _05754_ _05797_ _05700_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a21oi_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _01611_ _01655_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__xor2_1
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12027_ _04800_ _04801_ _04218_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__mux2_1
X_16904_ _07959_ _09126_ vssd1 vssd1 vccd1 vccd1 _09545_ sky130_fd_sc_hd__nor2_2
XFILLER_111_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17884_ _09391_ _09359_ _01463_ _10205_ _01462_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__o32a_1
XFILLER_39_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16835_ _09474_ _09475_ vssd1 vssd1 vccd1 vccd1 _09476_ sky130_fd_sc_hd__nor2_1
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19554_ _03022_ _03023_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__and3b_1
X_13978_ _06714_ _06674_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__xnor2_1
X_16766_ _09278_ _09280_ _09281_ _09277_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__a22oi_2
XFILLER_207_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _02200_ _02201_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__and2_1
X_12929_ _05650_ _05655_ _05664_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__o21ai_1
X_15717_ _07967_ _08097_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__or2_1
X_16697_ rbzero.wall_tracer.texu\[2\] _09085_ vssd1 vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__or2_1
X_19485_ _02963_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_1
XFILLER_207_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18436_ _02132_ _02133_ _02134_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__o21ai_1
X_15648_ _07996_ _07958_ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__nor2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18367_ _01474_ _09350_ _01934_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__nor3_1
X_15579_ _07970_ _08222_ _08223_ _07951_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__a31o_1
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17318_ _09887_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18298_ _01977_ _01997_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__xnor2_1
X_17249_ _08944_ _08948_ _04016_ vssd1 vssd1 vccd1 vccd1 _09826_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20260_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__buf_1
XFILLER_190_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ clknet_leaf_19_i_clk _01414_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21576_ net497 _01345_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_50 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20527_ rbzero.texV\[6\] _03327_ _03332_ _03420_ vssd1 vssd1 vccd1 vccd1 _01402_
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20218__240 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__inv_2
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__inv_2
XFILLER_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20458_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03362_
+ sky130_fd_sc_hd__nor2_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ rbzero.map_rom.f4 rbzero.map_rom.f3 _03973_ _03979_ vssd1 vssd1 vccd1 vccd1
+ _03980_ sky130_fd_sc_hd__a31o_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14950_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.trackDistX\[8\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__mux2_1
XFILLER_134_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13901_ _06619_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__xnor2_2
XFILLER_130_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14881_ _03969_ _04017_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__nor2_2
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13832_ _05974_ _06161_ _05940_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__or3_1
X_16620_ _09241_ _09242_ _09262_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__a21o_1
XFILLER_210_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20264__282 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__inv_2
XFILLER_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ rbzero.debug_overlay.playerY\[-5\] _07895_ vssd1 vssd1 vccd1 vccd1 _09195_
+ sky130_fd_sc_hd__or2_1
X_13763_ _06491_ _06492_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and2_1
X_10975_ _03835_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12714_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__nand2_1
X_15502_ _07945_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__buf_4
X_19270_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_floor\[5\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XFILLER_71_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16482_ _08189_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__clkbuf_4
X_13694_ _06429_ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__xor2_1
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18221_ _01920_ _01825_ _01823_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a21oi_1
X_15433_ rbzero.debug_overlay.playerX\[-2\] vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__inv_2
X_12645_ _05396_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15364_ _08008_ _07932_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__nor2_1
X_18152_ _01838_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12576_ _05324_ _05325_ _05328_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__nand3_1
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14315_ _06997_ _06726_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__o21a_1
X_17103_ _09599_ vssd1 vssd1 vccd1 vccd1 _09743_ sky130_fd_sc_hd__inv_2
XFILLER_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11527_ _04247_ _04302_ _04303_ _04305_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__o221a_1
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18083_ _01686_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__xor2_1
XFILLER_157_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15295_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__or2_1
XFILLER_102_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17034_ _09103_ vssd1 vssd1 vccd1 vccd1 _09674_ sky130_fd_sc_hd__clkbuf_4
X_14246_ _06944_ _06969_ _06975_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__and3_1
XFILLER_171_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ rbzero.tex_r0\[55\] _04221_ _04222_ _04219_ vssd1 vssd1 vccd1 vccd1 _04238_
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ rbzero.tex_r1\[15\] rbzero.tex_r1\[16\] _03527_ vssd1 vssd1 vccd1 vccd1 _03536_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14177_ _06905_ _06913_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__nand2_1
XFILLER_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11389_ _04161_ _04022_ gpout0.hpos\[3\] _04162_ _04168_ vssd1 vssd1 vccd1 vccd1
+ _04169_ sky130_fd_sc_hd__a221o_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13128_ _05798_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__nor2_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ rbzero.pov.spi_buffer\[25\] rbzero.pov.ready_buffer\[25\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor3_4
X_17936_ _01636_ _01637_ _01638_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nand3_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20347__357 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__inv_2
XFILLER_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17867_ _01561_ _01562_ _01568_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__and3_1
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16818_ _09459_ _08067_ _07895_ vssd1 vssd1 vccd1 vccd1 _09460_ sky130_fd_sc_hd__mux2_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17798_ _01500_ _01501_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__xnor2_2
XFILLER_66_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19537_ rbzero.wall_tracer.rayAddendY\[10\] _07695_ _07830_ _03012_ vssd1 vssd1 vccd1
+ vccd1 _03013_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16749_ _09245_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03037_ clknet_0__03037_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03037_
+ sky130_fd_sc_hd__clkbuf_16
X_19468_ _02904_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02949_
+ sky130_fd_sc_hd__or2_1
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19399_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__nor2_1
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21430_ net351 _01199_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21361_ net282 _01130_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20092__127 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__inv_2
XFILLER_163_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21292_ clknet_leaf_53_i_clk _01061_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_87_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10760_ rbzero.tex_g0\[44\] rbzero.tex_g0\[43\] _03718_ vssd1 vssd1 vccd1 vccd1 _03723_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10691_ _03686_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ net71 rbzero.wall_tracer.state\[7\] _05190_ vssd1 vssd1 vccd1 vccd1 _05192_
+ sky130_fd_sc_hd__and3_1
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21628_ clknet_leaf_19_i_clk _01397_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _05101_ _05126_ _05128_ _05085_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a2bb2o_1
X_21559_ net480 _01328_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14100_ _06822_ _06835_ _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a21boi_1
X_11312_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__inv_2
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15080_ _07728_ _07734_ _07740_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__a21o_1
X_12292_ net25 _05052_ _05060_ _05034_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__o211a_1
XFILLER_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14031_ _06766_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__nand2_1
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11243_ rbzero.wall_tracer.state\[14\] _04021_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_
+ sky130_fd_sc_hd__and3_2
XFILLER_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ rbzero.otherx\[3\] _03936_ _03919_ rbzero.otherx\[0\] vssd1 vssd1 vccd1 vccd1
+ _03963_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18770_ _02456_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__clkbuf_1
X_15982_ _08626_ _08039_ _08040_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__and3_1
XFILLER_121_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17721_ _10156_ _10158_ vssd1 vssd1 vccd1 vccd1 _10286_ sky130_fd_sc_hd__nor2_1
XFILLER_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14933_ _07621_ _07630_ _07631_ _07620_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__o211a_1
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17652_ _08445_ _08418_ vssd1 vssd1 vccd1 vccd1 _10217_ sky130_fd_sc_hd__nand2_1
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14864_ _07580_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16603_ _07932_ _08129_ _08047_ _09245_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__o22ai_1
X_13815_ _06548_ _06549_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14795_ _07473_ _07478_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__nand2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17583_ _09994_ _10002_ vssd1 vssd1 vccd1 vccd1 _10149_ sky130_fd_sc_hd__or2_1
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19322_ _02817_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__clkbuf_1
X_13746_ _06469_ _06471_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__nand2_1
X_16534_ _09161_ _09166_ _09177_ vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__or3b_1
XFILLER_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10958_ _03826_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19253_ _02779_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13677_ _06398_ _06412_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__nor2_1
X_16465_ _09098_ _09108_ vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10889_ _03790_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__clkbuf_1
X_18204_ _01903_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__or2_1
X_12628_ rbzero.map_rom.b6 _05374_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__and2_1
X_15416_ _07933_ _08060_ _07903_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__a21o_1
X_16396_ _08161_ _08431_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__nor2_1
X_19184_ rbzero.spi_registers.new_leak\[3\] _02733_ vssd1 vssd1 vccd1 vccd1 _02737_
+ sky130_fd_sc_hd__or2_1
XFILLER_157_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18135_ _01826_ _01835_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__nand2_1
X_15347_ _07545_ _07991_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07992_
+ sky130_fd_sc_hd__mux2_2
XFILLER_200_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12559_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nor2_1
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18066_ _01754_ _01647_ _01766_ _01767_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a211o_1
X_15278_ _07922_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__buf_2
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14229_ _06964_ _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__and2_1
XFILLER_160_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17017_ _09617_ _09656_ vssd1 vssd1 vccd1 vccd1 _09657_ sky130_fd_sc_hd__xnor2_2
XFILLER_176_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ rbzero.pov.spi_buffer\[17\] rbzero.pov.ready_buffer\[17\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_101_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _01619_ _01621_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__and2_1
X_18899_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] _02560_
+ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__and3_1
XFILLER_113_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20930_ clknet_leaf_75_i_clk _00699_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20861_ clknet_leaf_55_i_clk _00630_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20792_ clknet_leaf_20_i_clk _00561_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20100__134 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__inv_2
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21413_ net334 _01182_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21344_ net265 _01113_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21275_ clknet_leaf_65_i_clk _01044_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _04263_ vssd1 vssd1 vccd1 vccd1 _04706_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ rbzero.tex_g1\[7\] rbzero.tex_g1\[6\] _04336_ vssd1 vssd1 vccd1 vccd1 _04638_
+ sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _06293_ _06296_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__xnor2_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _03740_ vssd1 vssd1 vccd1 vccd1 _03750_
+ sky130_fd_sc_hd__mux2_1
X_14580_ _07273_ _07278_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__xor2_2
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11792_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _04262_ vssd1 vssd1 vccd1 vccd1 _04570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13531_ _06253_ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__xnor2_1
X_10743_ _03713_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16250_ _08283_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__clkbuf_4
X_13462_ _05752_ _06153_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__nand2_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10674_ _03677_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_1
X_20376__383 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__inv_2
XFILLER_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15201_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__or2_1
XFILLER_201_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12413_ _05146_ net61 _05179_ net36 vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__o211a_1
XFILLER_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16181_ _08816_ _08821_ _08825_ _08822_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__o31a_1
X_13393_ _06039_ _06048_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20075__111 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__inv_2
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15132_ _07788_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__inv_2
X_12344_ _05082_ _05083_ _04021_ _05085_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__and4_1
XFILLER_193_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15063_ _07723_ _07724_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__xnor2_1
X_19940_ rbzero.pov.ready_buffer\[57\] _03164_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__o21a_1
XFILLER_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12275_ net21 net20 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__nor2_2
XFILLER_126_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ _06745_ _06750_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__xnor2_1
X_11226_ _04011_ _04007_ _03478_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__a21bo_4
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19871_ rbzero.debug_overlay.playerX\[3\] _03176_ _02822_ vssd1 vssd1 vccd1 vccd1
+ _03181_ sky130_fd_sc_hd__a21o_1
XFILLER_96_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18822_ _09889_ _02501_ _02399_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a21boi_1
XFILLER_136_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11157_ _03940_ _03941_ _03943_ _03944_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a221o_1
XFILLER_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18753_ rbzero.wall_tracer.trackDistY\[-6\] _02440_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02442_ sky130_fd_sc_hd__mux2_1
XFILLER_95_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15965_ _08492_ _08566_ _08583_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__and3_1
X_11088_ _03894_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17704_ _10265_ _10268_ vssd1 vssd1 vccd1 vccd1 _10269_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14916_ _04035_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__buf_2
XFILLER_110_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18684_ _02377_ _02379_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _08509_ _08540_ vssd1 vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__nor2_1
XFILLER_48_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17635_ _09096_ _09480_ _09484_ vssd1 vssd1 vccd1 vccd1 _10200_ sky130_fd_sc_hd__or3_1
X_14847_ _07567_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _09117_ _10129_ vssd1 vssd1 vccd1 vccd1 _10132_ sky130_fd_sc_hd__nor2_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14778_ _07486_ _07433_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__nand2_1
XFILLER_204_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ _02808_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16517_ rbzero.wall_tracer.visualWallDist\[7\] _04015_ _09030_ _08416_ vssd1 vssd1
+ vccd1 vccd1 _09161_ sky130_fd_sc_hd__and4_1
X_13729_ _06453_ _06452_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__or2b_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17497_ _09368_ _09217_ _09929_ _09927_ vssd1 vssd1 vccd1 vccd1 _10063_ sky130_fd_sc_hd__o31a_1
XFILLER_189_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19236_ rbzero.spi_registers.vshift\[4\] _02762_ _02769_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00762_ sky130_fd_sc_hd__o211a_1
XFILLER_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16448_ _07941_ _08075_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__or4_1
XFILLER_158_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19167_ rbzero.spi_registers.new_other\[4\] _02712_ vssd1 vssd1 vccd1 vccd1 _02725_
+ sky130_fd_sc_hd__or2_1
X_16379_ _08327_ _08370_ _09023_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__a21oi_2
XFILLER_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18118_ _01715_ _01730_ _01818_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a21o_1
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19098_ _02682_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18049_ _01743_ _01750_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21060_ net150 _00829_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20011_ _04892_ _04992_ _04884_ _04883_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or4bb_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20913_ clknet_leaf_75_i_clk _00682_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20844_ clknet_leaf_12_i_clk _00613_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20775_ clknet_leaf_36_i_clk _00544_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10390_ rbzero.tex_r1\[24\] rbzero.tex_r1\[25\] _03516_ vssd1 vssd1 vccd1 vccd1 _03526_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21327_ net248 _01096_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _03474_ _04820_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a21o_1
X_21258_ clknet_leaf_62_i_clk _01027_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11011_ _03717_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__clkbuf_4
XFILLER_81_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21189_ clknet_leaf_76_i_clk _00958_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _05695_ _05673_ _05696_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__or4_2
X_15750_ _08394_ _08315_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__xor2_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _05963_ _07437_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__and2_1
X_11913_ _04687_ _04688_ _04139_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__mux2_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15681_ _08313_ _08324_ _08325_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__a21oi_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12893_ _04031_ _05329_ _05330_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a31o_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17420_ _09117_ _09693_ vssd1 vssd1 vccd1 vccd1 _09987_ sky130_fd_sc_hd__nor2_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _07367_ _07315_ _07368_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__o21ai_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ rbzero.tex_g1\[35\] rbzero.tex_g1\[34\] _04350_ vssd1 vssd1 vccd1 vccd1 _04621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _07297_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__nor2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _09908_ _09917_ vssd1 vssd1 vccd1 vccd1 _09918_ sky130_fd_sc_hd__xor2_4
XFILLER_207_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11775_ _04224_ _04550_ _04551_ _04552_ _04141_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__o221a_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16302_ _08941_ _08811_ _08946_ vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__a21oi_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _06236_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nand2_1
X_10726_ _03704_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14494_ _07229_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__and2b_1
X_17282_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09855_ sky130_fd_sc_hd__and2_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19021_ rbzero.pov.spi_buffer\[42\] rbzero.pov.ready_buffer\[42\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
X_13445_ _06179_ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16233_ _08830_ _08868_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10657_ _03668_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ _05889_ _05900_ _05910_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a21o_1
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ _08693_ _08717_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__nor2_1
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10588_ rbzero.tex_g1\[60\] rbzero.tex_g1\[61\] _03549_ vssd1 vssd1 vccd1 vccd1 _03632_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12327_ _05087_ _04325_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15115_ _07758_ _07761_ _07771_ _03912_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__a31o_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16095_ _08697_ _08712_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15046_ rbzero.debug_overlay.vplaneX\[-7\] _07705_ vssd1 vssd1 vccd1 vccd1 _07709_
+ sky130_fd_sc_hd__nand2_1
X_19923_ rbzero.debug_overlay.playerY\[1\] _03216_ _03145_ vssd1 vssd1 vccd1 vccd1
+ _03220_ sky130_fd_sc_hd__o21ai_1
X_12258_ net25 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__inv_2
XFILLER_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11209_ rbzero.wall_tracer.state\[1\] _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nand2_1
XFILLER_69_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19854_ rbzero.debug_overlay.playerX\[0\] _08028_ vssd1 vssd1 vccd1 vccd1 _03167_
+ sky130_fd_sc_hd__or2_1
XFILLER_69_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18805_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__nand2_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19785_ _03121_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16997_ _09626_ _09635_ vssd1 vssd1 vccd1 vccd1 _09637_ sky130_fd_sc_hd__or2_1
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18736_ rbzero.wall_tracer.trackDistY\[-8\] _02426_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02427_ sky130_fd_sc_hd__mux2_1
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _08591_ _08592_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18667_ _02351_ _02362_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ _08520_ _08521_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__and2_1
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17618_ _10165_ _10166_ _10026_ vssd1 vssd1 vccd1 vccd1 _10183_ sky130_fd_sc_hd__nand3b_1
XFILLER_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18598_ _02167_ _02168_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a21boi_1
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17549_ _08283_ _09555_ vssd1 vssd1 vccd1 vccd1 _10115_ sky130_fd_sc_hd__nor2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20560_ _09331_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__inv_2
XFILLER_177_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19219_ _09753_ _02758_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__and2_1
XFILLER_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20491_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03390_
+ sky130_fd_sc_hd__nand2_1
XFILLER_158_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21112_ net202 _00881_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20212__235 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__inv_2
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19618__71 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
XFILLER_119_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21043_ clknet_leaf_77_i_clk _00812_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19633__85 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__inv_2
XFILLER_80_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ clknet_leaf_92_i_clk _00596_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11560_ rbzero.tex_r1\[10\] _04338_ _04304_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a21o_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20758_ clknet_leaf_35_i_clk _00527_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.side
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ rbzero.tex_r0\[34\] rbzero.tex_r0\[33\] _03591_ vssd1 vssd1 vccd1 vccd1 _03592_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11491_ _04129_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__buf_4
X_20689_ clknet_leaf_26_i_clk _00473_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13230_ _05826_ _05934_ _05965_ _05966_ _05928_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__o221a_1
XFILLER_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10442_ _03553_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13161_ _05800_ _05896_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__o21a_1
X_10373_ _03517_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__buf_2
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13092_ _05757_ _05773_ _05792_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__mux2_1
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12043_ _04811_ _04813_ _04815_ _04816_ _04005_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a311o_1
X_16920_ _07598_ _09283_ _05210_ _09433_ vssd1 vssd1 vccd1 vccd1 _09561_ sky130_fd_sc_hd__or4_1
XFILLER_105_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20187__212 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__inv_2
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16851_ _09488_ _09491_ vssd1 vssd1 vccd1 vccd1 _09492_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15802_ _07974_ _08376_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__or2_2
X_19570_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__buf_1
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16782_ _09418_ _09422_ vssd1 vssd1 vccd1 vccd1 _09424_ sky130_fd_sc_hd__nor2_1
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13994_ _06729_ _06730_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__nand2_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ _02114_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__inv_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _08275_ _08377_ vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__nor2_2
X_12945_ _05677_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__or2_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _08802_ _09668_ _01524_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _08282_ _08194_ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__nor2_1
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ rbzero.wall_tracer.visualWallDist\[-3\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05613_ sky130_fd_sc_hd__a21o_1
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _09963_ _09969_ vssd1 vssd1 vccd1 vccd1 _09970_ sky130_fd_sc_hd__xor2_1
X_14615_ _07107_ _07349_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__a21o_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _04602_ _04603_ _04304_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux2_1
X_18383_ _02070_ _02080_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__or2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _08237_ _08239_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__nor2_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _09900_ _09893_ _09898_ _09899_ vssd1 vssd1 vccd1 vccd1 _09902_ sky130_fd_sc_hd__a211o_1
X_14546_ _07281_ _07282_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__nor2_1
X_11758_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _04341_ vssd1 vssd1 vccd1 vccd1 _04536_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10709_ rbzero.tex_g1\[3\] rbzero.tex_g1\[4\] _03691_ vssd1 vssd1 vccd1 vccd1 _03696_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17265_ _09830_ _09832_ _09831_ vssd1 vssd1 vccd1 vccd1 _09840_ sky130_fd_sc_hd__a21boi_1
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14477_ _07211_ _07212_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__and2_1
X_11689_ _04462_ _04463_ _04464_ rbzero.debug_overlay.vplaneX\[-4\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__a221o_1
X_19004_ rbzero.pov.spi_buffer\[34\] rbzero.pov.ready_buffer\[34\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
X_16216_ _08377_ _08062_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__nor2_1
X_13428_ _06163_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__xnor2_1
X_17196_ _09780_ vssd1 vssd1 vccd1 vccd1 _09781_ sky130_fd_sc_hd__buf_4
XFILLER_115_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13359_ _05941_ _05980_ _05990_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__a21oi_1
XFILLER_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16147_ _08787_ _08790_ _08791_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__a21bo_1
XFILLER_182_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ _08675_ _08720_ _08721_ _08722_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15029_ _07682_ _07693_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__xnor2_1
X_19906_ rbzero.pov.ready_buffer\[49\] _02823_ _03192_ _03207_ vssd1 vssd1 vccd1 vccd1
+ _03208_ sky130_fd_sc_hd__a211o_1
XFILLER_142_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19837_ net38 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__o21a_2
XFILLER_151_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput2 i_gpout0_sel[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_6
X_19768_ _03112_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18719_ _09863_ _02410_ _02411_ _09827_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__o31ai_1
X_19699_ _03076_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03299_ _03299_ vssd1 vssd1 vccd1 vccd1 clknet_0__03299_ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21661_ clknet_leaf_80_i_clk _01430_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20612_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__or2_1
XFILLER_51_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21592_ net133 _01361_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20543_ _03430_ _03431_ _03432_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__nand3_1
XFILLER_192_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20474_ _03374_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__xor2_1
XFILLER_119_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21026_ clknet_leaf_66_i_clk _00795_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10991_ rbzero.tex_b0\[62\] rbzero.tex_b0\[61\] _03843_ vssd1 vssd1 vccd1 vccd1 _03844_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12730_ rbzero.wall_tracer.rayAddendX\[-4\] rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\]
+ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__or4_1
XFILLER_128_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ rbzero.debug_overlay.playerX\[0\] _03919_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05410_ sky130_fd_sc_hd__mux2_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14400_ _06696_ _06708_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__nor2_1
X_11612_ _04230_ _04386_ _04390_ _04242_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__a211o_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _08014_ _08023_ _08024_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__a21bo_1
X_12592_ _05306_ _05343_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__xor2_2
XFILLER_129_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14331_ _06689_ _06663_ _07011_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__or3_1
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ gpout0.vpos\[5\] _04322_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _04323_
+ sky130_fd_sc_hd__a21o_4
XFILLER_156_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14262_ _06996_ _06998_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17050_ _09683_ _09688_ vssd1 vssd1 vccd1 vccd1 _09690_ sky130_fd_sc_hd__or2_1
X_11474_ _04253_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__buf_4
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ _05848_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__inv_2
X_16001_ _08642_ _08643_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__and2b_1
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _03544_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ _06895_ _06925_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__a21bo_1
XFILLER_87_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13144_ _05844_ _05880_ _05798_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__a21oi_2
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10356_ _03508_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13075_ _05802_ _05808_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__mux2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17952_ _01653_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__xor2_1
XFILLER_105_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12026_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _04250_ vssd1 vssd1 vccd1 vccd1 _04801_
+ sky130_fd_sc_hd__mux2_1
X_16903_ _09409_ _09543_ vssd1 vssd1 vccd1 vccd1 _09544_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17883_ _01584_ _01585_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__xor2_1
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16834_ _09379_ _09471_ _09473_ vssd1 vssd1 vccd1 vccd1 _09475_ sky130_fd_sc_hd__and3_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19612__66 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19553_ _03019_ _03025_ _03020_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a21boi_1
X_16765_ _09119_ _09270_ _09406_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__a21bo_1
X_13977_ _06240_ _06662_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or2_1
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18504_ _02200_ _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__nor2_1
XFILLER_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15716_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12928_ _05650_ _05655_ _05664_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or3_1
XFILLER_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19484_ _02905_ _04471_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1
+ _02964_ sky130_fd_sc_hd__or3b_1
X_16696_ _09082_ _09338_ vssd1 vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18435_ _02017_ _02019_ _02018_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a21boi_1
X_15647_ _08290_ _08291_ vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__xnor2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20241__261 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__inv_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _05477_ _05595_ _05560_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__mux2_4
XFILLER_181_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18366_ _02063_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nand2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ _07893_ _05372_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__or2_2
X_17317_ rbzero.wall_tracer.trackDistX\[-3\] _09886_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09887_ sky130_fd_sc_hd__mux2_1
X_14529_ _07264_ _07265_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__and2b_1
X_18297_ _01979_ _01996_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _09823_ _09821_ _09822_ _05531_ vssd1 vssd1 vccd1 vccd1 _09825_ sky130_fd_sc_hd__a31o_1
X_20159__188 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__inv_2
XFILLER_127_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17179_ rbzero.traced_texa\[7\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a22o_1
XFILLER_192_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20324__336 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__inv_2
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21644_ clknet_leaf_19_i_clk _01413_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21575_ net496 _01344_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_40 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 _10027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20526_ _03418_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20457_ _03272_ _03360_ _03361_ _03327_ rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1
+ _01391_ sky130_fd_sc_hd__a32o_1
XFILLER_134_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20370__378 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__inv_2
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11190_ _03919_ _03925_ _03976_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a31o_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _06635_ _06636_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21009_ clknet_leaf_49_i_clk _00778_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_floor
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14880_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.trackDistX\[-12\]
+ _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__mux2_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_i_clk clknet_1_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ _06253_ _06267_ _06251_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__a21bo_1
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16550_ _09088_ _09193_ vssd1 vssd1 vccd1 vccd1 _09194_ sky130_fd_sc_hd__xnor2_4
X_13762_ _06461_ _06458_ _06460_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__and3_1
X_20299__313 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__inv_2
X_10974_ rbzero.tex_b1\[5\] rbzero.tex_b1\[6\] _03828_ vssd1 vssd1 vccd1 vccd1 _03835_
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ _08122_ _08145_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__or2b_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _05442_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and2_1
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16481_ _09116_ _09124_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13693_ _05945_ _06409_ _06078_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18220_ _01822_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__inv_2
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15432_ rbzero.debug_overlay.playerX\[-2\] _08027_ vssd1 vssd1 vccd1 vccd1 _08077_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_54_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12644_ _05395_ rbzero.map_rom.a6 _05284_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _01850_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__nor2_1
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _05324_ _05325_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__a21o_1
X_15363_ _07945_ _08001_ _08006_ _08007_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__a22o_4
XFILLER_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17102_ _09739_ _09741_ vssd1 vssd1 vccd1 vccd1 _09742_ sky130_fd_sc_hd__xnor2_1
X_14314_ _06996_ _06998_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__nand2_1
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ _04209_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__buf_6
X_18082_ _01781_ _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15294_ _05197_ rbzero.wall_tracer.stepDistX\[-5\] vssd1 vssd1 vccd1 vccd1 _07939_
+ sky130_fd_sc_hd__nor2_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17033_ _09669_ _09672_ vssd1 vssd1 vccd1 vccd1 _09673_ sky130_fd_sc_hd__xnor2_2
X_14245_ _06962_ _06979_ _06981_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__and3b_1
X_11457_ rbzero.tex_r0\[54\] _04214_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__and2_1
X_10408_ _03535_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
X_14176_ _06911_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__and2_1
XFILLER_124_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11388_ _04147_ gpout0.hpos\[2\] gpout0.hpos\[3\] _04162_ _04167_ vssd1 vssd1 vccd1
+ vccd1 _04168_ sky130_fd_sc_hd__o221a_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _03499_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
X_13127_ _05859_ _05863_ _05811_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__mux2_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _02622_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__clkbuf_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _05759_ _05772_ _05775_ _05699_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__nor4b_2
X_17935_ _10110_ _09977_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__nor2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12009_ rbzero.tex_b1\[59\] rbzero.tex_b1\[58\] _04350_ vssd1 vssd1 vccd1 vccd1 _04784_
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17866_ _01561_ _01562_ _01568_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16817_ rbzero.debug_overlay.playerY\[-3\] vssd1 vssd1 vccd1 vccd1 _09459_ sky130_fd_sc_hd__clkinv_2
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17797_ _10239_ _08057_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nor2_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19536_ _03010_ _03011_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__xnor2_1
X_16748_ _09245_ _08059_ _09389_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__or3_1
X_20165__192 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__inv_2
XFILLER_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19467_ _02904_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02948_
+ sky130_fd_sc_hd__nand2_1
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16679_ _09181_ _09158_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__or2b_1
XFILLER_185_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18418_ _01928_ _02004_ _02003_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a21oi_2
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19398_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__and2_1
XFILLER_107_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _10248_ _09991_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__nor2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21360_ net281 _01129_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21291_ clknet_leaf_42_i_clk _01060_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ rbzero.tex_g1\[12\] rbzero.tex_g1\[13\] _03680_ vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21627_ clknet_leaf_20_i_clk _01396_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _05127_ _05099_ _05107_ net1 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21558_ net479 _01327_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ _04075_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__or2_1
XFILLER_181_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20509_ _09750_ _03404_ _03405_ _03250_ rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1
+ _01399_ sky130_fd_sc_hd__a32o_1
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _05042_ _05054_ _05059_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a21o_1
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21489_ net410 _01258_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14030_ _06762_ _06764_ _06765_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a21o_1
X_11242_ _04004_ _04022_ _04024_ _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__and4b_2
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11173_ rbzero.othery\[2\] _03933_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15981_ _07923_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__clkinv_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17720_ _10195_ _10284_ vssd1 vssd1 vccd1 vccd1 _10285_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14932_ rbzero.wall_tracer.visualWallDist\[2\] _07618_ vssd1 vssd1 vccd1 vccd1 _07631_
+ sky130_fd_sc_hd__or2_1
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20307__320 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__inv_2
X_17651_ _10095_ _10097_ _10093_ vssd1 vssd1 vccd1 vccd1 _10216_ sky130_fd_sc_hd__a21bo_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ rbzero.wall_tracer.stepDistY\[8\] _07579_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07580_ sky130_fd_sc_hd__mux2_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16602_ _07938_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__buf_2
X_13814_ _06423_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__xor2_1
X_17582_ _09994_ _10002_ vssd1 vssd1 vccd1 vccd1 _10148_ sky130_fd_sc_hd__nand2_1
X_14794_ _00004_ _07524_ _07525_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19321_ rbzero.spi_registers.new_vshift\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16533_ _09175_ _09176_ vssd1 vssd1 vccd1 vccd1 _09177_ sky130_fd_sc_hd__xor2_1
X_13745_ _06471_ _06472_ _06481_ _06474_ _06480_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a32o_1
X_10957_ rbzero.tex_b1\[13\] rbzero.tex_b1\[14\] _03817_ vssd1 vssd1 vccd1 vccd1 _03826_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19252_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_sky\[4\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_177_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16464_ _09106_ _09107_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__nor2_1
XFILLER_204_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13676_ _06398_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__xor2_1
XFILLER_143_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ rbzero.tex_b1\[46\] rbzero.tex_b1\[47\] _03784_ vssd1 vssd1 vccd1 vccd1 _03790_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18203_ _01802_ _01803_ _01901_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__and3_1
X_15415_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.side
+ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__mux2_1
X_19183_ rbzero.floor_leak\[2\] _02732_ _02736_ _02722_ vssd1 vssd1 vccd1 vccd1 _00742_
+ sky130_fd_sc_hd__o211a_1
X_12627_ _05380_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__clkbuf_1
X_16395_ _09031_ _09039_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__xnor2_2
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18134_ _01833_ _01834_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__and2_1
X_15346_ _05345_ _05466_ _07893_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__mux2_1
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12558_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] _05300_
+ _05310_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a221o_1
XFILLER_156_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20353__362 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__inv_2
X_11509_ _04210_ _04284_ _04288_ _04242_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a211o_1
XFILLER_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _01764_ _01765_ _01646_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ _07916_ _07921_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__or2_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12489_ rbzero.wall_tracer.trackDistY\[-11\] _05242_ rbzero.wall_tracer.trackDistY\[-12\]
+ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__o211a_1
X_17016_ _09654_ _09655_ vssd1 vssd1 vccd1 vccd1 _09656_ sky130_fd_sc_hd__nand2_1
X_14228_ _06935_ _06963_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__or2_1
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14159_ _06864_ _06895_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__xor2_1
XFILLER_140_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _02613_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _01498_ _01620_ _01618_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18898_ rbzero.spi_registers.spi_counter\[0\] _02564_ _02567_ vssd1 vssd1 vccd1 vccd1
+ _02568_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17849_ _05532_ _01552_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__nand2_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20860_ clknet_leaf_55_i_clk _00629_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19519_ _02983_ _02987_ _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__nand3_1
X_20791_ clknet_leaf_16_i_clk _00560_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21412_ net333 _01181_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21343_ net264 _01112_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21274_ clknet_leaf_63_i_clk _01043_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20181__207 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__inv_2
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ rbzero.tex_g1\[5\] rbzero.tex_g1\[4\] _04336_ vssd1 vssd1 vccd1 vccd1 _04637_
+ sky130_fd_sc_hd__mux2_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _03749_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11791_ rbzero.tex_g0\[55\] _04347_ _04348_ _04217_ vssd1 vssd1 vccd1 vccd1 _04569_
+ sky130_fd_sc_hd__a31o_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20989_ clknet_leaf_50_i_clk _00758_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _06219_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__xor2_1
XFILLER_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10742_ rbzero.tex_g0\[52\] rbzero.tex_g0\[51\] _03706_ vssd1 vssd1 vccd1 vccd1 _03713_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13461_ _06172_ _06187_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__and2b_1
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10673_ rbzero.tex_g1\[20\] rbzero.tex_g1\[21\] _03669_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15200_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__nand2_1
X_12412_ _05146_ _04666_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__nand2_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16180_ _08822_ _08824_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__nand2_1
X_13392_ _06111_ _06128_ _06109_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__a21o_1
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15131_ _07783_ _07784_ _07786_ _07787_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__o211a_1
XFILLER_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12343_ _04323_ _05084_ _05107_ net68 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a22oi_1
XFILLER_166_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12274_ _05032_ net20 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__and2_1
XFILLER_126_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15062_ _07710_ _07714_ _07711_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__o21ai_1
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14013_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__nand2_1
X_11225_ gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__inv_2
XFILLER_107_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19870_ rbzero.debug_overlay.playerX\[3\] _03176_ vssd1 vssd1 vccd1 vccd1 _03180_
+ sky130_fd_sc_hd__nor2_1
XFILLER_136_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03039_ clknet_0__03039_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03039_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18821_ _02499_ _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__xnor2_1
X_11156_ rbzero.debug_overlay.playerX\[4\] rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1
+ vccd1 _03945_ sky130_fd_sc_hd__xor2_1
XFILLER_95_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18752_ _02398_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__buf_4
X_15964_ _08586_ _08608_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__xor2_1
X_11087_ rbzero.tex_b0\[16\] rbzero.tex_b0\[15\] _03887_ vssd1 vssd1 vccd1 vccd1 _03894_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17703_ _10130_ _10266_ _10267_ vssd1 vssd1 vccd1 vccd1 _10268_ sky130_fd_sc_hd__o21a_1
XFILLER_49_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14915_ rbzero.wall_tracer.visualWallDist\[-3\] _07618_ vssd1 vssd1 vccd1 vccd1 _07619_
+ sky130_fd_sc_hd__or2_1
X_18683_ _02235_ _02249_ _02378_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ _08487_ _08506_ _08508_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__and3_1
XFILLER_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _10090_ _10108_ _10198_ vssd1 vssd1 vccd1 vccd1 _10199_ sky130_fd_sc_hd__a21o_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14846_ rbzero.wall_tracer.stepDistY\[4\] _07566_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07567_ sky130_fd_sc_hd__mux2_1
XFILLER_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17565_ _08872_ _08873_ vssd1 vssd1 vccd1 vccd1 _10131_ sky130_fd_sc_hd__nand2_1
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14777_ _07473_ _07507_ _07509_ _05814_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__o211ai_1
XFILLER_189_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11989_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _04212_ vssd1 vssd1 vccd1 vccd1 _04764_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19304_ rbzero.spi_registers.new_other\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_95_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16516_ _09002_ _09019_ _09159_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__a21bo_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ _06436_ _06459_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__xor2_1
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17496_ _10060_ _10061_ vssd1 vssd1 vccd1 vccd1 _10062_ sky130_fd_sc_hd__xor2_1
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19235_ rbzero.spi_registers.new_vshift\[4\] _02763_ vssd1 vssd1 vccd1 vccd1 _02769_
+ sky130_fd_sc_hd__or2_1
XFILLER_177_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16447_ _08961_ _08966_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__nand2_1
X_13659_ _06381_ _06386_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19166_ rbzero.othery\[3\] _02710_ _02724_ _02722_ vssd1 vssd1 vccd1 vccd1 _00737_
+ sky130_fd_sc_hd__o211a_1
X_20277__293 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__inv_2
X_16378_ _08297_ _08326_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__nor2_1
XFILLER_145_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18117_ _01728_ _01729_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__nor2_1
X_15329_ _07970_ _07549_ _07973_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__o21ai_4
X_19097_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.spi_buffer\[3\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_172_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18048_ _01748_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_86_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20010_ _04890_ _04989_ _02703_ _04990_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__or4b_1
XFILLER_141_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19999_ rbzero.pov.ready_buffer\[3\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-6\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__a221o_1
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20912_ clknet_leaf_75_i_clk _00681_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20843_ clknet_leaf_9_i_clk _00612_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20774_ clknet_leaf_37_i_clk _00543_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21326_ net247 _01095_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21257_ clknet_leaf_62_i_clk _01026_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_150_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _03853_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21188_ clknet_leaf_13_i_clk _00957_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ _05697_ _05692_ _05648_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__or3_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _05741_ _07397_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__nand2_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _04271_ vssd1 vssd1 vccd1 vccd1 _04688_
+ sky130_fd_sc_hd__mux2_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15680_ _08298_ _08312_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__nor2_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12892_ rbzero.wall_tracer.visualWallDist\[3\] _04030_ vssd1 vssd1 vccd1 vccd1 _05629_
+ sky130_fd_sc_hd__nor2_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14631_ _07314_ _07367_ _07311_ _07313_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__o211ai_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _04379_ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__or2_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17350_ _09915_ _09916_ vssd1 vssd1 vccd1 vccd1 _09917_ sky130_fd_sc_hd__nor2_2
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _07044_ _07089_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ rbzero.tex_g0\[30\] _04211_ _04125_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a21o_1
XFILLER_207_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _08808_ _08810_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__nor2_1
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13513_ _06248_ _06249_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__nor2_1
X_17281_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09854_ sky130_fd_sc_hd__nor2_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ rbzero.tex_g0\[60\] rbzero.tex_g0\[59\] _03624_ vssd1 vssd1 vccd1 vccd1 _03704_
+ sky130_fd_sc_hd__mux2_1
X_14493_ _07045_ _07046_ _07048_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__a21bo_1
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19020_ _02641_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16232_ _08194_ _08579_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__or2_1
X_13444_ _05910_ _06176_ _06085_ _06180_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a31oi_1
XFILLER_186_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10656_ rbzero.tex_g1\[28\] rbzero.tex_g1\[29\] _03658_ vssd1 vssd1 vccd1 vccd1 _03668_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _08666_ _08668_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__xnor2_4
X_13375_ _06061_ _05940_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10587_ _03631_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15114_ _07758_ _07761_ _07771_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__a21oi_1
X_12326_ _05082_ net28 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__and2_1
XFILLER_127_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16094_ _08695_ _08738_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__xnor2_2
XFILLER_127_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15045_ rbzero.debug_overlay.vplaneX\[-7\] _07705_ vssd1 vssd1 vccd1 vccd1 _07708_
+ sky130_fd_sc_hd__or2_1
X_19922_ rbzero.debug_overlay.playerY\[0\] _03198_ _03219_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00998_ sky130_fd_sc_hd__o211a_1
X_12257_ _05021_ net64 _05024_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a211o_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _03987_ _03996_ _03955_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o21a_1
X_12188_ _04666_ _04903_ _04904_ _04905_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a41o_2
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19853_ rbzero.debug_overlay.playerX\[-1\] _03139_ _03166_ net60 vssd1 vssd1 vccd1
+ vccd1 _00982_ sky130_fd_sc_hd__a211o_1
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18804_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__or2_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11139_ rbzero.debug_overlay.playerX\[1\] _03924_ _03925_ rbzero.debug_overlay.playerY\[0\]
+ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__a221o_1
X_16996_ _09626_ _09635_ vssd1 vssd1 vccd1 vccd1 _09636_ sky130_fd_sc_hd__nand2_1
X_19784_ rbzero.pov.spi_buffer\[65\] rbzero.pov.spi_buffer\[66\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18735_ _09863_ _02424_ _02425_ _09843_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__o31ai_1
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15947_ _07601_ _04014_ _07990_ _07927_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__and4_1
XFILLER_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18666_ _02353_ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _08445_ _08250_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__nand2_1
XFILLER_188_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14829_ _07527_ _07504_ _07449_ _07459_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__o2bb2a_1
X_17617_ _10179_ _10180_ _10175_ _10177_ vssd1 vssd1 vccd1 vccd1 _10182_ sky130_fd_sc_hd__o211a_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18597_ _02169_ _02170_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__or2b_1
XFILLER_205_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17548_ _09117_ _09693_ _09992_ _10113_ vssd1 vssd1 vccd1 vccd1 _10114_ sky130_fd_sc_hd__o31a_1
XFILLER_205_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ _09952_ _10040_ _10044_ vssd1 vssd1 vccd1 vccd1 _10045_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19218_ rbzero.spi_registers.new_floor\[4\] rbzero.color_floor\[4\] _02751_ vssd1
+ vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20490_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03389_
+ sky130_fd_sc_hd__or2_1
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19149_ rbzero.spi_registers.new_other\[7\] _02712_ vssd1 vssd1 vccd1 vccd1 _02715_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21111_ net201 _00880_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21042_ clknet_leaf_77_i_clk _00811_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ clknet_leaf_93_i_clk _00595_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20293__308 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__inv_2
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20757_ clknet_leaf_41_i_clk _00526_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_51_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10510_ _03557_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__clkbuf_4
X_11490_ _04207_ _04233_ _04243_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a31o_1
XFILLER_196_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20688_ clknet_leaf_28_i_clk _00472_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10441_ rbzero.tex_r1\[0\] rbzero.tex_r1\[1\] _03549_ vssd1 vssd1 vccd1 vccd1 _03553_
+ sky130_fd_sc_hd__mux2_1
XFILLER_148_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10372_ rbzero.tex_r1\[33\] rbzero.tex_r1\[34\] _03516_ vssd1 vssd1 vccd1 vccd1 _03517_
+ sky130_fd_sc_hd__mux2_1
X_13160_ _05811_ _05819_ _05814_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a21o_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12111_ gpout0.vpos\[2\] vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__buf_2
XFILLER_151_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13091_ _05826_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__and2_1
X_21309_ net230 _01078_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12042_ _04813_ _04809_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__nor2_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16850_ _09489_ _09490_ vssd1 vssd1 vccd1 vccd1 _09491_ sky130_fd_sc_hd__and2b_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ _08445_ _08227_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__nand2_2
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16781_ _09418_ _09422_ vssd1 vssd1 vccd1 vccd1 _09423_ sky130_fd_sc_hd__and2_1
X_13993_ _06724_ _06690_ _06728_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__o21bai_1
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18520_ _02215_ _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__xnor2_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _08376_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__buf_4
X_12944_ _05678_ _05679_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__mux2_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _02147_ _02148_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__xor2_2
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _08265_ _08307_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__xnor2_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _04030_ _05338_ _05339_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a31o_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17402_ _09967_ _09968_ vssd1 vssd1 vccd1 vccd1 _09969_ sky130_fd_sc_hd__xor2_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14614_ _05793_ _07350_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__and2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11826_ rbzero.tex_g1\[61\] rbzero.tex_g1\[60\] _04392_ vssd1 vssd1 vccd1 vccd1 _04603_
+ sky130_fd_sc_hd__mux2_1
X_18382_ _02070_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__nand2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _08238_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__buf_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _09898_ _09899_ _09900_ _09893_ vssd1 vssd1 vccd1 vccd1 _09901_ sky130_fd_sc_hd__o211ai_1
X_14545_ _07276_ _07280_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__nor2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ rbzero.tex_g0\[2\] _04211_ _04125_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a21o_1
XFILLER_144_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17264_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09839_ sky130_fd_sc_hd__and2_1
X_10708_ _03695_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__clkbuf_1
X_14476_ _07211_ _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nor2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11688_ rbzero.debug_overlay.vplaneX\[-1\] _04465_ _04466_ rbzero.debug_overlay.vplaneX\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a22o_1
XFILLER_186_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19003_ _02632_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16215_ _08858_ _08859_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__xor2_1
X_13427_ _05991_ _05978_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__nor2_1
X_10639_ _03659_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__clkbuf_1
X_17195_ _05413_ vssd1 vssd1 vccd1 vccd1 _09780_ sky130_fd_sc_hd__inv_2
XFILLER_155_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16146_ _08782_ _08783_ _08786_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__or3_1
X_13358_ _05920_ _05975_ _06093_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__or3b_1
X_12309_ _05034_ _05027_ _05069_ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a31o_2
X_16077_ _08008_ _08042_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__nor2_1
X_13289_ _05946_ _05973_ _06007_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or3_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15028_ _07683_ _07691_ _07692_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__a21boi_1
XFILLER_69_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19905_ _07954_ _03141_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nor2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19836_ rbzero.pov.ready_buffer\[63\] _07914_ _03146_ vssd1 vssd1 vccd1 vccd1 _03154_
+ sky130_fd_sc_hd__mux2_1
XFILLER_190_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19767_ rbzero.pov.spi_buffer\[57\] rbzero.pov.spi_buffer\[58\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 i_gpout0_sel[1] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_6
X_16979_ _09537_ _09518_ vssd1 vssd1 vccd1 vccd1 _09619_ sky130_fd_sc_hd__or2b_1
XFILLER_65_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18718_ _02408_ _02409_ _02407_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__o21a_1
XFILLER_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19698_ rbzero.pov.spi_buffer\[24\] rbzero.pov.spi_buffer\[25\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18649_ _02241_ _02245_ _02344_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a21bo_1
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03298_ _03298_ vssd1 vssd1 vccd1 vccd1 clknet_0__03298_ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21660_ clknet_leaf_78_i_clk _01429_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__nand2_1
X_21591_ net132 _01360_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20542_ _03430_ _03431_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__a21o_1
XFILLER_193_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20473_ _03367_ _03369_ _03368_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__a21boi_1
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20136__167 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__inv_2
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21025_ clknet_leaf_66_i_clk _00794_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _03717_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20301__315 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__inv_2
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _05409_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _04387_ _04388_ _04389_ _04226_ _04306_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__o221a_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ clknet_leaf_26_i_clk _00578_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _05337_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__and2_1
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14330_ _07061_ _07066_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__xor2_1
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11542_ gpout0.vpos\[8\] gpout0.vpos\[7\] gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1
+ _04322_ sky130_fd_sc_hd__and3_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14261_ _06997_ _06725_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11473_ _04123_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__buf_4
XFILLER_184_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16000_ _07994_ _08594_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__nor2_1
X_13212_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10424_ rbzero.tex_r1\[8\] rbzero.tex_r1\[9\] _03538_ vssd1 vssd1 vccd1 vccd1 _03544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14192_ _06805_ _06667_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__or3b_1
XFILLER_183_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13143_ _05837_ _05841_ _05807_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__mux2_1
X_10355_ rbzero.tex_r1\[41\] rbzero.tex_r1\[42\] _03505_ vssd1 vssd1 vccd1 vccd1 _03508_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13074_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__clkbuf_2
X_17951_ _01513_ _01533_ _01532_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a21oi_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12025_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _04250_ vssd1 vssd1 vccd1 vccd1 _04800_
+ sky130_fd_sc_hd__mux2_1
X_16902_ _08242_ _09129_ _08283_ vssd1 vssd1 vccd1 vccd1 _09543_ sky130_fd_sc_hd__a21oi_1
X_17882_ _09526_ _09359_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__nor2_1
XFILLER_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16833_ _09379_ _09471_ _09473_ vssd1 vssd1 vccd1 vccd1 _09474_ sky130_fd_sc_hd__a21oi_2
XFILLER_120_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19552_ rbzero.pov.spi_counter\[2\] rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\]
+ _03024_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and4bb_1
X_16764_ _09114_ _08204_ _09271_ vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__or3_1
X_13976_ _05982_ _06663_ _06712_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__or3_1
XFILLER_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ _07931_ _08109_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__nor2_1
X_18503_ _02060_ _02101_ _02058_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12927_ _05660_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__inv_2
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16695_ _09336_ _09337_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19483_ _02905_ _04471_ _02961_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o22ai_1
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15646_ _07912_ _08276_ vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__nor2_1
X_18434_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__and2_1
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ rbzero.wall_tracer.visualWallDist\[-9\] _05355_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__mux2_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _01996_ _01979_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__or2b_1
X_11809_ _04585_ _04586_ _04217_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__mux2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15577_ _07894_ _05494_ vssd1 vssd1 vccd1 vccd1 _08222_ sky130_fd_sc_hd__nand2_1
X_12789_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__buf_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _09863_ _09883_ _09884_ _09885_ vssd1 vssd1 vccd1 vccd1 _09886_ sky130_fd_sc_hd__o31ai_1
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _07261_ _07263_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__nand2_1
X_18296_ _01981_ _01995_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__xor2_1
XFILLER_174_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17247_ _09821_ _09822_ _09823_ vssd1 vssd1 vccd1 vccd1 _09824_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14459_ _07168_ _07183_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__or2b_1
XFILLER_190_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ rbzero.traced_texa\[6\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a22o_1
XFILLER_155_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16129_ _08772_ _08773_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__or2b_1
XFILLER_66_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ _02822_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03319_ clknet_0__03319_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03319_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21643_ clknet_leaf_36_i_clk _01412_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_30 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21574_ net495 _01343_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_41 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20525_ _03411_ _03414_ _03412_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a21boi_1
XFILLER_165_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20456_ _03357_ _03358_ _03359_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a21o_1
XFILLER_107_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21008_ clknet_leaf_52_i_clk _00777_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13830_ _06565_ _06566_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__nand2_1
X_20055__93 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__inv_2
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13761_ _06462_ _06496_ _06426_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a21bo_1
X_10973_ _03834_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15500_ _08137_ _08143_ _08144_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__a21o_1
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12712_ _05439_ _05441_ _05418_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a21bo_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16480_ _09118_ _09123_ vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13692_ _06384_ _06385_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15431_ _08074_ _08075_ _07965_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__or3_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12643_ rbzero.debug_overlay.playerY\[3\] _05393_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_93_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18150_ _01848_ _01849_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and2_1
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15362_ rbzero.wall_tracer.visualWallDist\[-7\] _04014_ _05207_ vssd1 vssd1 vccd1
+ vccd1 _08007_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12574_ _05326_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and2_1
X_17101_ _09082_ _09740_ vssd1 vssd1 vccd1 vccd1 _09741_ sky130_fd_sc_hd__xnor2_1
X_14313_ _07048_ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__nand2_1
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ rbzero.tex_r0\[30\] _04273_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__a21o_1
X_18081_ _01572_ _01659_ _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a21boi_1
X_15293_ _04013_ _07936_ _07937_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__a21oi_4
XFILLER_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17032_ _09545_ _09670_ _09671_ vssd1 vssd1 vccd1 vccd1 _09672_ sky130_fd_sc_hd__a21oi_2
X_14244_ _06946_ _06961_ _06980_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__a21oi_1
X_11456_ _04234_ _04235_ _04226_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__mux2_1
XFILLER_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20119__151 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__inv_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ rbzero.tex_r1\[16\] rbzero.tex_r1\[17\] _03527_ vssd1 vssd1 vccd1 vccd1 _03535_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14175_ _06886_ _06910_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__nand2_1
X_11387_ _04147_ gpout0.hpos\[2\] _04163_ _04164_ _04166_ vssd1 vssd1 vccd1 vccd1
+ _04167_ sky130_fd_sc_hd__a221o_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13126_ _05861_ _05862_ _05807_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__mux2_1
X_10338_ rbzero.tex_r1\[49\] rbzero.tex_r1\[50\] _03494_ vssd1 vssd1 vccd1 vccd1 _03499_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ rbzero.pov.spi_buffer\[24\] rbzero.pov.ready_buffer\[24\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _05700_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__inv_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _08895_ _10139_ _08626_ _09989_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ rbzero.tex_b1\[56\] _04291_ _04139_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a21o_1
XFILLER_113_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17865_ _01566_ _01567_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xnet99_2 clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
X_19604_ clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__buf_1
XFILLER_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16816_ _09341_ _09457_ vssd1 vssd1 vccd1 vccd1 _09458_ sky130_fd_sc_hd__xnor2_4
XFILLER_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17796_ _01497_ _01499_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__nand2_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19535_ _02906_ rbzero.wall_tracer.rayAddendY\[10\] vssd1 vssd1 vccd1 vccd1 _03011_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ _06080_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16747_ _09387_ _09388_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__nand2_1
XFILLER_35_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16678_ _09318_ _09320_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19466_ rbzero.wall_tracer.rayAddendY\[4\] _00013_ _02947_ vssd1 vssd1 vccd1 vccd1
+ _00814_ sky130_fd_sc_hd__o21a_1
XFILLER_179_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18417_ _02105_ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__xnor2_1
X_15629_ _05193_ _08273_ _04013_ vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__o21a_1
X_19397_ _02865_ _02875_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nand2_1
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18348_ _10266_ _02045_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__o21ba_1
XFILLER_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18279_ _01865_ _01873_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a21o_1
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21290_ clknet_leaf_42_i_clk _01059_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[8\] sky130_fd_sc_hd__dfxtp_1
Xinput50 i_vec_csb vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_6
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20330__341 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__inv_2
XFILLER_118_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20172_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__buf_1
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20248__268 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__inv_2
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19588__44 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21626_ clknet_leaf_20_i_clk _01395_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21557_ net478 _01326_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11310_ _04071_ _04074_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__and2_1
XFILLER_166_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20508_ _03401_ _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nand3_1
X_12290_ _05055_ _05056_ _05057_ _05058_ _05033_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__o311a_1
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21488_ net409 _01257_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11241_ _03475_ _04006_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nor2_1
XFILLER_175_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20439_ _03343_ _03344_ _03345_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__or3_1
XFILLER_162_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11172_ rbzero.otherx\[4\] rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 _03961_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_175_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15980_ _07912_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__or3_1
XFILLER_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14931_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.trackDistX\[2\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14862_ _07456_ _07577_ _07578_ _07487_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__o31a_4
X_17650_ _10073_ _10077_ _10075_ vssd1 vssd1 vccd1 vccd1 _10215_ sky130_fd_sc_hd__a21bo_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ _06426_ _06462_ _06422_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__o21bai_1
X_16601_ _07932_ _07938_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__or4_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17581_ _10122_ _10146_ vssd1 vssd1 vccd1 vccd1 _10147_ sky130_fd_sc_hd__xnor2_2
X_14793_ rbzero.wall_tracer.stepDistY\[-7\] _00004_ vssd1 vssd1 vccd1 vccd1 _07525_
+ sky130_fd_sc_hd__nor2_1
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19320_ _02816_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16532_ _09031_ _09039_ _09037_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__a21oi_1
XFILLER_182_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ _06474_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__xor2_1
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10956_ _03825_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19251_ _02778_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__clkbuf_1
X_16463_ _09102_ _09105_ vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__and2_1
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13675_ _06405_ _06410_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o21ba_1
X_10887_ _03789_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18202_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__inv_2
X_15414_ _08058_ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__buf_2
X_19182_ rbzero.spi_registers.new_leak\[2\] _02733_ vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__or2_1
X_12626_ _05379_ _03942_ _05284_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__mux2_1
X_16394_ _09037_ _09038_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__nor2_1
XFILLER_169_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18133_ _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__nand2_1
X_15345_ _05196_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__buf_4
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12557_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\]
+ rbzero.debug_overlay.facingY\[-3\] vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__o211a_1
XFILLER_157_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11508_ _04285_ _04286_ _04287_ _04226_ _04230_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__o221a_1
X_18064_ _01646_ _01764_ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and3_1
XFILLER_172_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ _07920_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__inv_2
X_12488_ rbzero.wall_tracer.trackDistX\[-12\] vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__inv_2
XFILLER_89_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17015_ _09618_ _09619_ _09653_ vssd1 vssd1 vccd1 vccd1 _09655_ sky130_fd_sc_hd__nand3_1
X_14227_ _06935_ _06963_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__nand2_1
XFILLER_160_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _04218_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__buf_4
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14158_ _06776_ _06677_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nor2_1
XFILLER_152_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _05835_ _05845_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nor2_4
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14089_ _06806_ _06808_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__xnor2_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ rbzero.pov.spi_buffer\[16\] rbzero.pov.ready_buffer\[16\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17917_ _08057_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__buf_2
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18897_ rbzero.spi_registers.spi_counter\[6\] rbzero.spi_registers.spi_counter\[5\]
+ rbzero.spi_registers.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__or3_1
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17848_ _01550_ _01551_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__xnor2_4
XFILLER_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17779_ _01473_ _01481_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or2_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19518_ rbzero.debug_overlay.vplaneY\[0\] _02980_ _02993_ _02995_ vssd1 vssd1 vccd1
+ vccd1 _02996_ sky130_fd_sc_hd__o22a_1
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20790_ clknet_leaf_21_i_clk _00559_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19449_ _02930_ _02931_ _02911_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__o21bai_1
XFILLER_195_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21411_ net332 _01180_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21342_ net263 _01111_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21273_ clknet_leaf_63_i_clk _01042_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_116_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ rbzero.tex_g0\[20\] rbzero.tex_g0\[19\] _03740_ vssd1 vssd1 vccd1 vccd1 _03749_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ rbzero.tex_g0\[54\] _04350_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__and2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ clknet_leaf_49_i_clk _00757_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _03712_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13460_ _06170_ _06171_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2b_1
XFILLER_158_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10672_ _03676_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _05150_ _05138_ _05152_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a31o_2
X_21609_ net126 _01378_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[60\] sky130_fd_sc_hd__dfxtp_1
X_13391_ _06126_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__nor2_1
XFILLER_182_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15130_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__or2_1
XFILLER_194_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12342_ _05101_ _05105_ _05109_ net28 vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__o22a_1
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _07721_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__nand2_1
X_12273_ net23 _05033_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__nor2_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14012_ _06746_ _06747_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__or2_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11224_ _04010_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_6
XFILLER_181_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03038_ clknet_0__03038_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03038_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18820_ _02492_ _02494_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__or2_1
XFILLER_150_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11155_ rbzero.debug_overlay.playerY\[1\] _03942_ vssd1 vssd1 vccd1 vccd1 _03944_
+ sky130_fd_sc_hd__or2_1
XFILLER_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18751_ _09863_ _02438_ _02439_ _09860_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o31ai_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15963_ _08605_ _08606_ _08607_ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__a21oi_1
X_11086_ _03893_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17702_ _10139_ _08873_ _08263_ _10134_ vssd1 vssd1 vccd1 vccd1 _10267_ sky130_fd_sc_hd__a2bb2o_1
X_14914_ _07594_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__clkbuf_2
X_15894_ _08512_ _08538_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__xor2_1
X_18682_ _02250_ _02287_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__and2b_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _10092_ _10107_ vssd1 vssd1 vccd1 vccd1 _10198_ sky130_fd_sc_hd__nor2_1
X_14845_ _05929_ _07456_ _07458_ _07487_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__o31a_2
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14776_ _07477_ _07475_ _07508_ _05884_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__a211o_1
X_17564_ _08872_ _08873_ _10129_ vssd1 vssd1 vccd1 vccd1 _10130_ sky130_fd_sc_hd__or3_1
X_11988_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _04212_ vssd1 vssd1 vccd1 vccd1 _04763_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19303_ _02807_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__clkbuf_1
X_13727_ _06423_ _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__nand2_1
XFILLER_182_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16515_ _09020_ _09000_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__or2b_1
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10939_ _03816_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17495_ _09096_ _09217_ vssd1 vssd1 vccd1 vccd1 _10061_ sky130_fd_sc_hd__nor2_1
XFILLER_149_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19234_ rbzero.spi_registers.vshift\[3\] _02762_ _02768_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00761_ sky130_fd_sc_hd__o211a_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13658_ _06352_ _06367_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__xnor2_1
X_16446_ _09008_ _09018_ _09016_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__a21o_1
XFILLER_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _05318_ _05308_ _05312_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__or3_1
X_16377_ _08998_ _09021_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19165_ rbzero.spi_registers.new_other\[3\] _02712_ vssd1 vssd1 vccd1 vccd1 _02724_
+ sky130_fd_sc_hd__or2_1
X_13589_ _06325_ _06301_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18116_ _01691_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__xnor2_1
X_15328_ _07971_ _05340_ _07972_ _05193_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__a211o_1
XFILLER_184_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19096_ _02681_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15259_ _07903_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__buf_4
X_18047_ _01503_ _01623_ _01624_ _01625_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19998_ rbzero.pov.ready_buffer\[2\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[-7\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__o221a_1
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18949_ rbzero.pov.spi_buffer\[8\] rbzero.pov.ready_buffer\[8\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20911_ clknet_leaf_75_i_clk _00680_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ clknet_leaf_8_i_clk _00611_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20773_ clknet_leaf_36_i_clk _00542_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21325_ net246 _01094_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21256_ clknet_leaf_81_i_clk _01025_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21187_ clknet_leaf_13_i_clk _00956_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20138_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__buf_1
XFILLER_89_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _05615_ _05639_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _04271_ vssd1 vssd1 vccd1 vccd1 _04687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__buf_2
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _07306_ _07307_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__and2_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ rbzero.tex_g1\[33\] rbzero.tex_g1\[32\] _04337_ vssd1 vssd1 vccd1 vccd1 _04619_
+ sky130_fd_sc_hd__mux2_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _07086_ _07088_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__nor2_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11773_ rbzero.tex_g0\[31\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__and3_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _06237_ _06238_ _06247_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__and3_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16300_ _08620_ _08670_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__xnor2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17280_ _09853_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__clkbuf_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _03703_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__clkbuf_1
X_14492_ _07165_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16231_ _08867_ _08875_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__nand2_1
X_13443_ _06041_ _06080_ _06084_ _05990_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__o22a_1
XFILLER_139_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10655_ _03667_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16162_ _08801_ _08805_ _08806_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__a21oi_4
XFILLER_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _06109_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__nor2_1
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10586_ rbzero.tex_g1\[61\] rbzero.tex_g1\[62\] _03549_ vssd1 vssd1 vccd1 vccd1 _03631_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15113_ _07769_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__nand2_1
X_12325_ _05087_ net64 _05091_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a211o_1
XFILLER_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16093_ _08716_ _08715_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__and2b_1
XFILLER_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15044_ rbzero.wall_tracer.rayAddendX\[-4\] _00013_ _07702_ _07707_ vssd1 vssd1 vccd1
+ vccd1 _00492_ sky130_fd_sc_hd__o22a_1
X_19921_ rbzero.pov.ready_buffer\[53\] _03141_ _03192_ _03218_ vssd1 vssd1 vccd1 vccd1
+ _03219_ sky130_fd_sc_hd__a211o_1
X_12256_ _05021_ _04738_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__nor2_1
XFILLER_141_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11207_ _03993_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__nand2_2
X_19852_ _08093_ _03164_ _03143_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a211oi_1
X_12187_ _04907_ _04908_ net13 _04917_ _04957_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__o41a_2
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _02485_ _10028_ rbzero.wall_tracer.trackDistY\[0\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00613_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ rbzero.debug_overlay.playerY\[3\] _03921_ _03926_ rbzero.map_rom.f3 vssd1
+ vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19783_ _03120_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16995_ _09633_ _09634_ vssd1 vssd1 vccd1 vccd1 _09635_ sky130_fd_sc_hd__and2_1
XFILLER_62_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18734_ _02421_ _02422_ _02423_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__o21a_1
XFILLER_37_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11069_ _03884_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15946_ rbzero.wall_tracer.visualWallDist\[-11\] _04014_ _05197_ _07992_ vssd1 vssd1
+ vccd1 vccd1 _08591_ sky130_fd_sc_hd__and4_1
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18665_ _02359_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__xnor2_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15877_ _08520_ _08521_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__xnor2_2
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17616_ _10175_ _10177_ _10179_ _10180_ vssd1 vssd1 vccd1 vccd1 _10181_ sky130_fd_sc_hd__a211oi_1
X_14828_ _00004_ _07552_ _07553_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18596_ _02166_ _02197_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a21bo_1
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17547_ _08873_ _09991_ _09696_ vssd1 vssd1 vccd1 vccd1 _10113_ sky130_fd_sc_hd__or3b_1
X_14759_ _07357_ _07370_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__and2b_1
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17478_ _10042_ _10043_ vssd1 vssd1 vccd1 vccd1 _10044_ sky130_fd_sc_hd__or2_1
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19217_ rbzero.color_floor\[3\] _02751_ _02757_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__a21o_1
X_16429_ _09068_ _09072_ _09073_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__a21o_1
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19148_ rbzero.otherx\[0\] _02710_ _02713_ _02714_ vssd1 vssd1 vccd1 vccd1 _00729_
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19079_ rbzero.pov.spi_buffer\[70\] rbzero.pov.ready_buffer\[70\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21110_ net200 _00879_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21041_ clknet_leaf_77_i_clk _00810_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20389__15 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20825_ clknet_leaf_0_i_clk _00594_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20756_ clknet_leaf_38_i_clk _00525_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20687_ clknet_3_5_0_i_clk _00471_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ _03552_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _03482_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12110_ _04869_ _04879_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__nor2_1
XFILLER_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21308_ net229 _01077_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _05591_ _05803_ _05796_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__mux2_1
XFILLER_152_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12041_ _04317_ _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__or2_1
X_21239_ clknet_leaf_80_i_clk _01008_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20113__146 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__inv_2
XFILLER_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15800_ _07904_ rbzero.wall_tracer.stepDistY\[-1\] _08272_ _08274_ vssd1 vssd1 vccd1
+ vccd1 _08445_ sky130_fd_sc_hd__a22o_4
Xclkbuf_leaf_70_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13992_ _06724_ _06610_ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__or3b_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16780_ _09419_ _09421_ vssd1 vssd1 vccd1 vccd1 _09422_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12943_ _05601_ _05638_ _05649_ _05628_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__o31a_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _05206_ _08215_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__or2_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _08356_ _09138_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__nor2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ rbzero.wall_tracer.visualWallDist\[-2\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05611_ sky130_fd_sc_hd__a21o_1
X_15662_ _08276_ _07989_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__nor2_1
XFILLER_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_85_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17401_ _09545_ _09670_ _09672_ _09669_ vssd1 vssd1 vccd1 vccd1 _09968_ sky130_fd_sc_hd__a22oi_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _07284_ _07321_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__xor2_1
X_11825_ rbzero.tex_g1\[63\] rbzero.tex_g1\[62\] _04337_ vssd1 vssd1 vccd1 vccd1 _04602_
+ sky130_fd_sc_hd__mux2_1
X_18381_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__and2_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ rbzero.wall_tracer.visualWallDist\[-12\] _04014_ vssd1 vssd1 vccd1 vccd1
+ _08238_ sky130_fd_sc_hd__nand2_2
XFILLER_187_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14544_ _07276_ _07280_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__and2_1
XFILLER_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09900_ sky130_fd_sc_hd__nand2_1
XFILLER_159_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11756_ rbzero.tex_g0\[3\] _04088_ _04127_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__and3_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ rbzero.tex_g1\[4\] rbzero.tex_g1\[5\] _03691_ vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__mux2_1
X_14475_ _07144_ _07156_ _07158_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__o21ba_1
X_17263_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09838_ sky130_fd_sc_hd__nor2_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11687_ _04437_ _04447_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__and2_2
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19002_ rbzero.pov.spi_buffer\[33\] rbzero.pov.ready_buffer\[33\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
X_13426_ _06160_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__xor2_1
XFILLER_186_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16214_ _08816_ _08823_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__nor2_1
XFILLER_179_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10638_ rbzero.tex_g1\[37\] rbzero.tex_g1\[38\] _03658_ vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__mux2_1
X_17194_ _04019_ _05412_ vssd1 vssd1 vccd1 vccd1 _09779_ sky130_fd_sc_hd__nor2_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16145_ _08768_ _08789_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__xnor2_1
X_13357_ _05991_ _05975_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__o21bai_1
XFILLER_154_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10569_ rbzero.tex_r0\[6\] rbzero.tex_r0\[5\] _03613_ vssd1 vssd1 vccd1 vccd1 _03622_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12308_ _05072_ _05074_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and3_1
XFILLER_143_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16076_ _08675_ _08720_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__xor2_1
X_13288_ _05983_ _06016_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__nor2_1
XFILLER_142_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15027_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__nand2_1
X_19904_ rbzero.debug_overlay.playerY\[-5\] _03198_ _03206_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00993_ sky130_fd_sc_hd__o211a_1
XFILLER_190_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12239_ _05004_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__nand2_1
XFILLER_190_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19835_ _03139_ _03152_ _03153_ _02765_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__o211a_1
X_20088__123 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__inv_2
XFILLER_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19766_ _03111_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16978_ _09536_ _09520_ vssd1 vssd1 vccd1 vccd1 _09618_ sky130_fd_sc_hd__or2b_1
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 i_gpout0_sel[2] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18717_ _02407_ _02408_ _02409_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__nor3_1
XFILLER_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15929_ _08124_ _08490_ _08084_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__a21oi_1
X_19697_ _03075_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18648_ _02045_ _02150_ _02152_ _02243_ _02343_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a311o_1
Xclkbuf_0__03297_ _03297_ vssd1 vssd1 vccd1 vccd1 clknet_0__03297_ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18579_ _01860_ _08423_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__nor2_1
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20610_ gpout4.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__nor2_1
XFILLER_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21590_ net131 _01359_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20541_ _03424_ _03428_ _03425_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20472_ _03372_ _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__or2_1
XFILLER_119_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21024_ clknet_leaf_65_i_clk _00793_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11610_ rbzero.tex_r1\[53\] rbzero.tex_r1\[52\] _04338_ vssd1 vssd1 vccd1 vccd1 _04389_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20808_ clknet_leaf_27_i_clk _00577_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12590_ _05309_ _05343_ _05305_ _05299_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a211o_1
XFILLER_204_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ gpout0.vpos\[3\] _04315_ _04316_ gpout0.vpos\[4\] _04320_ vssd1 vssd1 vccd1
+ vccd1 _04321_ sky130_fd_sc_hd__o221ai_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20739_ clknet_leaf_14_i_clk _00508_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ _06134_ _06667_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__or2_1
X_11472_ _04225_ _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__or2_1
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13211_ _05946_ _05947_ _05888_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__or3_1
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10423_ _03543_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_1
X_14191_ _06895_ _06925_ _06927_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13142_ _05830_ _05878_ _05778_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__mux2_1
X_10354_ _03507_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13073_ _05797_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and2_1
X_17950_ _01632_ _01652_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__xnor2_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12024_ _04266_ _04798_ _04229_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__o21a_1
X_16901_ _09541_ vssd1 vssd1 vccd1 vccd1 _09542_ sky130_fd_sc_hd__inv_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17881_ _01581_ _01583_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nand2_1
XFILLER_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16832_ _09358_ _09360_ _09472_ vssd1 vssd1 vccd1 vccd1 _09473_ sky130_fd_sc_hd__o21a_1
XFILLER_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19551_ rbzero.pov.spi_counter\[5\] rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\]
+ rbzero.pov.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__and4bb_1
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16763_ _09383_ _09404_ vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__xnor2_1
X_13975_ _06659_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18502_ _02163_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _07940_ _08084_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__nor2_1
XFILLER_206_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12926_ _05574_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19482_ _02905_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _02962_
+ sky130_fd_sc_hd__and2_1
XFILLER_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16694_ _09198_ _09200_ _09197_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__a21o_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18433_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__nor2_1
XFILLER_59_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _07977_ _07923_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__nor2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12857_ _05589_ _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or3_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18364_ _01995_ _01981_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__or2b_1
X_11808_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _04341_ vssd1 vssd1 vccd1 vccd1 _04586_
+ sky130_fd_sc_hd__mux2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _04016_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__buf_4
X_15576_ _07566_ _08220_ _07970_ vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17315_ _09807_ _09458_ vssd1 vssd1 vccd1 vccd1 _09885_ sky130_fd_sc_hd__or2_1
X_14527_ _07261_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__nor2_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11739_ _04320_ _04508_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__and3_1
X_18295_ _01987_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17246_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ _09815_ vssd1 vssd1 vccd1 vccd1 _09823_ sky130_fd_sc_hd__a21o_1
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14458_ _07162_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13409_ _06139_ _06140_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nand2_1
X_14389_ _06698_ _07121_ _06760_ _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o31a_1
X_17177_ rbzero.traced_texa\[5\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a22o_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16128_ _08728_ _08731_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16059_ _08702_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xor2_1
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19818_ rbzero.debug_overlay.playerX\[-9\] vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__inv_2
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03318_ clknet_0__03318_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03318_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19749_ _03102_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21642_ clknet_leaf_36_i_clk _01411_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20142__172 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__inv_2
XFILLER_52_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21573_ net494 _01342_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_20 _09331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_42 _01673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ _03416_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__and2b_1
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20455_ _03357_ _03358_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nand3_1
XFILLER_119_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21007_ clknet_leaf_50_i_clk _00776_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _06426_ _06462_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__nand3b_1
X_10972_ rbzero.tex_b1\[6\] rbzero.tex_b1\[7\] _03828_ vssd1 vssd1 vccd1 vccd1 _03834_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20225__247 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__inv_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12711_ _05457_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__xnor2_2
X_13691_ _05824_ _06134_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__or2_1
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15430_ _07964_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12642_ _05203_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__buf_4
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _08002_ _08005_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__nand2_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[11\] vssd1
+ vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__or2_1
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17100_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerX\[-1\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09740_ sky130_fd_sc_hd__mux2_1
XFILLER_196_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14312_ _06724_ _06678_ _07047_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__o21bai_1
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11524_ _04217_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__buf_6
X_15292_ _07903_ rbzero.wall_tracer.stepDistY\[-5\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _07937_ sky130_fd_sc_hd__a21o_1
X_18080_ _01658_ _01656_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__or2b_1
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14243_ _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__xor2_1
X_17031_ _07959_ _09276_ _08111_ _09126_ vssd1 vssd1 vccd1 vccd1 _09671_ sky130_fd_sc_hd__o22a_1
X_11455_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _04214_ vssd1 vssd1 vccd1 vccd1 _04235_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10406_ _03534_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
X_14174_ _06886_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__or2_1
X_11386_ _04164_ gpout0.hpos\[1\] gpout0.hpos\[0\] _04165_ vssd1 vssd1 vccd1 vccd1
+ _04166_ sky130_fd_sc_hd__o211a_1
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13125_ _05728_ _05744_ _05791_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__mux2_1
X_10337_ _03498_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18982_ _02621_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13056_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__clkbuf_4
X_17933_ _08767_ _10139_ _01518_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__or3b_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ rbzero.tex_b1\[57\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__and3_1
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17864_ _01563_ _01565_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__or2_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16815_ _09342_ _09456_ vssd1 vssd1 vccd1 vccd1 _09457_ sky130_fd_sc_hd__xor2_4
XFILLER_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xnet99_3 clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
X_17795_ _09276_ _08493_ _08044_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__o22ai_1
X_19534_ _02906_ rbzero.wall_tracer.rayAddendY\[9\] _03003_ vssd1 vssd1 vccd1 vccd1
+ _03010_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16746_ _07996_ _08129_ _08047_ _08705_ vssd1 vssd1 vccd1 vccd1 _09388_ sky130_fd_sc_hd__o22ai_1
X_13958_ _06687_ _06694_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__or2_1
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12909_ _05610_ _05612_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nand2_2
X_19465_ _04035_ _02936_ _02937_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a31o_1
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677_ _09156_ _09182_ _09319_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13889_ _06621_ _06625_ _06576_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__o21a_1
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18416_ _01922_ _02114_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _05364_ _05461_ _07893_ vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__mux2_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19396_ _02878_ _02881_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18347_ _08802_ _01524_ _10139_ _09668_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__o22a_1
XFILLER_187_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15559_ _08202_ _08203_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__and2_2
XFILLER_174_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _01870_ _01872_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__nor2_1
XFILLER_163_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17229_ _09804_ _09805_ _09806_ _09807_ vssd1 vssd1 vccd1 vccd1 _09808_ sky130_fd_sc_hd__a211o_1
Xinput40 i_mode[2] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_4
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput51 i_vec_mosi vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_4
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21625_ clknet_leaf_20_i_clk _01394_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21556_ net477 _01325_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[7\] sky130_fd_sc_hd__dfxtp_1
X_20507_ _03401_ _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a21o_1
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21487_ net408 _01256_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ gpout0.hpos\[3\] _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__and2_1
XFILLER_140_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20438_ _03343_ _03344_ _03345_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o21ai_1
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11171_ rbzero.otherx\[2\] _03929_ rbzero.map_rom.a6 _03958_ _03959_ vssd1 vssd1
+ vccd1 vccd1 _03960_ sky130_fd_sc_hd__o221a_1
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14930_ _07621_ _07628_ _07629_ _07620_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__o211a_1
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _05902_ _07426_ _07394_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__o21ai_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _08075_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__buf_2
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _06426_ _06496_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nor2_1
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17580_ _10124_ _10145_ vssd1 vssd1 vccd1 vccd1 _10146_ sky130_fd_sc_hd__xnor2_2
XFILLER_91_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _07487_ _07456_ _07522_ _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__a211oi_4
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16531_ _09167_ _09174_ vssd1 vssd1 vccd1 vccd1 _09175_ sky130_fd_sc_hd__xnor2_1
X_13743_ _06475_ _06476_ _06477_ _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__a22o_1
X_10955_ rbzero.tex_b1\[14\] rbzero.tex_b1\[15\] _03817_ vssd1 vssd1 vccd1 vccd1 _03825_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19250_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_sky\[3\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16462_ _09102_ _09105_ vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__nor2_1
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13674_ _06400_ _06404_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__nor2_1
XFILLER_143_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10886_ rbzero.tex_b1\[47\] rbzero.tex_b1\[48\] _03784_ vssd1 vssd1 vccd1 vccd1 _03789_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18201_ _01802_ _01803_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a21o_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ _05209_ _08057_ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__or2_2
XFILLER_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19181_ rbzero.floor_leak\[1\] _02732_ _02735_ _02722_ vssd1 vssd1 vccd1 vccd1 _00741_
+ sky130_fd_sc_hd__o211a_1
X_12625_ rbzero.debug_overlay.playerY\[1\] _05378_ _05204_ vssd1 vssd1 vccd1 vccd1
+ _05379_ sky130_fd_sc_hd__mux2_1
X_16393_ _08352_ _08355_ _09036_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__and3_1
XFILLER_145_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18132_ _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__or2_1
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15344_ _07988_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__clkbuf_4
X_12556_ _05301_ _05305_ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__o21a_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _04273_ vssd1 vssd1 vccd1 vccd1 _04287_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18063_ _01762_ _01763_ _01755_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a21o_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12487_ rbzero.wall_tracer.trackDistX\[-11\] vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__inv_2
XFILLER_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15275_ _07903_ _07918_ _07919_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__a21o_1
XFILLER_184_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17014_ _09618_ _09619_ _09653_ vssd1 vssd1 vccd1 vccd1 _09654_ sky130_fd_sc_hd__a21o_1
X_14226_ _06805_ _06672_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__nor2_1
X_11438_ _04217_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__buf_6
XFILLER_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14157_ _06805_ _06663_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nor2_1
X_11369_ _04147_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nand2_1
XFILLER_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13108_ _05814_ _05840_ _05843_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a22o_1
XFILLER_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14088_ _06669_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__xnor2_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ _02612_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__clkbuf_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _05759_ _05772_ _05775_ _05699_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__or4b_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17916_ _01498_ _08057_ _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__or3_1
XFILLER_113_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18896_ rbzero.spi_registers.spi_counter\[2\] _02565_ vssd1 vssd1 vccd1 vccd1 _02566_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_117_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17847_ _10292_ _10295_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__nor2_2
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20208__231 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__inv_2
X_17778_ _01473_ _01481_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__and2_1
XFILLER_47_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19517_ _02980_ _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nand2_1
X_16729_ _09364_ _09370_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19448_ _02913_ _02916_ _02929_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__and3_1
XFILLER_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ _04034_ _02864_ _02865_ _02866_ _07706_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a221o_1
XFILLER_210_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21410_ net331 _01179_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21341_ net262 _01110_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21272_ clknet_leaf_65_i_clk _01041_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
X_20254__273 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__inv_2
XFILLER_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20987_ clknet_leaf_48_i_clk _00756_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10740_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _03706_ vssd1 vssd1 vccd1 vccd1 _03712_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10671_ rbzero.tex_g1\[21\] rbzero.tex_g1\[22\] _03669_ vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ net36 _05165_ _05176_ net37 vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o211a_1
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21608_ net149 _01377_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _06124_ _06125_ _06121_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a21oi_1
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20337__348 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__inv_2
XFILLER_167_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _05100_ _05106_ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o21ai_1
X_21539_ net460 _01308_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15060_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__nand2_1
X_12272_ _05035_ _05040_ net25 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__and3b_1
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14011_ _06746_ _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__nand2_1
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11223_ _04007_ _04008_ _04009_ _03477_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or4b_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03037_ clknet_0__03037_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03037_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ rbzero.debug_overlay.playerY\[1\] _03942_ vssd1 vssd1 vccd1 vccd1 _03943_
+ sky130_fd_sc_hd__nand2_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18750_ _02435_ _02436_ _02437_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__o21a_1
X_15962_ _08587_ _08604_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__nor2_1
X_11085_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _03887_ vssd1 vssd1 vccd1 vccd1 _03893_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17701_ _10139_ vssd1 vssd1 vccd1 vccd1 _10266_ sky130_fd_sc_hd__clkbuf_4
X_14913_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.trackDistX\[-3\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__mux2_1
X_18681_ _02293_ _02298_ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a21o_1
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _08535_ _08536_ _08537_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _10069_ _10083_ _10196_ vssd1 vssd1 vccd1 vccd1 _10197_ sky130_fd_sc_hd__a21o_1
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14844_ _07565_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__clkbuf_1
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20082__118 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__inv_2
XFILLER_64_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17563_ _05211_ _09699_ _10128_ vssd1 vssd1 vccd1 vccd1 _10129_ sky130_fd_sc_hd__o21a_1
X_14775_ _07477_ _07479_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__nor2_1
X_11987_ _04247_ _04759_ _04760_ _04761_ _04254_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__o221a_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19302_ rbzero.spi_registers.new_other\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16514_ _09040_ _08430_ _09041_ _09157_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__o31ai_2
XFILLER_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13726_ _06426_ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__nor2_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10938_ rbzero.tex_b1\[22\] rbzero.tex_b1\[23\] _03806_ vssd1 vssd1 vccd1 vccd1 _03816_
+ sky130_fd_sc_hd__mux2_1
X_17494_ _10058_ _10059_ vssd1 vssd1 vccd1 vccd1 _10060_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19233_ rbzero.spi_registers.new_vshift\[3\] _02763_ vssd1 vssd1 vccd1 vccd1 _02768_
+ sky130_fd_sc_hd__or2_1
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16445_ _09056_ _09058_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__nand2_1
X_13657_ _06388_ _06390_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__xnor2_1
X_10869_ rbzero.tex_b1\[55\] rbzero.tex_b1\[56\] _03773_ vssd1 vssd1 vccd1 vccd1 _03780_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _05308_ _05312_ _05318_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__o21ai_1
X_19164_ rbzero.othery\[2\] _02710_ _02723_ _02722_ vssd1 vssd1 vccd1 vccd1 _00736_
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _09000_ _09020_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__xnor2_2
X_13588_ _06281_ _06283_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__nor2_1
XFILLER_185_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18115_ _01814_ _01815_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__nor2_1
XFILLER_157_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15327_ _07971_ _05488_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__nor2_1
X_19095_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.spi_buffer\[2\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
X_12539_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] _05291_
+ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a31o_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18046_ _01746_ _01747_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__xor2_1
XFILLER_145_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14209_ _06932_ _06945_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__or2b_1
XFILLER_144_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15189_ rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\] rbzero.wall_tracer.rayAddendX\[4\]
+ rbzero.wall_tracer.rayAddendX\[3\] _07785_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__o41a_1
XFILLER_193_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19997_ rbzero.pov.ready_buffer\[1\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[-8\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__o221a_1
XFILLER_154_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18948_ _02603_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18879_ rbzero.wall_tracer.trackDistY\[11\] rbzero.wall_tracer.stepDistY\[11\] vssd1
+ vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__xor2_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20910_ clknet_leaf_79_i_clk _00679_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_20284__299 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__inv_2
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20841_ clknet_leaf_8_i_clk _00610_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20772_ clknet_leaf_35_i_clk _00541_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21324_ net245 _01093_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21255_ clknet_leaf_81_i_clk _01024_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21186_ clknet_leaf_13_i_clk _00955_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _04684_ _04685_ _04265_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__mux2_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _05562_ _05565_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and2_1
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _04230_ _04613_ _04617_ _04232_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a211o_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14560_ _07291_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__nand2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _04129_ vssd1 vssd1 vccd1 vccd1 _04550_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _06237_ _06238_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _03624_ vssd1 vssd1 vccd1 vccd1 _03703_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14491_ _07137_ _07045_ _07166_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__a21o_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16230_ _08871_ _08874_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__nor2_1
X_13442_ _06078_ _06067_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__or2_1
XFILLER_186_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ rbzero.tex_g1\[29\] rbzero.tex_g1\[30\] _03658_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ _06037_ _06092_ _06108_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ _08737_ _08761_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__xnor2_2
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10585_ _03630_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__or2_1
X_12324_ _05087_ _04738_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__nor2_1
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16092_ _08725_ _08734_ _08736_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__a21oi_4
XFILLER_115_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ net23 net24 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__nand2_1
X_15043_ _07703_ _07704_ _07705_ _07706_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__a31o_1
X_19920_ _03216_ _03217_ _02822_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11206_ _03933_ rbzero.map_rom.i_row\[4\] _03990_ _03994_ vssd1 vssd1 vccd1 vccd1
+ _03995_ sky130_fd_sc_hd__or4_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19851_ rbzero.pov.ready_buffer\[67\] _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__nor2_1
X_12186_ _04904_ _04925_ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a21oi_2
XFILLER_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18802_ _05532_ _02483_ _02484_ _02399_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__o31a_1
X_11137_ rbzero.debug_overlay.playerX\[1\] vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__inv_2
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19782_ rbzero.pov.spi_buffer\[64\] rbzero.pov.spi_buffer\[65\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
XFILLER_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16994_ _09631_ _09632_ vssd1 vssd1 vccd1 vccd1 _09634_ sky130_fd_sc_hd__nand2_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18733_ _02421_ _02422_ _02423_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__nor3_1
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11068_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _03876_ vssd1 vssd1 vccd1 vccd1 _03884_
+ sky130_fd_sc_hd__mux2_1
X_15945_ _08522_ _08523_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__xnor2_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18664_ _08257_ _09215_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__nor2_1
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15876_ _07601_ _04014_ _05197_ _07992_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__and4_1
XFILLER_209_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _10180_ sky130_fd_sc_hd__nor2_1
X_14827_ rbzero.wall_tracer.stepDistY\[-1\] _07461_ vssd1 vssd1 vccd1 vccd1 _07553_
+ sky130_fd_sc_hd__nor2_1
X_18595_ _02198_ _02164_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__or2b_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17546_ _09686_ _09980_ _10111_ vssd1 vssd1 vccd1 vccd1 _10112_ sky130_fd_sc_hd__a21bo_1
X_14758_ _07477_ _07489_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__a21oi_1
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__or2_1
X_17477_ _09933_ _09936_ _10041_ vssd1 vssd1 vccd1 vccd1 _10043_ sky130_fd_sc_hd__and3_1
X_14689_ _07106_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__or2_1
X_19216_ rbzero.spi_registers.new_floor\[3\] rbzero.spi_registers.got_new_floor _02711_
+ _03911_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a31o_1
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16428_ _09071_ _09069_ _09070_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__and3_1
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19147_ _05190_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__buf_2
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16359_ _07967_ _08035_ _08046_ _08674_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__o22ai_1
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19078_ _02671_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18029_ _01715_ _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21040_ clknet_leaf_77_i_clk _00809_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20366__374 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__inv_2
XFILLER_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20065__102 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__inv_2
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ clknet_leaf_4_i_clk _00593_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20755_ clknet_leaf_38_i_clk _00524_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20686_ clknet_leaf_29_i_clk _00470_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10370_ _03515_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21307_ net228 _01076_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12040_ _04163_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__buf_2
X_21238_ clknet_leaf_80_i_clk _01007_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19609__63 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_132_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21169_ clknet_leaf_64_i_clk _00938_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19624__77 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__inv_2
X_13991_ _06698_ _06726_ _06671_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__o31a_1
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _08302_ _08374_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__xor2_2
X_12942_ _05604_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__clkinv_2
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _08299_ _08305_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__xor2_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _04000_ _05488_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nand2_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17400_ _09965_ _09966_ vssd1 vssd1 vccd1 vccd1 _09967_ sky130_fd_sc_hd__xnor2_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07218_ _07323_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__xor2_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _02075_ _02077_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__nand2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _04597_ _04600_ _04332_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__mux2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _08231_ _08236_ _05209_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__a21o_4
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09899_ sky130_fd_sc_hd__and2_1
XFILLER_186_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14543_ _07160_ _07199_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__xor2_1
XFILLER_42_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11755_ _04531_ _04532_ _04138_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_1
XFILLER_42_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17262_ _09837_ vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__clkbuf_1
X_10706_ _03694_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14474_ _07203_ _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _04430_ _04431_ _04450_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and3_2
X_19001_ _02631_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__clkbuf_1
X_16213_ _08855_ _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__nand2_1
X_13425_ _05978_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__nor2_1
X_10637_ _03646_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__clkbuf_4
X_17193_ _09774_ _09776_ vssd1 vssd1 vccd1 vccd1 _09778_ sky130_fd_sc_hd__nand2_1
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16144_ _08769_ _08788_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__xnor2_1
X_13356_ _05945_ _05949_ _05939_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a21oi_1
X_10568_ _03621_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12307_ _05062_ _05075_ _05035_ net25 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__o211a_1
XFILLER_170_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16075_ _07989_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__or3_1
XFILLER_114_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10499_ _03585_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
X_13287_ _06010_ _06012_ _06023_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__a21o_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _07684_ _07689_ _07690_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__o21ai_2
X_19903_ rbzero.pov.ready_buffer\[48\] _02823_ _03193_ _03205_ vssd1 vssd1 vccd1 vccd1
+ _03206_ sky130_fd_sc_hd__a211o_1
X_12238_ _04996_ _05005_ _04986_ _05007_ net19 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__o2111a_1
XFILLER_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _04907_ _04905_ _04938_ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a31o_1
X_19834_ _07901_ _03143_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__nand2_1
XFILLER_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19765_ rbzero.pov.spi_buffer\[56\] rbzero.pov.spi_buffer\[57\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
X_16977_ _09498_ _09512_ _09510_ vssd1 vssd1 vccd1 vccd1 _09617_ sky130_fd_sc_hd__a21o_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 i_gpout0_sel[3] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_6
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18716_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__and2_1
X_15928_ _08096_ _08572_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__or2_1
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ rbzero.pov.spi_buffer\[23\] rbzero.pov.spi_buffer\[24\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
XFILLER_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03296_ _03296_ vssd1 vssd1 vccd1 vccd1 clknet_0__03296_ sky130_fd_sc_hd__clkbuf_16
X_18647_ _10248_ _02150_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__and2_1
X_15859_ _08496_ _08502_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__nor2_1
XFILLER_80_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18578_ _02273_ _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__xor2_1
XFILLER_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17529_ _08178_ _08493_ _08044_ _10094_ vssd1 vssd1 vccd1 vccd1 _10095_ sky130_fd_sc_hd__o22ai_1
XFILLER_162_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20540_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03431_
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20471_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03373_
+ sky130_fd_sc_hd__and2_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21023_ clknet_leaf_65_i_clk _00792_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20807_ clknet_leaf_14_i_clk _00576_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11540_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] _04319_ vssd1 vssd1 vccd1
+ vccd1 _04320_ sky130_fd_sc_hd__o31a_2
XFILLER_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20738_ clknet_leaf_1_i_clk _00507_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _04250_ vssd1 vssd1 vccd1 vccd1 _04251_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20669_ clknet_leaf_11_i_clk _00453_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ rbzero.tex_r1\[9\] rbzero.tex_r1\[10\] _03538_ vssd1 vssd1 vccd1 vccd1 _03543_
+ sky130_fd_sc_hd__mux2_1
X_13210_ _05865_ _05870_ _05875_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nor3b_2
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14190_ _06769_ _06677_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__o21ba_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10353_ rbzero.tex_r1\[42\] rbzero.tex_r1\[43\] _03505_ vssd1 vssd1 vccd1 vccd1 _03507_
+ sky130_fd_sc_hd__mux2_1
X_13141_ _05827_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__clkinv_2
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _05740_ _05777_ _05790_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__or3_1
XFILLER_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12023_ rbzero.tex_b1\[35\] rbzero.tex_b1\[34\] _04337_ vssd1 vssd1 vccd1 vccd1 _04798_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16900_ _08170_ _09419_ _09540_ vssd1 vssd1 vccd1 vccd1 _09541_ sky130_fd_sc_hd__or3_1
X_17880_ _09522_ _09029_ _01582_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__or3_1
XFILLER_120_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16831_ _09352_ _09361_ vssd1 vssd1 vccd1 vccd1 _09472_ sky130_fd_sc_hd__or2b_1
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19550_ rbzero.pov.spi_counter\[0\] _03019_ rbzero.pov.spi_counter\[1\] vssd1 vssd1
+ vccd1 vccd1 _03023_ sky130_fd_sc_hd__a21o_1
XFILLER_111_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16762_ _09386_ _09403_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__xor2_1
X_13974_ _06031_ _06707_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__nor2_1
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18501_ _02164_ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15713_ _08355_ _08357_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__and2_1
X_12925_ _05650_ _05655_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__or3_2
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19481_ _02905_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _02961_
+ sky130_fd_sc_hd__nor2_1
X_16693_ _09334_ _09335_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__or2b_1
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18432_ _02128_ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nand2_1
XFILLER_61_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15644_ _08191_ _08265_ _08277_ _08267_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__a22o_1
X_12856_ rbzero.wall_tracer.rayAddendX\[-3\] _05592_ _05560_ vssd1 vssd1 vccd1 vccd1
+ _05593_ sky130_fd_sc_hd__mux2_2
XFILLER_62_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _01951_ _01963_ _02061_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a21o_1
X_11807_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _04341_ vssd1 vssd1 vccd1 vccd1 _04585_
+ sky130_fd_sc_hd__mux2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20202__226 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__inv_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _07560_ _07562_ _07564_ _08171_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__or4_1
X_12787_ _05530_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _09880_ _09881_ _09882_ vssd1 vssd1 vccd1 vccd1 _09884_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14526_ _07070_ _07079_ _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__a21oi_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18294_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__xor2_1
X_11738_ _04510_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__or2_1
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17245_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09822_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14457_ _07184_ _07193_ _07191_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__a21oi_1
X_11669_ _04422_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__nand2_2
XFILLER_128_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ _06091_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and2b_1
XFILLER_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17176_ rbzero.traced_texa\[4\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a22o_1
X_14388_ _07122_ _07124_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__or2b_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ _08768_ _08770_ _08771_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__o21a_1
XFILLER_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13339_ _06044_ _06047_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__and2b_1
XFILLER_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16058_ _07601_ _08148_ _07990_ _07962_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__and4_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15009_ rbzero.wall_tracer.stepDistX\[11\] _07589_ _05201_ vssd1 vssd1 vccd1 vccd1
+ _07675_ sky130_fd_sc_hd__mux2_1
XFILLER_97_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19817_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03317_ clknet_0__03317_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03317_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19748_ rbzero.pov.spi_buffer\[48\] rbzero.pov.spi_buffer\[49\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
X_19603__58 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19679_ rbzero.pov.spi_buffer\[15\] rbzero.pov.spi_buffer\[16\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ clknet_leaf_20_i_clk _01410_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20177__203 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__inv_2
X_21572_ net493 _01341_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_10 _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_21 _09483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_32 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_43 _04140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20523_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03417_
+ sky130_fd_sc_hd__nand2_1
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20454_ _03351_ _03355_ _03352_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o21ai_1
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_84_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21006_ clknet_leaf_51_i_clk _00775_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10971_ _03833_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12710_ _05416_ _05442_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nand2_1
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13690_ _06394_ _06416_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _05391_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15360_ _08004_ rbzero.debug_overlay.playerY\[-7\] _05374_ vssd1 vssd1 vccd1 vccd1
+ _08005_ sky130_fd_sc_hd__mux2_1
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[11\] vssd1
+ vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__nand2_1
XFILLER_211_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14311_ _06067_ _06678_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__or3b_1
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ rbzero.tex_r0\[31\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__and3_1
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15291_ _07933_ _07536_ _07935_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__o21ai_2
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17030_ _09276_ _08111_ vssd1 vssd1 vccd1 vccd1 _09670_ sky130_fd_sc_hd__nor2_2
X_14242_ _06967_ _06968_ _06976_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__a211oi_1
X_11454_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _04214_ vssd1 vssd1 vccd1 vccd1 _04234_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ rbzero.tex_r1\[17\] rbzero.tex_r1\[18\] _03527_ vssd1 vssd1 vccd1 vccd1 _03534_
+ sky130_fd_sc_hd__mux2_1
X_14173_ _06887_ _06901_ _06909_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__o21a_1
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11385_ rbzero.row_render.size\[0\] vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__inv_2
XFILLER_125_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ _05645_ _05796_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__o21ai_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10336_ rbzero.tex_r1\[50\] rbzero.tex_r1\[51\] _03494_ vssd1 vssd1 vccd1 vccd1 _03498_
+ sky130_fd_sc_hd__mux2_1
X_18981_ rbzero.pov.spi_buffer\[23\] rbzero.pov.ready_buffer\[23\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XFILLER_140_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13055_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__buf_2
X_17932_ _10134_ _10131_ _01527_ _01525_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__a31o_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12006_ _04779_ _04780_ _04304_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__mux2_1
XFILLER_39_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17863_ _01563_ _01565_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__nand2_1
XFILLER_87_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16814_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09456_ sky130_fd_sc_hd__or2_2
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xnet99_4 clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
X_17794_ _08188_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__buf_2
XFILLER_19_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19533_ _02906_ _04034_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or3_1
X_16745_ _07996_ _08705_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__or4_1
X_13957_ _06681_ _06688_ _06691_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_47_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12908_ _05618_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__xor2_4
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19464_ _02944_ _02945_ _04029_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__o21ai_1
X_16676_ _09153_ _09155_ vssd1 vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__nor2_1
X_13888_ _06622_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15627_ _07549_ _08270_ _08271_ _07933_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__a211o_2
X_18415_ _02112_ _02113_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__and2_1
XFILLER_59_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12839_ rbzero.wall_tracer.visualWallDist\[10\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05576_ sky130_fd_sc_hd__a21o_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19395_ _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__nand2_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ _08802_ _09668_ _01524_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__or3_2
XFILLER_194_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _05208_ rbzero.wall_tracer.stepDistX\[0\] vssd1 vssd1 vccd1 vccd1 _08203_
+ sky130_fd_sc_hd__nand2_1
X_14509_ _07235_ _07244_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__a21oi_1
X_18277_ _01975_ _01976_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__nor2_1
X_15489_ _04013_ rbzero.wall_tracer.stepDistY\[-12\] vssd1 vssd1 vccd1 vccd1 _08134_
+ sky130_fd_sc_hd__or2_1
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17228_ _05203_ vssd1 vssd1 vccd1 vccd1 _09807_ sky130_fd_sc_hd__clkbuf_4
Xinput30 i_gpout4_sel[4] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_135_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 i_reg_csb vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_6
Xinput52 i_vec_sclk vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17159_ rbzero.traced_texa\[-10\] _09766_ _09767_ _07601_ vssd1 vssd1 vccd1 vccd1
+ _00547_ sky130_fd_sc_hd__a22o_1
XFILLER_192_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21624_ clknet_leaf_22_i_clk _01393_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21555_ net476 _01324_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20506_ _03396_ _03399_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__nand2_1
X_21486_ net407 _01255_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ _03338_ _03341_ _03339_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__a21boi_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11170_ rbzero.otherx\[2\] _03929_ _03935_ rbzero.othery\[4\] vssd1 vssd1 vccd1 vccd1
+ _03959_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_161_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20231__252 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__inv_2
XFILLER_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _07433_ _07445_ _07446_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__nor3_1
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _06497_ _06498_ _06547_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ _07511_ _07437_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__nor2_1
XFILLER_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16530_ _09168_ _09173_ vssd1 vssd1 vccd1 vccd1 _09174_ sky130_fd_sc_hd__xnor2_1
X_13742_ _06475_ _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__xnor2_1
X_19594__49 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
X_10954_ _03824_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16461_ _07941_ _09103_ _09010_ _09104_ vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__o31a_1
X_13673_ _06408_ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__xor2_1
XFILLER_73_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10885_ _03788_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18200_ _01804_ _01900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__xor2_1
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15412_ rbzero.wall_tracer.visualWallDist\[2\] _04015_ vssd1 vssd1 vccd1 vccd1 _08057_
+ sky130_fd_sc_hd__nand2_2
X_19180_ rbzero.spi_registers.new_leak\[1\] _02733_ vssd1 vssd1 vccd1 vccd1 _02735_
+ sky130_fd_sc_hd__or2_1
X_12624_ _03925_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__xnor2_1
X_16392_ _08352_ _08355_ _09036_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18131_ _01582_ _01706_ _01708_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__o21a_1
X_15343_ _05206_ _07984_ _07987_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__o21ai_4
X_12555_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or2_2
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11506_ rbzero.tex_r0\[2\] _04214_ _04219_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__a21o_1
X_18062_ _01755_ _01762_ _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nand3_1
X_15274_ rbzero.wall_tracer.visualWallDist\[-5\] _04012_ rbzero.wall_tracer.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__a21o_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ rbzero.wall_tracer.trackDistX\[-10\] vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__inv_2
XFILLER_176_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17013_ _09638_ _09652_ vssd1 vssd1 vccd1 vccd1 _09653_ sky130_fd_sc_hd__xnor2_1
X_14225_ _06946_ _06949_ _06961_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__a21oi_1
X_20314__327 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__inv_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ _04125_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__buf_6
XFILLER_99_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14156_ _06865_ _06867_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11368_ rbzero.row_render.size\[1\] rbzero.row_render.size\[0\] vssd1 vssd1 vccd1
+ vccd1 _04148_ sky130_fd_sc_hd__nor2_1
XFILLER_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ _05811_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__buf_2
XFILLER_152_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10319_ rbzero.tex_r1\[58\] rbzero.tex_r1\[59\] _03483_ vssd1 vssd1 vccd1 vccd1 _03489_
+ sky130_fd_sc_hd__mux2_1
X_14087_ _06666_ _06668_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__nor2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ rbzero.pov.spi_buffer\[15\] rbzero.pov.ready_buffer\[15\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XFILLER_140_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11299_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _04079_ sky130_fd_sc_hd__nand2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _05684_ _05689_ _05703_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a2bb2o_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17915_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18895_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] _02564_
+ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a21o_1
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17846_ _01548_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__nor2_4
XFILLER_113_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17777_ _01479_ _01480_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14989_ rbzero.wall_tracer.stepDistX\[1\] _07560_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07665_ sky130_fd_sc_hd__mux2_1
XFILLER_187_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19516_ _02905_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 _02994_
+ sky130_fd_sc_hd__or2_1
X_16728_ _09367_ _09369_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__xor2_1
XFILLER_207_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19447_ _02913_ _02916_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a21oi_1
X_16659_ _09132_ _09144_ _09301_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__a21bo_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19378_ rbzero.debug_overlay.vplaneY\[-6\] _02849_ _04034_ vssd1 vssd1 vccd1 vccd1
+ _02866_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18329_ _01971_ _02027_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__xor2_2
XFILLER_72_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21340_ net261 _01109_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21271_ clknet_leaf_65_i_clk _01040_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_118_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20289__304 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__inv_2
XFILLER_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20986_ clknet_leaf_50_i_clk _00755_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ _03675_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21607_ net148 _01376_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ net41 _05084_ _05107_ net43 net29 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a221o_1
X_21538_ net459 _01307_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12271_ _05036_ _05037_ _05038_ _05039_ net22 net21 vssd1 vssd1 vccd1 vccd1 _05040_
+ sky130_fd_sc_hd__mux4_1
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21469_ net390 _01238_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _06680_ _06662_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__nor2_1
XFILLER_181_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ gpout0.hpos\[7\] gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__or2_1
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11153_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15961_ _08582_ _08568_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__xnor2_2
X_11084_ _03892_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17700_ _09117_ _09991_ vssd1 vssd1 vccd1 vccd1 _10265_ sky130_fd_sc_hd__nor2_1
X_14912_ _05278_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__buf_4
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15892_ _08513_ _08534_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__nor2_1
X_18680_ _02208_ _02299_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__and2b_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17631_ _10080_ _10082_ vssd1 vssd1 vccd1 vccd1 _10196_ sky130_fd_sc_hd__nor2_1
X_14843_ rbzero.wall_tracer.stepDistY\[3\] _07564_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07565_ sky130_fd_sc_hd__mux2_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17562_ _05211_ rbzero.wall_tracer.stepDistX\[11\] vssd1 vssd1 vccd1 vccd1 _10128_
+ sky130_fd_sc_hd__nand2_1
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14774_ _07477_ _07470_ _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__a21oi_1
XFILLER_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11986_ rbzero.tex_b1\[10\] _04273_ _04304_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a21o_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16513_ _09030_ _09043_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__nand2_1
X_19301_ _02806_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__clkbuf_1
X_13725_ _06458_ _06460_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__a21o_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10937_ _03815_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17493_ _09245_ _09243_ _09028_ _09164_ vssd1 vssd1 vccd1 vccd1 _10059_ sky130_fd_sc_hd__or4_1
XFILLER_205_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16444_ _08549_ _08957_ _09060_ _09087_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__a31o_1
X_19232_ rbzero.spi_registers.vshift\[2\] _02762_ _02767_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00760_ sky130_fd_sc_hd__o211a_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13656_ _06350_ _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ _03779_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ rbzero.spi_registers.new_other\[2\] _02712_ vssd1 vssd1 vccd1 vccd1 _02723_
+ sky130_fd_sc_hd__or2_1
X_12607_ _05351_ _05353_ _05356_ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__or4_1
XFILLER_157_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _09002_ _09019_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__xnor2_1
X_13587_ _06304_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nand2_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _03743_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
X_18114_ _01805_ _01806_ _01813_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__and3_1
XFILLER_185_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15326_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__clkinv_2
X_19094_ _02680_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__clkbuf_1
X_12538_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__and2_1
XFILLER_200_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ _09674_ _09973_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__nor2_1
X_15257_ _07900_ _07901_ _05495_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__mux2_1
XFILLER_173_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12469_ rbzero.wall_tracer.trackDistX\[4\] vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__inv_2
X_14208_ _06934_ _06939_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o21ai_1
XFILLER_160_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15188_ _07818_ _07819_ _07828_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__nor3_1
XFILLER_158_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14139_ _06859_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ rbzero.pov.ready_buffer\[0\] _03252_ _03253_ rbzero.debug_overlay.vplaneY\[-9\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__o221a_1
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18947_ rbzero.pov.spi_buffer\[7\] rbzero.pov.ready_buffer\[7\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18878_ _02546_ _02547_ _02545_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__o21ai_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17829_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__nand2_1
XFILLER_67_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20840_ clknet_leaf_8_i_clk _00609_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20771_ clknet_leaf_35_i_clk _00540_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21323_ net244 _01092_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21254_ clknet_leaf_61_i_clk _01023_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20205_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__buf_1
X_21185_ clknet_leaf_13_i_clk _00954_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20343__353 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__inv_2
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _04379_ _04614_ _04615_ _04616_ _04209_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o221a_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _04547_ _04548_ _04126_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__mux2_1
XFILLER_198_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ clknet_leaf_69_i_clk _00738_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_202_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13510_ _06244_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__nand2_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _03702_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14490_ _07220_ _07226_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__xor2_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13441_ _06083_ _06086_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__and2b_1
XFILLER_201_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10653_ _03666_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _08803_ _08804_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__or2_1
X_13372_ _06037_ _06092_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__and3_1
XFILLER_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10584_ rbzero.tex_g1\[62\] rbzero.tex_g1\[63\] _03549_ vssd1 vssd1 vccd1 vccd1 _03630_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15111_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__nand2_1
X_12323_ net29 net30 vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__nand2_1
XFILLER_154_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16091_ _08661_ _08735_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__or2_1
XFILLER_108_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15042_ _07695_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__buf_4
X_12254_ _05021_ net61 _05022_ net24 vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__o211a_1
XFILLER_182_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11205_ rbzero.map_rom.f4 rbzero.map_rom.d6 _03921_ _03977_ vssd1 vssd1 vccd1 vccd1
+ _03994_ sky130_fd_sc_hd__or4_1
X_19850_ _03146_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__clkbuf_4
X_12185_ _04930_ _04934_ _04942_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__o31a_1
XFILLER_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18801_ _02480_ _02481_ _02479_ _02476_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__o211a_1
X_11136_ rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__clkinv_2
X_19781_ _03119_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16993_ _09631_ _09632_ vssd1 vssd1 vccd1 vccd1 _09633_ sky130_fd_sc_hd__or2_1
XFILLER_114_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18732_ _02414_ _02416_ _02415_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a21boi_1
X_11067_ _03883_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__clkbuf_1
X_15944_ _08555_ _08554_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__xor2_1
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18663_ _02354_ _02358_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15875_ _07974_ _08519_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__nor2_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _07486_ _07455_ _07551_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__a21oi_4
X_17614_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _10179_ sky130_fd_sc_hd__and2_1
X_18594_ _02288_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _07477_ _07490_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__nor2_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17545_ _10110_ _09417_ _09982_ vssd1 vssd1 vccd1 vccd1 _10111_ sky130_fd_sc_hd__or3_1
X_11969_ _04742_ _04743_ _04345_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__mux2_1
X_13708_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17476_ _09933_ _09936_ _10041_ vssd1 vssd1 vccd1 vccd1 _10042_ sky130_fd_sc_hd__a21oi_2
X_14688_ _07378_ _07413_ _06239_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ _02756_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__clkbuf_1
X_13639_ _06332_ _06331_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__xor2_1
X_16427_ _09069_ _09070_ _09071_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__a21o_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19146_ rbzero.spi_registers.new_other\[6\] _02712_ vssd1 vssd1 vccd1 vccd1 _02713_
+ sky130_fd_sc_hd__or2_1
X_16358_ _07967_ _08674_ _08034_ _08045_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__or4_1
XFILLER_192_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__04835_ _04835_ vssd1 vssd1 vccd1 vccd1 clknet_0__04835_ sky130_fd_sc_hd__clkbuf_16
X_15309_ _07952_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__and2_1
XFILLER_195_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19077_ rbzero.pov.spi_buffer\[69\] rbzero.pov.ready_buffer\[69\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02671_ sky130_fd_sc_hd__mux2_1
X_16289_ _08908_ _08930_ _08931_ _08933_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__and4_1
XFILLER_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18028_ _01728_ _01729_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__xor2_1
XFILLER_195_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19979_ rbzero.pov.ready_buffer\[28\] _03252_ _03253_ rbzero.debug_overlay.facingY\[-3\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__o221a_1
XFILLER_140_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20823_ clknet_leaf_3_i_clk _00592_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20754_ clknet_leaf_38_i_clk _00523_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_126_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20685_ clknet_leaf_27_i_clk _00469_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_210_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21306_ net227 _01075_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21237_ clknet_leaf_80_i_clk _01006_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21168_ clknet_leaf_64_i_clk _00937_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13990_ _06134_ _06677_ _06697_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__o21bai_1
X_21099_ net189 _00868_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _05605_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__clkinv_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _08188_ _08239_ _08302_ _08304_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__o31a_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _05561_ _05459_ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__o21a_2
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _07106_ _07337_ _07347_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nand3_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _04598_ _04599_ _04218_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__mux2_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15591_ _07970_ _08233_ _08234_ _08235_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__o31ai_2
XFILLER_199_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09898_ sky130_fd_sc_hd__nor2_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14542_ _07273_ _07278_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__or2b_1
XFILLER_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11754_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _04129_ vssd1 vssd1 vccd1 vccd1 _04532_
+ sky130_fd_sc_hd__mux2_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17261_ rbzero.wall_tracer.trackDistX\[-9\] _09836_ _05414_ vssd1 vssd1 vccd1 vccd1
+ _09837_ sky130_fd_sc_hd__mux2_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ rbzero.tex_g1\[5\] rbzero.tex_g1\[6\] _03691_ vssd1 vssd1 vccd1 vccd1 _03694_
+ sky130_fd_sc_hd__mux2_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14473_ _07204_ _07209_ _07154_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11685_ _04022_ _04440_ _04450_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__and3_2
XFILLER_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19000_ net513 rbzero.pov.ready_buffer\[32\] _02627_ vssd1 vssd1 vccd1 vccd1 _02631_
+ sky130_fd_sc_hd__mux2_1
X_16212_ _08227_ _08331_ _08856_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__a21o_1
X_13424_ _06119_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__clkbuf_4
X_10636_ _03657_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__clkbuf_1
X_17192_ _09774_ _09776_ vssd1 vssd1 vccd1 vccd1 _09777_ sky130_fd_sc_hd__or2_1
XFILLER_167_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16143_ _08266_ _08039_ _08040_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__and3_1
X_13355_ _06036_ _06035_ _06030_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a21bo_1
X_10567_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _03613_ vssd1 vssd1 vccd1 vccd1 _03621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12306_ _04154_ _03477_ net20 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__mux2_1
XFILLER_155_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16074_ _08692_ _08718_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__xnor2_2
X_13286_ _05973_ _06011_ _06009_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__o21a_1
XFILLER_154_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10498_ rbzero.tex_r0\[40\] rbzero.tex_r0\[39\] _03580_ vssd1 vssd1 vccd1 vccd1 _03585_
+ sky130_fd_sc_hd__mux2_1
XFILLER_114_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15025_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nand2_1
XFILLER_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19902_ _07917_ _03141_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__nor2_1
X_12237_ net16 _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or2_1
XFILLER_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19833_ rbzero.pov.ready_buffer\[62\] _07900_ _03146_ vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__mux2_1
X_12168_ _04021_ _04922_ _04905_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__and3_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _03910_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19764_ _03110_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
X_12099_ _04862_ _04866_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__o21a_1
XFILLER_84_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16976_ _09614_ _09615_ vssd1 vssd1 vccd1 vccd1 _09616_ sky130_fd_sc_hd__nor2_1
XFILLER_110_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__nor2_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _07945_ rbzero.wall_tracer.stepDistX\[-12\] _08135_ vssd1 vssd1 vccd1 vccd1
+ _08572_ sky130_fd_sc_hd__a21boi_2
Xinput6 i_gpout0_sel[4] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_4
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19695_ _03074_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03295_ _03295_ vssd1 vssd1 vccd1 vccd1 clknet_0__03295_ sky130_fd_sc_hd__clkbuf_16
X_18646_ _02340_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__xnor2_1
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _08496_ _08502_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__xor2_1
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ _05884_ _07507_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__nor2_1
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18577_ _09141_ _01475_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__nor2_1
XFILLER_149_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ _08432_ _08433_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17528_ _08202_ vssd1 vssd1 vccd1 vccd1 _10094_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17459_ _10023_ _10025_ vssd1 vssd1 vccd1 vccd1 _10026_ sky130_fd_sc_hd__xor2_4
XFILLER_178_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20095__129 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__inv_2
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20470_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03372_
+ sky130_fd_sc_hd__nor2_1
X_19129_ _02699_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21022_ clknet_leaf_65_i_clk _00791_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_2_0_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ clknet_leaf_14_i_clk _00575_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20737_ clknet_leaf_89_i_clk _00506_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _04211_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__buf_6
X_20668_ clknet_leaf_11_i_clk _00452_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_52_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ _03542_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20599_ _03462_ _03463_ rbzero.wall_tracer.rayAddendY\[-6\] _09762_ vssd1 vssd1 vccd1
+ vccd1 _01431_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_104_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__buf_2
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10352_ _03506_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13071_ _05804_ _05805_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__mux2_1
XFILLER_124_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _04379_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__or2_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16830_ _09381_ _09348_ vssd1 vssd1 vccd1 vccd1 _09471_ sky130_fd_sc_hd__or2b_1
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13973_ _06705_ _06709_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__nand2_1
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16761_ _09393_ _09402_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18500_ _02166_ _02197_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12924_ _05567_ _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__nor2_1
X_15712_ _08329_ _08356_ _08354_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16692_ _09331_ _09333_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__nand2_1
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19480_ rbzero.wall_tracer.rayAddendY\[5\] _07855_ _02955_ _02960_ vssd1 vssd1 vccd1
+ vccd1 _00815_ sky130_fd_sc_hd__a211o_1
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18431_ _02127_ _02129_ _09807_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a21oi_1
X_15643_ _08285_ _08286_ _08287_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__a21bo_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ rbzero.wall_tracer.visualWallDist\[-11\] rbzero.wall_tracer.rayAddendY\[-3\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__mux2_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11806_ _04217_ _04583_ _04123_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__o21a_1
X_18362_ _01960_ _01962_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__nor2_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15574_ _08218_ _08208_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__nand2_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ rbzero.wall_tracer.mapX\[5\] _05529_ _05414_ vssd1 vssd1 vccd1 vccd1 _05530_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _07077_ _07078_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__and2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _09880_ _09881_ _09882_ vssd1 vssd1 vccd1 vccd1 _09883_ sky130_fd_sc_hd__and3_1
XFILLER_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ rbzero.debug_overlay.playerX\[-3\] _04463_ _04511_ _04513_ _04515_ vssd1
+ vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a2111o_1
X_18293_ _01745_ _01988_ _01868_ _01869_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22oi_2
XFILLER_159_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ _07191_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__nor2_1
X_17244_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09821_ sky130_fd_sc_hd__or2_1
X_11668_ _03476_ _04441_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a21bo_4
XFILLER_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ _06131_ _06142_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__a21o_1
XFILLER_174_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17175_ rbzero.traced_texa\[3\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__a22o_1
X_10619_ rbzero.tex_g1\[46\] rbzero.tex_g1\[47\] _03647_ vssd1 vssd1 vccd1 vccd1 _03649_
+ sky130_fd_sc_hd__mux2_1
X_14387_ _07121_ _07123_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__xnor2_1
X_11599_ rbzero.tex_r1\[57\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__and3_1
XFILLER_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _07981_ _08042_ _08720_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__or3_1
X_13338_ _06069_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nand2_1
X_16057_ rbzero.wall_tracer.visualWallDist\[-11\] _04014_ _07990_ _07936_ vssd1 vssd1
+ vccd1 vccd1 _08702_ sky130_fd_sc_hd__and4_1
X_13269_ _06004_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nand2_1
XFILLER_131_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _07674_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ net38 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__o21ai_2
XFILLER_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03316_ clknet_0__03316_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03316_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19747_ _03101_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
X_16959_ _09597_ _09598_ vssd1 vssd1 vccd1 vccd1 _09600_ sky130_fd_sc_hd__and2_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19678_ _03065_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18629_ _02296_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_21640_ clknet_leaf_19_i_clk _01409_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21571_ net492 _01340_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_11 _07041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_22 _09611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_33 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20522_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03416_
+ sky130_fd_sc_hd__nor2_1
XFILLER_123_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_44 _05211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20453_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _03358_
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21005_ clknet_leaf_51_i_clk _00774_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10970_ rbzero.tex_b1\[7\] rbzero.tex_b1\[8\] _03828_ vssd1 vssd1 vccd1 vccd1 _03833_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ _05382_ _05384_ _05381_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__o21bai_1
XFILLER_203_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12571_ rbzero.wall_tracer.rayAddendY\[10\] rbzero.wall_tracer.rayAddendY\[9\] rbzero.debug_overlay.facingY\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__o21ai_1
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _07045_ _07046_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__xor2_1
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11522_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _04213_ vssd1 vssd1 vccd1 vccd1 _04302_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _07933_ _07934_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__nand2_1
XFILLER_211_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _06974_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
XFILLER_156_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11453_ _04210_ _04220_ _04231_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__a211o_1
XFILLER_109_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _03533_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
X_14172_ _06907_ _06908_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__nand2_1
XFILLER_137_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11384_ rbzero.row_render.size\[1\] vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__inv_2
XFILLER_178_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ _05648_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__or4_1
X_10335_ _03497_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18980_ _02620_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13054_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__clkbuf_4
X_17931_ _10110_ _09693_ _01519_ _01633_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__o31ai_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12005_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _04337_ vssd1 vssd1 vccd1 vccd1 _04780_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17862_ _01564_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__inv_2
XFILLER_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16813_ _09451_ _09453_ vssd1 vssd1 vccd1 vccd1 _09455_ sky130_fd_sc_hd__and2_1
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17793_ _08188_ _09276_ _08493_ _08044_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__or4_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19532_ rbzero.debug_overlay.vplaneY\[-1\] _02987_ vssd1 vssd1 vccd1 vccd1 _03008_
+ sky130_fd_sc_hd__nor2_1
X_16744_ _09268_ _09384_ _09385_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__a21o_1
X_13956_ _06679_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nor2_1
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12907_ _05562_ _05566_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__and3_1
XFILLER_62_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19463_ _02942_ _02943_ _07676_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__o21ai_1
X_13887_ _06201_ _06052_ _06623_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__and3_1
X_16675_ _09239_ _09317_ vssd1 vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20126__158 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__inv_2
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18414_ _02106_ _02107_ _02111_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__nand3_1
X_15626_ _07487_ _07455_ _07548_ _07551_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__a22o_1
X_12838_ _05569_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__and2_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ rbzero.debug_overlay.vplaneY\[0\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__nand2_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18345_ _02042_ _02043_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__and2_1
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _08199_ _08201_ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__nand2_4
X_12769_ _05506_ _05507_ _05504_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a21o_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14508_ _07236_ _07243_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__nor2_1
X_15488_ _07460_ _08132_ _07933_ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__mux2_1
X_18276_ _01973_ _01974_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__and2_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 i_gpout3_sel[0] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_8
XFILLER_147_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17227_ _09804_ _09805_ vssd1 vssd1 vccd1 vccd1 _09806_ sky130_fd_sc_hd__nor2_1
Xinput31 i_gpout4_sel[5] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_4
X_14439_ _06689_ _06740_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__nor2_1
XFILLER_190_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput42 i_reg_mosi vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_6
XFILLER_190_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17158_ rbzero.traced_texa\[-11\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22o_1
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _08742_ _08752_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__nor2_1
XFILLER_66_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17089_ _09726_ _09728_ vssd1 vssd1 vccd1 vccd1 _09729_ sky130_fd_sc_hd__xor2_2
XFILLER_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21623_ clknet_leaf_22_i_clk _01392_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21554_ net475 _01323_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20505_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03402_
+ sky130_fd_sc_hd__nand2_1
XFILLER_166_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21485_ net406 _01254_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20436_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03344_
+ sky130_fd_sc_hd__and2_1
XFILLER_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19579__36 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XFILLER_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _06499_ _06465_ _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__or3_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _07459_ _07519_ _07521_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__and3_1
XFILLER_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13741_ _05946_ _05899_ _06007_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__or3_1
X_10953_ rbzero.tex_b1\[15\] rbzero.tex_b1\[16\] _03817_ vssd1 vssd1 vccd1 vccd1 _03824_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13672_ _06041_ _06406_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__or2_1
X_16460_ _08360_ _09009_ vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__nand2_1
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10884_ rbzero.tex_b1\[48\] rbzero.tex_b1\[49\] _03784_ vssd1 vssd1 vccd1 vccd1 _03788_
+ sky130_fd_sc_hd__mux2_1
X_15411_ _08043_ _08055_ vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__xnor2_1
X_12623_ _05375_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__nor2_1
X_16391_ _09034_ _09035_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__xor2_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18130_ _01829_ _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__xnor2_1
X_15342_ rbzero.debug_overlay.playerX\[-8\] _05496_ _07986_ _05196_ vssd1 vssd1 vccd1
+ vccd1 _07987_ sky130_fd_sc_hd__a211o_1
XFILLER_197_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12554_ _05289_ _05295_ _05300_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__and4_1
XFILLER_200_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ rbzero.tex_r0\[3\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__and3_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18061_ _01760_ _01761_ _01756_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a21o_1
X_15273_ _07917_ rbzero.debug_overlay.playerY\[-5\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _07918_ sky130_fd_sc_hd__mux2_1
XFILLER_185_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12485_ rbzero.wall_tracer.trackDistX\[-9\] vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__03319_ clknet_0__03319_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03319_
+ sky130_fd_sc_hd__clkbuf_16
X_14224_ _06953_ _06960_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17012_ _09650_ _09651_ vssd1 vssd1 vccd1 vccd1 _09652_ sky130_fd_sc_hd__nor2_1
X_11436_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _04214_ vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_165_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14155_ _06890_ _06891_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__xnor2_1
X_11367_ rbzero.row_render.size\[2\] vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__inv_2
XFILLER_99_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13106_ _05841_ _05842_ _05807_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__mux2_1
X_10318_ _03488_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14086_ _06802_ _06811_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__xnor2_1
X_18963_ _02611_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
X_11298_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _04078_ sky130_fd_sc_hd__or2_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13037_ _05716_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__nor2_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _08257_ _08044_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__nor2_1
XFILLER_152_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18894_ _02560_ _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__nor2_1
XFILLER_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17845_ _01441_ _01547_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__and2_1
XFILLER_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17776_ _07974_ _08427_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__nor2_1
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14988_ _00008_ _07555_ _07664_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__a21oi_1
X_19515_ _02906_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 _02993_
+ sky130_fd_sc_hd__and2_1
XFILLER_93_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16727_ _09368_ _08427_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__nor2_1
X_13939_ _06605_ _06611_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__and2_1
XFILLER_74_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19446_ _02927_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__nand2_1
X_16658_ _09143_ _09140_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__or2b_1
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_i_clk clknet_opt_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15609_ _05193_ _08172_ _08174_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__a21o_1
X_19377_ rbzero.debug_overlay.vplaneY\[-6\] _02849_ vssd1 vssd1 vccd1 vccd1 _02865_
+ sky130_fd_sc_hd__or2_1
X_16589_ _09003_ _09006_ _09173_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18328_ _10110_ _02026_ _01967_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__o21a_1
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18259_ _01953_ _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21270_ clknet_leaf_65_i_clk _01039_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20083_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__buf_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20109__142 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__inv_2
X_20985_ clknet_leaf_51_i_clk _00754_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20261__279 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__inv_2
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21606_ net147 _01375_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21537_ net458 _01306_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _04891_ _04992_ _04890_ _04892_ _05024_ _05021_ vssd1 vssd1 vccd1 vccd1 _05039_
+ sky130_fd_sc_hd__mux4_1
XFILLER_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21468_ net389 _01237_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11221_ gpout0.hpos\[5\] gpout0.hpos\[4\] gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1
+ _04008_ sky130_fd_sc_hd__and3_1
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20419_ _03325_ _03328_ _03329_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nand3b_1
XFILLER_150_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20155__184 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__inv_2
XFILLER_162_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21399_ net320 _01168_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11152_ rbzero.debug_overlay.playerX\[5\] rbzero.wall_tracer.mapX\[5\] vssd1 vssd1
+ vccd1 vccd1 _03941_ sky130_fd_sc_hd__nand2_1
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15960_ _08587_ _08604_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__xor2_2
X_11083_ rbzero.tex_b0\[18\] rbzero.tex_b0\[17\] _03887_ vssd1 vssd1 vccd1 vccd1 _03892_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14911_ _07591_ _07614_ _07615_ _04039_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__o211a_1
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _08505_ _08489_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__xnor2_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ _10042_ _10194_ vssd1 vssd1 vccd1 vccd1 _10195_ sky130_fd_sc_hd__xor2_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _07459_ _07453_ _07468_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__o21bai_4
XFILLER_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ _10125_ _10126_ vssd1 vssd1 vccd1 vccd1 _10127_ sky130_fd_sc_hd__or2_1
X_14773_ _07477_ _07476_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__nor2_1
X_11985_ rbzero.tex_b1\[11\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__and3_1
XFILLER_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19300_ rbzero.spi_registers.new_other\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
X_16512_ _09153_ _09155_ vssd1 vssd1 vccd1 vccd1 _09156_ sky130_fd_sc_hd__xor2_1
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13724_ _06391_ _06419_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__xnor2_1
X_10936_ rbzero.tex_b1\[23\] rbzero.tex_b1\[24\] _03806_ vssd1 vssd1 vccd1 vccd1 _03815_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17492_ _09245_ _09029_ _09165_ _09243_ vssd1 vssd1 vccd1 vccd1 _10058_ sky130_fd_sc_hd__o22ai_1
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20320__332 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__inv_2
XFILLER_147_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19231_ rbzero.spi_registers.new_vshift\[2\] _02763_ vssd1 vssd1 vccd1 vccd1 _02767_
+ sky130_fd_sc_hd__or2_1
XFILLER_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16443_ _09059_ _08547_ vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__and2b_1
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13655_ _06351_ _06369_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__xor2_1
XFILLER_90_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ rbzero.tex_b1\[56\] rbzero.tex_b1\[57\] _03773_ vssd1 vssd1 vccd1 vccd1 _03779_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12606_ _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__xnor2_2
X_19162_ rbzero.othery\[1\] _02710_ _02720_ _02722_ vssd1 vssd1 vccd1 vccd1 _00735_
+ sky130_fd_sc_hd__o211a_1
X_13586_ _06305_ _06321_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a21oi_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16374_ _09008_ _09018_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__xor2_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ rbzero.tex_g0\[26\] rbzero.tex_g0\[25\] _03740_ vssd1 vssd1 vccd1 vccd1 _03743_
+ sky130_fd_sc_hd__mux2_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18113_ _01805_ _01806_ _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12537_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__xor2_2
X_15325_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__buf_4
XFILLER_185_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19093_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.spi_buffer\[1\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _01744_ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ _05220_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.trackDistY\[5\]
+ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a2bb2o_1
X_15256_ rbzero.debug_overlay.playerX\[-6\] vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__inv_2
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14207_ _06942_ _06943_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__nand2_1
X_11419_ gpout0.hpos\[6\] _04184_ _04182_ gpout0.hpos\[7\] _04198_ vssd1 vssd1 vccd1
+ vccd1 _04199_ sky130_fd_sc_hd__o221a_1
XFILLER_126_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15187_ _07829_ _07832_ _07840_ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__o21bai_1
X_12399_ _04006_ _03475_ _04992_ _04892_ _05143_ net34 vssd1 vssd1 vccd1 vccd1 _05166_
+ sky130_fd_sc_hd__mux4_1
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14138_ _06860_ _06874_ _06872_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a21o_1
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19995_ rbzero.pov.ready_buffer\[21\] _03252_ _03253_ _07821_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01036_ sky130_fd_sc_hd__o221a_1
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ _06805_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__and3b_1
X_18946_ _02602_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18877_ _02549_ _02316_ rbzero.wall_tracer.trackDistY\[10\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00623_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17828_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__nor2_1
XFILLER_39_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17759_ _01462_ _09029_ _09165_ _09526_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__o22a_1
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20770_ clknet_leaf_33_i_clk _00539_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19429_ _04471_ rbzero.debug_overlay.vplaneY\[-7\] _02910_ _02911_ vssd1 vssd1 vccd1
+ vccd1 _02913_ sky130_fd_sc_hd__or4_1
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21322_ net243 _01091_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21253_ clknet_leaf_81_i_clk _01022_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_190_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21184_ clknet_leaf_76_i_clk _00953_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _04341_ vssd1 vssd1 vccd1 vccd1 _04548_
+ sky130_fd_sc_hd__mux2_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ clknet_leaf_68_i_clk _00737_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ rbzero.tex_g0\[62\] rbzero.tex_g0\[61\] _03624_ vssd1 vssd1 vccd1 vccd1 _03702_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20899_ clknet_leaf_84_i_clk _00668_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _06115_ _06176_ _06085_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__and3_1
XFILLER_186_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ rbzero.tex_g1\[30\] rbzero.tex_g1\[31\] _03658_ vssd1 vssd1 vccd1 vccd1 _03666_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _06097_ _06098_ _06106_ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__a31o_1
XFILLER_210_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _03629_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ net31 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__inv_2
XFILLER_177_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15110_ _07756_ _07761_ _07762_ _07768_ vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a31o_1
XFILLER_103_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16090_ _08570_ _08579_ _08571_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__o21a_1
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15041_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__or2_1
X_12253_ _05021_ _04666_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__nand2_1
XFILLER_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ _03988_ _03989_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__or3b_1
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ net13 _04953_ _04954_ _04922_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a22o_1
XFILLER_150_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18800_ _02482_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__inv_2
XFILLER_150_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11135_ rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__clkinv_2
XFILLER_123_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19780_ rbzero.pov.spi_buffer\[63\] rbzero.pov.spi_buffer\[64\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16992_ _08335_ _09217_ _09489_ _09490_ vssd1 vssd1 vccd1 vccd1 _09632_ sky130_fd_sc_hd__o31a_1
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18731_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__and2_1
X_11066_ rbzero.tex_b0\[26\] rbzero.tex_b0\[25\] _03876_ vssd1 vssd1 vccd1 vccd1 _03883_
+ sky130_fd_sc_hd__mux2_1
X_15943_ _08526_ _08528_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__xnor2_2
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18662_ _02255_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15874_ _08518_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__clkbuf_4
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17613_ rbzero.wall_tracer.trackDistX\[1\] _09817_ _10173_ _10178_ vssd1 vssd1 vccd1
+ vccd1 _00590_ sky130_fd_sc_hd__o22a_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _07473_ _07527_ _07499_ _07376_ _05834_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__a32o_2
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _02163_ _02199_ _02289_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a21oi_1
XFILLER_184_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _09114_ vssd1 vssd1 vccd1 vccd1 _10110_ sky130_fd_sc_hd__clkbuf_4
X_14756_ _07351_ _07361_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__nor2_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11968_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _04290_ vssd1 vssd1 vccd1 vccd1 _04743_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ _05846_ _06009_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__or2_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _03646_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17475_ _08416_ _09704_ _09924_ _09922_ vssd1 vssd1 vccd1 vccd1 _10041_ sky130_fd_sc_hd__o31a_1
X_14687_ _07106_ _07419_ _07420_ _07423_ _05742_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__a311oi_2
X_11899_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _04290_ vssd1 vssd1 vccd1 vccd1 _04675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_149_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19214_ _09753_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__and2_1
X_16426_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerX\[-8\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__mux2_1
X_13638_ _06347_ _06373_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__a21boi_2
X_19145_ rbzero.spi_registers.got_new_other _02711_ vssd1 vssd1 vccd1 vccd1 _02712_
+ sky130_fd_sc_hd__nand2_2
XFILLER_146_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16357_ _08289_ _08294_ _09001_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__a21bo_1
X_13569_ _06097_ _06098_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__and2_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15308_ rbzero.debug_overlay.playerY\[-5\] _07906_ rbzero.debug_overlay.playerY\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19076_ _02670_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16288_ _08901_ _08932_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__nor2_1
XFILLER_195_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18027_ _01592_ _01601_ _01599_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a21oi_1
XFILLER_161_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15239_ rbzero.wall_tracer.rayAddendX\[11\] _07887_ vssd1 vssd1 vccd1 vccd1 _07888_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19978_ _03242_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__buf_2
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18929_ rbzero.spi_registers.spi_counter\[6\] _02589_ _02592_ vssd1 vssd1 vccd1 vccd1
+ _00632_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20822_ clknet_leaf_4_i_clk _00591_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20753_ clknet_leaf_38_i_clk _00522_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20684_ clknet_leaf_27_i_clk _00468_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21305_ net226 _01074_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21236_ clknet_leaf_80_i_clk _01005_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21167_ clknet_leaf_64_i_clk _00936_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21098_ net188 _00867_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20049_ _04891_ _03281_ _04890_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a21oi_1
X_20267__285 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__inv_2
X_12940_ _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__xor2_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _04030_ _05367_ _05368_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a31o_1
XFILLER_206_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14610_ _07343_ _07344_ _07346_ _07107_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__o211ai_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11822_ rbzero.tex_g1\[53\] rbzero.tex_g1\[52\] _04212_ vssd1 vssd1 vccd1 vccd1 _04599_
+ sky130_fd_sc_hd__mux2_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _07970_ _08222_ _08223_ _08002_ vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__a31oi_4
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14541_ _07276_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nor2_1
X_11753_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _04129_ vssd1 vssd1 vccd1 vccd1 _04531_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _03693_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__clkbuf_1
X_17260_ _09812_ _09833_ _09834_ _09835_ vssd1 vssd1 vccd1 vccd1 _09836_ sky130_fd_sc_hd__o31ai_1
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14472_ _07148_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11684_ _04004_ _04438_ _04450_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__and3_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16211_ _08377_ _08054_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__nor2_1
X_13423_ _05983_ _06159_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__nor2_1
X_10635_ rbzero.tex_g1\[38\] rbzero.tex_g1\[39\] _03647_ vssd1 vssd1 vccd1 vccd1 _03657_
+ sky130_fd_sc_hd__mux2_1
X_17191_ rbzero.wall_tracer.mapX\[5\] _05512_ _09775_ vssd1 vssd1 vccd1 vccd1 _09776_
+ sky130_fd_sc_hd__o21a_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13354_ _06051_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16142_ _08782_ _08783_ _08786_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__o21ai_1
X_10566_ _03620_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ net22 _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or2_1
X_13285_ _06014_ _06018_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__xor2_2
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16073_ _08693_ _08717_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__xor2_2
X_10497_ _03584_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12236_ _04813_ _04811_ _04006_ _03475_ _04961_ _04960_ vssd1 vssd1 vccd1 vccd1 _05006_
+ sky130_fd_sc_hd__mux4_1
X_15024_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] _07688_
+ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__a21oi_1
X_19901_ rbzero.debug_overlay.playerY\[-6\] _03198_ _03204_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00992_ sky130_fd_sc_hd__o211a_1
XFILLER_155_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19832_ _03139_ _03150_ _03151_ _02765_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__o211a_1
X_12167_ net41 net43 net8 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__mux2_1
XFILLER_111_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11118_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _03557_ vssd1 vssd1 vccd1 vccd1 _03910_
+ sky130_fd_sc_hd__mux2_1
X_19763_ rbzero.pov.spi_buffer\[55\] rbzero.pov.spi_buffer\[56\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
X_12098_ _04868_ _04851_ _04855_ _04869_ net7 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a32o_1
X_16975_ _09514_ _09607_ _09613_ vssd1 vssd1 vccd1 vccd1 _09615_ sky130_fd_sc_hd__and3_1
XFILLER_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18714_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ _02403_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a21oi_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ rbzero.tex_b0\[34\] rbzero.tex_b0\[33\] _03865_ vssd1 vssd1 vccd1 vccd1 _03874_
+ sky130_fd_sc_hd__mux2_1
X_15926_ _08109_ _08491_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__or2_1
X_19694_ rbzero.pov.spi_buffer\[22\] rbzero.pov.spi_buffer\[23\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 i_gpout0_sel[5] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03294_ _03294_ vssd1 vssd1 vccd1 vccd1 clknet_0__03294_ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18645_ _10094_ _09611_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__nand2_1
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _08497_ _08501_ _08499_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__a21boi_1
XFILLER_188_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14808_ _00004_ _07536_ _07537_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18576_ _08151_ _09138_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__nor2_1
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _08161_ _08165_ vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__or2_1
XFILLER_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17527_ _08178_ _08202_ _08493_ _08044_ vssd1 vssd1 vccd1 vccd1 _10093_ sky130_fd_sc_hd__or4_1
X_14739_ _07378_ _07360_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__and2_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17458_ _09474_ _09733_ _10024_ vssd1 vssd1 vccd1 vccd1 _10025_ sky130_fd_sc_hd__a21oi_4
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16409_ _08437_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__inv_2
XFILLER_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17389_ _09673_ _09676_ vssd1 vssd1 vccd1 vccd1 _09956_ sky130_fd_sc_hd__nor2_1
XFILLER_119_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19128_ rbzero.spi_registers.ss_buffer\[1\] rbzero.spi_registers.ss_buffer\[0\] _05189_
+ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_118_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19059_ rbzero.pov.spi_buffer\[60\] rbzero.pov.ready_buffer\[60\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21021_ clknet_leaf_68_i_clk _00790_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ clknet_leaf_14_i_clk _00574_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20736_ clknet_leaf_89_i_clk _00505_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_211_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20667_ clknet_leaf_10_i_clk _00451_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10420_ rbzero.tex_r1\[10\] rbzero.tex_r1\[11\] _03538_ vssd1 vssd1 vccd1 vccd1 _03542_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20598_ _02827_ _02836_ _02835_ _07830_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__a31o_1
X_10351_ rbzero.tex_r1\[43\] rbzero.tex_r1\[44\] _03505_ vssd1 vssd1 vccd1 vccd1 _03506_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__clkbuf_4
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12021_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _04250_ vssd1 vssd1 vccd1 vccd1 _04796_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21219_ clknet_leaf_68_i_clk _00988_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16760_ _09400_ _09401_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__nor2_1
XFILLER_98_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13972_ _05825_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__nor2_1
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15711_ _08059_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__buf_4
X_12923_ _05659_ _05569_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__and2_1
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16691_ _09331_ _09333_ vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__nor2_1
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18430_ _01799_ _02024_ _02025_ _02023_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
X_15642_ _07977_ _07913_ _07924_ _07995_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__or4_1
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ rbzero.wall_tracer.rayAddendX\[-4\] _05590_ _05560_ vssd1 vssd1 vccd1 vccd1
+ _05591_ sky130_fd_sc_hd__mux2_4
XFILLER_185_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18361_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__nor2_1
X_11805_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _04211_ vssd1 vssd1 vccd1 vccd1 _04583_
+ sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _07566_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__inv_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ rbzero.debug_overlay.playerX\[5\] _05528_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05529_ sky130_fd_sc_hd__mux2_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _09872_ _09875_ _09873_ vssd1 vssd1 vccd1 vccd1 _09882_ sky130_fd_sc_hd__o21ai_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14524_ _07237_ _07260_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__xnor2_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18292_ _01990_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__xor2_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ rbzero.debug_overlay.playerX\[2\] _04451_ _04465_ rbzero.debug_overlay.playerX\[-1\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a221o_1
XFILLER_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17243_ _05242_ _09781_ _09820_ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14455_ _07187_ _07190_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__nor2_1
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ gpout0.hpos\[8\] _04442_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__nand2_1
X_13406_ _06130_ _06129_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__and2b_1
X_17174_ _07706_ vssd1 vssd1 vccd1 vccd1 _09770_ sky130_fd_sc_hd__buf_2
X_10618_ _03648_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__clkbuf_1
X_14386_ _06698_ _06760_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nor2_1
X_11598_ _04375_ _04376_ _04219_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
XFILLER_127_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16125_ _08180_ _08042_ _08769_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__o21a_1
X_13337_ _06070_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__xor2_2
X_10549_ _03611_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16056_ _08644_ _08645_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ _05983_ _05982_ _06003_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15007_ rbzero.wall_tracer.stepDistX\[10\] _07586_ _05201_ vssd1 vssd1 vccd1 vccd1
+ _07674_ sky130_fd_sc_hd__mux2_1
X_12219_ gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__buf_2
XFILLER_155_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13199_ _05931_ _05903_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__o21ai_1
XFILLER_123_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19815_ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__buf_2
XFILLER_111_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03315_ clknet_0__03315_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03315_
+ sky130_fd_sc_hd__clkbuf_16
X_16958_ _09597_ _09598_ vssd1 vssd1 vccd1 vccd1 _09599_ sky130_fd_sc_hd__nor2_1
X_19746_ rbzero.pov.spi_buffer\[47\] rbzero.pov.spi_buffer\[48\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03101_ sky130_fd_sc_hd__mux2_1
X_15909_ _08475_ _08553_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__xor2_1
X_19677_ rbzero.pov.spi_buffer\[14\] rbzero.pov.spi_buffer\[15\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16889_ _08178_ _08111_ vssd1 vssd1 vccd1 vccd1 _09530_ sky130_fd_sc_hd__nor2_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18628_ _02288_ _02290_ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__o21a_1
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18559_ _10239_ _09350_ _09481_ _10094_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__o22a_1
XFILLER_178_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21570_ net491 _01339_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[21\] sky130_fd_sc_hd__dfxtp_1
X_20103__137 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__inv_2
XANTENNA_12 _07552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20521_ rbzero.texV\[5\] _03327_ _03332_ _03415_ vssd1 vssd1 vccd1 vccd1 _01401_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_23 _09739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_34 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _09458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20452_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _03357_
+ sky130_fd_sc_hd__or2_1
XFILLER_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21004_ clknet_leaf_49_i_clk _00773_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20184__209 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__inv_2
XFILLER_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20379__386 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__inv_2
XFILLER_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12570_ _05288_ _05319_ _05320_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o211ai_2
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11521_ _04299_ _04300_ _04266_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
X_20078__114 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__inv_2
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20719_ clknet_leaf_15_i_clk _00009_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14240_ _06844_ _06973_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__nor2_1
XFILLER_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ _04119_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__buf_6
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10403_ rbzero.tex_r1\[18\] rbzero.tex_r1\[19\] _03527_ vssd1 vssd1 vccd1 vccd1 _03533_
+ sky130_fd_sc_hd__mux2_1
X_14171_ _06887_ _06901_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__xor2_1
XFILLER_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11383_ gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__clkbuf_4
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10334_ rbzero.tex_r1\[51\] rbzero.tex_r1\[52\] _03494_ vssd1 vssd1 vccd1 vccd1 _03497_
+ sky130_fd_sc_hd__mux2_1
X_13122_ _05857_ _05858_ _05807_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__mux2_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13053_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__or3_1
XFILLER_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17930_ _01514_ _01518_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nand2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12004_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _04337_ vssd1 vssd1 vccd1 vccd1 _04779_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17861_ _09249_ _10200_ _01458_ _01460_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__o22a_1
XFILLER_121_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16812_ _09451_ _09453_ vssd1 vssd1 vccd1 vccd1 _09454_ sky130_fd_sc_hd__nor2_1
XFILLER_113_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17792_ _10257_ _10263_ _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a21oi_2
XFILLER_94_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19531_ rbzero.wall_tracer.rayAddendY\[9\] _07718_ _07831_ _03005_ _03007_ vssd1
+ vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__o221a_1
XFILLER_207_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16743_ _09269_ _09273_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__and2_1
X_13955_ _06680_ _06672_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__nor2_1
XFILLER_98_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12906_ _05610_ _05612_ _05615_ _05601_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a211o_1
X_19462_ _02942_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__and2_1
XFILLER_98_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16674_ _09315_ _09316_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__nor2_1
X_13886_ _05974_ _05983_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__nand2_1
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18413_ _02106_ _02107_ _02111_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a21o_1
X_15625_ _07551_ vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__inv_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _05563_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__nand2_2
X_19393_ rbzero.debug_overlay.vplaneY\[0\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__or2_1
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _09141_ _01620_ _02041_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__o21ai_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _08002_ _08200_ _07945_ vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__a21oi_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12768_ _05511_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or2b_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14507_ _07236_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nand2_1
XFILLER_187_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18275_ _01973_ _01974_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__nor2_1
X_11719_ rbzero.debug_overlay.playerY\[-5\] _04454_ _04458_ rbzero.debug_overlay.playerY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a22o_1
X_15487_ rbzero.wall_tracer.rayAddendY\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] _07893_
+ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__mux2_1
X_12699_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__xnor2_4
X_17226_ _08939_ _08850_ _08936_ vssd1 vssd1 vccd1 vccd1 _09805_ sky130_fd_sc_hd__and3_1
Xinput10 i_gpout1_sel[2] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_4
XFILLER_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14438_ _07172_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput21 i_gpout3_sel[1] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_8
Xinput32 i_gpout5_sel[0] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_2
XFILLER_156_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput43 i_reg_sclk vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_4
XFILLER_122_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17157_ rbzero.traced_texa\[-12\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-12\]
+ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a22o_1
X_14369_ _05931_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__buf_2
XFILLER_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16108_ _08742_ _08752_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__xor2_1
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17088_ _09517_ _09582_ _09727_ vssd1 vssd1 vccd1 vccd1 _09728_ sky130_fd_sc_hd__a21oi_2
XFILLER_170_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16039_ _07958_ _08491_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__or2_1
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19729_ _03047_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21622_ clknet_leaf_22_i_clk _01391_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21553_ net474 _01322_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20504_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03401_
+ sky130_fd_sc_hd__or2_1
XFILLER_166_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21484_ net405 _01253_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20435_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03343_
+ sky130_fd_sc_hd__nor2_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ _05944_ _06016_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__nor2_1
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10952_ _03823_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _06061_ _06407_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__nand2_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _03787_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15410_ _08047_ _08054_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__nor2_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ _03942_ _05374_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__nor2_1
XFILLER_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16390_ _08062_ _08425_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__nor2_1
XFILLER_145_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15341_ _05495_ _07985_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__nor2_1
XFILLER_145_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12553_ _05303_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__and2_1
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ _04282_ _04283_ _04226_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__mux2_1
X_18060_ _01756_ _01760_ _01761_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__nand3_1
X_15272_ rbzero.debug_overlay.playerY\[-5\] _07906_ vssd1 vssd1 vccd1 vccd1 _07917_
+ sky130_fd_sc_hd__xor2_1
Xclkbuf_1_0__f__03318_ clknet_0__03318_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03318_
+ sky130_fd_sc_hd__clkbuf_16
X_12484_ rbzero.wall_tracer.trackDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__inv_2
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17011_ _09647_ _09649_ vssd1 vssd1 vccd1 vccd1 _09651_ sky130_fd_sc_hd__and2_1
X_14223_ _06958_ _06959_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__and2b_1
X_11435_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _04214_ vssd1 vssd1 vccd1 vccd1 _04215_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14154_ _06666_ _06672_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__nor2_1
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11366_ _04137_ _04139_ _04140_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__or4_1
XFILLER_153_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _05690_ _05681_ _05791_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__mux2_1
X_10317_ rbzero.tex_r1\[59\] rbzero.tex_r1\[60\] _03483_ vssd1 vssd1 vccd1 vccd1 _03488_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14085_ _06687_ _06694_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__xor2_1
X_11297_ rbzero.texV\[4\] _04076_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__xor2_1
X_18962_ rbzero.pov.spi_buffer\[14\] rbzero.pov.ready_buffer\[14\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20132__163 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__inv_2
X_13036_ _05598_ _05717_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__xnor2_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _08242_ _09129_ _08129_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a21oi_2
XFILLER_191_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18893_ _02562_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__inv_2
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17844_ _01441_ _01547_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__nor2_1
XFILLER_113_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17775_ _01477_ _01478_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__nand2_1
X_14987_ rbzero.wall_tracer.stepDistX\[0\] _07650_ vssd1 vssd1 vccd1 vccd1 _07664_
+ sky130_fd_sc_hd__nor2_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19514_ _02990_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__nor2_1
X_16726_ _08823_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__buf_2
X_13938_ _06240_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19445_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__nand2_1
XFILLER_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16657_ _09297_ _09298_ _09282_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__a21o_1
X_13869_ _06548_ _06549_ _06551_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__or3_1
Xclkbuf_0__03045_ _03045_ vssd1 vssd1 vccd1 vccd1 clknet_0__03045_ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _08183_ _08185_ _07598_ _08002_ _05208_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__a2111o_1
X_19376_ _02862_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__xnor2_1
X_16588_ _09223_ _09230_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18327_ _10134_ _01878_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__nand2_1
XFILLER_148_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15539_ _07894_ _05335_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__nor2_1
XFILLER_176_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _01956_ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__xor2_1
XFILLER_191_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ rbzero.wall_tracer.mapX\[8\] _05525_ _09790_ vssd1 vssd1 vccd1 vccd1 _09791_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18189_ _01887_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nand3_1
XFILLER_128_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20215__238 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__inv_2
XFILLER_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ clknet_leaf_49_i_clk _00753_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19584__40 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21605_ net146 _01374_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21536_ net457 _01305_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21467_ net388 _01236_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[46\] sky130_fd_sc_hd__dfxtp_1
X_11220_ _04004_ _04005_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20418_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03329_
+ sky130_fd_sc_hd__nand2_1
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21398_ net319 _01167_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11151_ rbzero.debug_overlay.playerX\[5\] rbzero.wall_tracer.mapX\[5\] vssd1 vssd1
+ vccd1 vccd1 _03940_ sky130_fd_sc_hd__or2_1
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20349_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__buf_1
XFILLER_134_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11082_ _03891_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14910_ rbzero.wall_tracer.visualWallDist\[-4\] _07595_ vssd1 vssd1 vccd1 vccd1 _07615_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _08513_ _08534_ vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__xor2_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14841_ _07563_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__clkbuf_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _09700_ _09998_ vssd1 vssd1 vccd1 vccd1 _10126_ sky130_fd_sc_hd__and2_2
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _05814_ _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__or2_1
X_11984_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _04263_ vssd1 vssd1 vccd1 vccd1 _04759_
+ sky130_fd_sc_hd__mux2_1
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16511_ _08998_ _09021_ _09154_ vssd1 vssd1 vccd1 vccd1 _09155_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13723_ _06436_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__or2b_1
X_10935_ _03814_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17491_ _10055_ _10056_ vssd1 vssd1 vccd1 vccd1 _10057_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19230_ rbzero.spi_registers.vshift\[1\] _02762_ _02766_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00759_ sky130_fd_sc_hd__o211a_1
X_20162__189 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__inv_2
X_16442_ _09083_ _09084_ _09086_ _07642_ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__o211a_1
XFILLER_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13654_ _06388_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__and2_1
XFILLER_147_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10866_ _03778_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _05290_ _05293_ _05294_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a21o_1
X_19161_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__clkbuf_4
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _09016_ _09017_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__nor2_1
X_13585_ _06308_ _06320_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__and2b_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _03742_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _01811_ _01812_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__nand2_1
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _07944_ _07968_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__xor2_1
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19092_ _02679_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__clkbuf_1
X_12536_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__or2_1
XFILLER_173_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18043_ _09292_ _09695_ _08802_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a21oi_2
XFILLER_172_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15255_ _07898_ _07899_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ rbzero.wall_tracer.trackDistX\[5\] vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__inv_2
X_14206_ _06934_ _06939_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__xor2_1
X_11418_ _04004_ _04186_ _04184_ gpout0.hpos\[6\] _04197_ vssd1 vssd1 vccd1 vccd1
+ _04198_ sky130_fd_sc_hd__a221o_1
XFILLER_144_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15186_ rbzero.wall_tracer.rayAddendX\[6\] _07695_ _07839_ _03913_ vssd1 vssd1 vccd1
+ vccd1 _07840_ sky130_fd_sc_hd__a22o_1
X_12398_ _05153_ _05149_ _05154_ _05164_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__o31a_1
XFILLER_141_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14137_ _06872_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__and2b_1
XFILLER_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__buf_4
XFILLER_99_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19994_ rbzero.pov.ready_buffer\[20\] _03252_ _03253_ _07742_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01035_ sky130_fd_sc_hd__o221a_1
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14068_ _06009_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__buf_2
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18945_ rbzero.pov.spi_buffer\[6\] rbzero.pov.ready_buffer\[6\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13019_ _05736_ _05735_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__or2_1
XFILLER_140_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18876_ _05532_ _02548_ _02406_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__o21a_1
XFILLER_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _10264_ _10272_ _10271_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17758_ _09522_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__buf_2
XFILLER_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16709_ _05210_ _09350_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__or2_2
X_17689_ _10235_ _10253_ vssd1 vssd1 vccd1 vccd1 _10254_ sky130_fd_sc_hd__xor2_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19428_ _04471_ rbzero.debug_overlay.vplaneY\[-7\] _02910_ _02911_ vssd1 vssd1 vccd1
+ vccd1 _02912_ sky130_fd_sc_hd__o22ai_1
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19359_ rbzero.wall_tracer.rayAddendY\[-4\] _00013_ _02845_ _02848_ vssd1 vssd1 vccd1
+ vccd1 _00806_ sky130_fd_sc_hd__o22a_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21321_ net242 _01090_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20139__169 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__inv_2
XFILLER_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21252_ clknet_leaf_82_i_clk _01021_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_128_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21183_ clknet_leaf_74_i_clk _00952_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19636__88 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__inv_2
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ clknet_leaf_68_i_clk _00736_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _03701_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ clknet_leaf_84_i_clk _00667_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ _03665_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _06102_ _06105_ _06099_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__a21oi_1
X_10582_ rbzero.tex_g1\[63\] net47 _03549_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12321_ _05087_ net61 _05088_ net30 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__o211a_1
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21519_ net440 _01288_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__nand2_1
X_12252_ net20 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20350__359 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__inv_2
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ rbzero.map_rom.f3 rbzero.map_rom.d6 _03990_ _03991_ vssd1 vssd1 vccd1 vccd1
+ _03992_ sky130_fd_sc_hd__o211a_1
X_12183_ net11 net10 _04904_ _04867_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__and4b_1
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11134_ rbzero.debug_overlay.playerX\[0\] _03919_ rbzero.map_rom.i_row\[4\] _03920_
+ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_82_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16991_ _09627_ _09630_ vssd1 vssd1 vccd1 vccd1 _09631_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15942_ _08531_ _08532_ vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__xnor2_2
X_11065_ _03882_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__clkbuf_1
X_18730_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__nor2_1
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18661_ _02355_ _02356_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__nand2_1
XFILLER_188_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _05195_ _08226_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__or2_1
XFILLER_110_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _09889_ _10176_ _10177_ _09780_ vssd1 vssd1 vccd1 vccd1 _10178_ sky130_fd_sc_hd__a31o_1
XFILLER_97_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14824_ _00004_ _07549_ _07550_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a21oi_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__nor2_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20244__264 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__inv_2
XFILLER_205_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17543_ _10090_ _10108_ vssd1 vssd1 vccd1 vccd1 _10109_ sky130_fd_sc_hd__xor2_1
X_14755_ _07107_ _07349_ _07337_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__a21bo_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _04356_ vssd1 vssd1 vccd1 vccd1 _04742_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _05823_ _05909_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__or2_1
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10918_ _03805_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17474_ _09954_ _09919_ vssd1 vssd1 vccd1 vccd1 _10040_ sky130_fd_sc_hd__or2b_1
X_14686_ _05779_ _07337_ _07347_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_20_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _04247_ _04671_ _04672_ _04673_ _04229_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__o221a_1
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19213_ rbzero.spi_registers.new_floor\[2\] rbzero.color_floor\[2\] _02751_ vssd1
+ vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
X_16425_ rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerX\[-9\] _07894_
+ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__mux2_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13637_ _06372_ _06349_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__or2b_1
XFILLER_189_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10849_ _03769_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19144_ _02708_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__clkbuf_4
X_16356_ _08295_ _08288_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__or2b_1
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13568_ _06291_ _06298_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__xor2_2
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ rbzero.debug_overlay.playerY\[-4\] rbzero.debug_overlay.playerY\[-5\] _07906_
+ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__or3_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19075_ rbzero.pov.spi_buffer\[68\] rbzero.pov.ready_buffer\[68\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
X_12519_ _05261_ _05259_ _05256_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_35_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16287_ _08900_ _08885_ _08888_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__and3_1
X_13499_ _05752_ _06153_ _06207_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and3_1
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _01726_ _01727_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nand2_1
X_15238_ _07885_ _07821_ _07886_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__mux2_1
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _07819_ _07822_ _07818_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__a21o_1
XFILLER_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19977_ _03239_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__buf_2
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18928_ rbzero.spi_registers.spi_counter\[6\] _02589_ _02557_ vssd1 vssd1 vccd1 vccd1
+ _02592_ sky130_fd_sc_hd__o21ai_1
XFILLER_171_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18859_ _02530_ _02531_ _02532_ _05203_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__o31a_1
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19641__91 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__inv_2
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20821_ clknet_leaf_5_i_clk _00590_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20752_ clknet_leaf_38_i_clk _00521_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20683_ clknet_leaf_27_i_clk _00467_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21304_ net225 _01073_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21235_ clknet_leaf_78_i_clk _01004_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21166_ clknet_leaf_63_i_clk _00935_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21097_ net187 _00866_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[37\] sky130_fd_sc_hd__dfxtp_1
X_20048_ _04891_ _03281_ _03284_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__o21ba_1
XFILLER_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12870_ rbzero.wall_tracer.visualWallDist\[0\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05607_ sky130_fd_sc_hd__a21o_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ rbzero.tex_g1\[55\] rbzero.tex_g1\[54\] _04212_ vssd1 vssd1 vccd1 vccd1 _04598_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _07274_ _07275_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__and2_1
XFILLER_42_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _04345_ _04527_ _04528_ _04529_ _04253_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__o221a_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ rbzero.tex_g1\[6\] rbzero.tex_g1\[7\] _03691_ vssd1 vssd1 vccd1 vccd1 _03693_
+ sky130_fd_sc_hd__mux2_1
X_14471_ _07206_ _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__or2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11683_ rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__buf_4
XFILLER_42_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _08377_ _08329_ _08854_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__or3b_1
X_13422_ _05995_ _06113_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__and2_1
XFILLER_186_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ _03656_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__clkbuf_1
X_17190_ rbzero.wall_tracer.mapX\[5\] _05512_ _05527_ vssd1 vssd1 vccd1 vccd1 _09775_
+ sky130_fd_sc_hd__a21o_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _08594_ _08075_ _08784_ _08785_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__o31a_1
X_13353_ _06075_ _06089_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__xnor2_1
X_10565_ rbzero.tex_r0\[8\] rbzero.tex_r0\[7\] _03613_ vssd1 vssd1 vccd1 vccd1 _03620_
+ sky130_fd_sc_hd__mux2_1
X_12304_ _04813_ _04811_ _04006_ _03475_ net20 net21 vssd1 vssd1 vccd1 vccd1 _05073_
+ sky130_fd_sc_hd__mux4_1
X_16072_ _08695_ _08715_ _08716_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__a21oi_2
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ _06001_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__xnor2_1
X_10496_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _03580_ vssd1 vssd1 vccd1 vccd1 _03584_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15023_ _07685_ _07686_ _07687_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__and3b_1
XFILLER_68_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19900_ rbzero.pov.ready_buffer\[47\] _02823_ _03193_ _03203_ vssd1 vssd1 vccd1 vccd1
+ _03204_ sky130_fd_sc_hd__a211o_1
X_12235_ _04154_ _03477_ _04966_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__mux2_1
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19831_ _08000_ _03143_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__nand2_1
X_12166_ net39 _04918_ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a21o_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11117_ _03909_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19762_ _03109_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
X_12097_ net6 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__inv_2
X_16974_ _09514_ _09607_ _09613_ vssd1 vssd1 vccd1 vccd1 _09614_ sky130_fd_sc_hd__a21oi_4
XFILLER_111_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18713_ _02405_ _09819_ rbzero.wall_tracer.trackDistY\[-11\] _02406_ vssd1 vssd1
+ vccd1 vccd1 _00602_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ _03873_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__clkbuf_1
X_15925_ _08084_ vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__buf_4
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19693_ _03073_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__clkbuf_1
Xinput8 i_gpout1_sel[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_6
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20168__195 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__inv_2
XFILLER_92_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15856_ _08499_ _08500_ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__and2_1
X_18644_ _02335_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__03293_ _03293_ vssd1 vssd1 vccd1 vccd1 clknet_0__03293_ sky130_fd_sc_hd__clkbuf_16
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ rbzero.wall_tracer.stepDistY\[-5\] _07461_ vssd1 vssd1 vccd1 vccd1 _07537_
+ sky130_fd_sc_hd__nor2_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15787_ _08430_ _08431_ vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__nor2_1
X_18575_ _02146_ _02148_ _02145_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a21bo_1
XFILLER_75_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _05687_ _05719_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__or2_2
XFILLER_205_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14738_ _05844_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__buf_2
X_17526_ _09975_ _09985_ _10091_ vssd1 vssd1 vccd1 vccd1 _10092_ sky130_fd_sc_hd__a21oi_2
XFILLER_75_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17457_ _09730_ _09732_ vssd1 vssd1 vccd1 vccd1 _10024_ sky130_fd_sc_hd__nor2_1
X_14669_ _07376_ _07392_ _07405_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__or3_1
XFILLER_33_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16408_ _09050_ _09052_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__xor2_2
X_17388_ _09919_ _09954_ vssd1 vssd1 vccd1 vccd1 _09955_ sky130_fd_sc_hd__xnor2_2
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19127_ _02698_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__clkbuf_1
X_16339_ _05194_ _08982_ _08983_ _08224_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__a31o_1
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19058_ _02661_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18009_ _01581_ _01585_ _01583_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a21boi_1
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21020_ clknet_leaf_69_i_clk _00789_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20385__11 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
XFILLER_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20804_ clknet_leaf_17_i_clk _00573_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20735_ clknet_leaf_91_i_clk _00504_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20666_ clknet_leaf_25_i_clk _00450_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20597_ _02827_ _02836_ _02835_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a21oi_1
XFILLER_104_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10350_ _03482_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12020_ _04254_ _04790_ _04794_ _04371_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a211o_1
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21218_ clknet_leaf_71_i_clk _00987_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21149_ clknet_leaf_83_i_clk _00918_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13971_ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15710_ _08354_ _08329_ _08058_ vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__or3_1
X_12922_ _04001_ _05494_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nand2_1
X_16690_ _09332_ _07949_ _07895_ vssd1 vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__mux2_1
XFILLER_100_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _07959_ _07932_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__nor2_1
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ rbzero.wall_tracer.visualWallDist\[-12\] rbzero.wall_tracer.rayAddendY\[-4\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__mux2_1
XFILLER_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _02056_ _02057_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and2_1
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11804_ _04224_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__or2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _08002_ rbzero.wall_tracer.stepDistY\[4\] vssd1 vssd1 vccd1 vccd1 _08217_
+ sky130_fd_sc_hd__and2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12784_ _05526_ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09881_ sky130_fd_sc_hd__nand2_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14523_ _07242_ _07240_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__and2_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18291_ _10248_ _09977_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__nor2_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ rbzero.debug_overlay.playerX\[0\] _04459_ _04460_ rbzero.debug_overlay.playerX\[-2\]
+ _04042_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a221o_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _09812_ _09815_ _09816_ _09817_ _09819_ vssd1 vssd1 vccd1 vccd1 _09820_ sky130_fd_sc_hd__o311a_1
XFILLER_109_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14454_ _07187_ _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__and2_1
XFILLER_175_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11666_ _04435_ _04437_ _04439_ _04440_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o41a_1
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ _06138_ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__xor2_1
XFILLER_168_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20356__365 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__inv_2
XFILLER_179_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17173_ rbzero.traced_texa\[2\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__a22o_1
X_10617_ rbzero.tex_g1\[47\] rbzero.tex_g1\[48\] _03647_ vssd1 vssd1 vccd1 vccd1 _03648_
+ sky130_fd_sc_hd__mux2_1
X_14385_ _06724_ _06708_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__or2_1
X_11597_ rbzero.tex_r1\[61\] rbzero.tex_r1\[60\] _04338_ vssd1 vssd1 vccd1 vccd1 _04376_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16124_ _07980_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__or3_1
X_13336_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__xnor2_2
X_10548_ rbzero.tex_r0\[16\] rbzero.tex_r0\[15\] _03602_ vssd1 vssd1 vccd1 vccd1 _03611_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16055_ _08679_ _08699_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__xnor2_1
X_13267_ _05983_ _05981_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__or3_1
X_10479_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _03569_ vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15006_ _07673_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__clkbuf_1
X_12218_ _04886_ _04887_ _04961_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__mux2_1
XFILLER_130_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13198_ _05778_ _05934_ _05928_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__o21a_1
XFILLER_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19814_ rbzero.pov.ready _02821_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__and2_1
X_12149_ net50 _04907_ _04910_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a31o_1
XFILLER_111_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03314_ clknet_0__03314_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03314_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19745_ _03100_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
X_16957_ rbzero.debug_overlay.playerY\[-2\] rbzero.debug_overlay.playerX\[-2\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09598_ sky130_fd_sc_hd__mux2_1
XFILLER_110_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15908_ _07988_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__or3_1
X_19676_ _03064_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16888_ _08204_ _08570_ vssd1 vssd1 vccd1 vccd1 _09529_ sky130_fd_sc_hd__nor2_1
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18627_ _02291_ _02300_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__or2b_1
XFILLER_53_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _08480_ _08481_ _08483_ vssd1 vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__a21bo_1
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18558_ _10239_ _09481_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _09522_ _08151_ _10074_ vssd1 vssd1 vccd1 vccd1 _10075_ sky130_fd_sc_hd__or3_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18489_ _01860_ _09141_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__or4_1
XFILLER_127_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_13 _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20520_ _03413_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 _09762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_46 _09458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20451_ rbzero.texV\[-6\] _03175_ _03332_ _03356_ vssd1 vssd1 vccd1 vccd1 _01390_
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20382_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__buf_1
XFILLER_173_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21003_ clknet_leaf_50_i_clk _00772_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20383__9 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11520_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _04263_ vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__mux2_1
XFILLER_169_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20718_ clknet_leaf_9_i_clk _00008_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11451_ _04223_ _04227_ _04228_ _04219_ _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__o221a_1
XFILLER_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20649_ clknet_leaf_6_i_clk _00433_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10402_ _03532_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14170_ _06905_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__nor2_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11382_ rbzero.row_render.size\[3\] vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__inv_2
XFILLER_180_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13121_ _05761_ _05762_ _05796_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__mux2_1
XFILLER_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10333_ _03496_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13052_ _05694_ _05771_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nand2_1
XFILLER_124_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12003_ _04774_ _04777_ _04332_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__mux2_1
X_17860_ _01461_ _01470_ _01468_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a21o_1
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16811_ _09321_ _09323_ _09452_ vssd1 vssd1 vccd1 vccd1 _09453_ sky130_fd_sc_hd__o21a_1
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17791_ _10258_ _10262_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__and2_1
X_19530_ _04034_ _03006_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__or2_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13954_ _06689_ _06690_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__or2_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16742_ _09269_ _09273_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__or2_1
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12905_ _05609_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__xor2_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19461_ _02916_ _02929_ _02930_ _02911_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_74_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16673_ _09311_ _09312_ _09314_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__a21oi_1
X_13885_ _05978_ _06067_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__or2_1
XFILLER_47_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18412_ _02109_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__or2_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ rbzero.wall_tracer.visualWallDist\[9\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05573_ sky130_fd_sc_hd__a21o_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ rbzero.wall_tracer.stepDistX\[-1\] vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__clkinv_2
XFILLER_50_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _02868_ _02871_ _02869_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a21bo_1
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18343_ _09141_ _01620_ _02041_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__or3_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ rbzero.wall_tracer.stepDistY\[0\] vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__inv_2
XFILLER_187_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12767_ rbzero.map_rom.f1 _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__or2_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14506_ _07237_ _07240_ _07242_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__a21boi_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18274_ _01646_ _01883_ _10271_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a21oi_1
X_11718_ _04480_ _04490_ _04492_ _04496_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__o22a_1
XFILLER_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15486_ _08127_ _08130_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__nor2_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _05416_ _05442_ _05443_ _05444_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a311o_1
XFILLER_187_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14437_ _07110_ _07173_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__xnor2_1
X_17225_ _08937_ _09803_ vssd1 vssd1 vccd1 vccd1 _09804_ sky130_fd_sc_hd__xor2_1
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput11 i_gpout1_sel[3] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_4
X_11649_ _04422_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nor2_1
Xinput22 i_gpout3_sel[2] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_6
Xinput33 i_gpout5_sel[1] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_2
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 i_reset_lock_a vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_4
X_17156_ _07679_ vssd1 vssd1 vccd1 vccd1 _09767_ sky130_fd_sc_hd__buf_2
X_14368_ _07104_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__inv_2
XFILLER_196_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _08743_ _08750_ _08751_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__a21oi_1
X_13319_ _05922_ _06054_ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a21o_1
XFILLER_157_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17087_ _09579_ _09581_ vssd1 vssd1 vccd1 vccd1 _09727_ sky130_fd_sc_hd__and2b_1
XFILLER_196_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14299_ _06842_ _06881_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__xor2_1
XFILLER_66_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16038_ _08680_ _08681_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17989_ _01688_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nand2_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19728_ _03091_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19659_ _03055_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21621_ clknet_leaf_20_i_clk _01390_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21552_ net473 _01321_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20503_ _09750_ _03399_ _03400_ _03250_ rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1
+ _01398_ sky130_fd_sc_hd__a32o_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21483_ net404 _01252_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20434_ rbzero.texV\[-9\] _03175_ _03332_ _03342_ vssd1 vssd1 vccd1 vccd1 _01387_
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ rbzero.tex_b1\[16\] rbzero.tex_b1\[17\] _03817_ vssd1 vssd1 vccd1 vccd1 _03823_
+ sky130_fd_sc_hd__mux2_1
XFILLER_112_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ _06406_ _06078_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__or2_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10882_ rbzero.tex_b1\[49\] rbzero.tex_b1\[50\] _03784_ vssd1 vssd1 vccd1 vccd1 _03787_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ rbzero.map_rom.c6 _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__and2_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15340_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _05304_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__nor2_1
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _04273_ vssd1 vssd1 vccd1 vccd1 _04283_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15271_ _05495_ _07914_ _07915_ _05195_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__o211a_2
XFILLER_184_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12483_ rbzero.wall_tracer.trackDistX\[-7\] vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__inv_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03317_ clknet_0__03317_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03317_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17010_ _09647_ _09649_ vssd1 vssd1 vccd1 vccd1 _09650_ sky130_fd_sc_hd__nor2_1
X_14222_ _06955_ _06957_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__nand2_1
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14153_ _06741_ _06888_ _06889_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a21bo_1
X_11365_ _04141_ _04142_ _04143_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__or4_1
XFILLER_99_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ _05634_ _05636_ _05796_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__mux2_1
XFILLER_153_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10316_ _03487_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14084_ _06799_ _06814_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18961_ _02610_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__clkbuf_1
X_11296_ _04073_ _04072_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__nand2_1
XFILLER_106_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13035_ _05760_ _05763_ _05767_ _05769_ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o2111ai_2
X_17912_ _01516_ _01522_ _01614_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a21oi_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18892_ _02561_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__or3b_1
XFILLER_121_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17843_ _01442_ _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17774_ _08202_ _01476_ _08417_ _08445_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14986_ _00008_ _07552_ _07663_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19513_ _02973_ _02979_ _02989_ _03913_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a31o_1
X_16725_ _09365_ _09366_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__nand2_1
X_13937_ _06161_ _06667_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__nor2_2
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19444_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__or2_1
X_13868_ _06604_ _06554_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__xnor2_2
XFILLER_35_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16656_ _09282_ _09297_ _09298_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__nand3_1
XFILLER_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03044_ _03044_ vssd1 vssd1 vccd1 vccd1 clknet_0__03044_ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12819_ rbzero.wall_tracer.mapY\[10\] _05404_ _05555_ vssd1 vssd1 vccd1 vccd1 _05557_
+ sky130_fd_sc_hd__a21bo_1
X_15607_ _08245_ _08251_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__xor2_2
X_19375_ _02851_ _02855_ _02852_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__o21ai_1
X_13799_ _06057_ _06061_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__nor2_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16587_ _09224_ _09229_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18326_ _01905_ _02013_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__or2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15538_ _08181_ _08182_ _07970_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__a21o_1
XFILLER_124_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15469_ _08111_ _08022_ _08113_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__o21ai_1
X_18257_ _01498_ _08423_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__nor2_1
XFILLER_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17208_ _09779_ _09789_ _09790_ _09781_ rbzero.wall_tracer.mapX\[8\] vssd1 vssd1
+ vccd1 vccd1 _00573_ sky130_fd_sc_hd__a32o_1
XFILLER_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18188_ _01753_ _01769_ _01768_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a21bo_1
XFILLER_190_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _07530_ _09763_ rbzero.row_render.size\[2\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00530_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_143_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20983_ clknet_leaf_50_i_clk _00752_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21604_ net145 _01373_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21535_ net456 _01304_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21466_ net387 _01235_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20417_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03328_
+ sky130_fd_sc_hd__or2_1
X_21397_ net318 _01166_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11150_ _03923_ _03928_ _03932_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or4_2
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _03887_ vssd1 vssd1 vccd1 vccd1 _03891_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ rbzero.wall_tracer.stepDistY\[2\] _07562_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07563_ sky130_fd_sc_hd__mux2_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _05844_ _05952_ _07469_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__and3_1
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11983_ _04755_ _04756_ _04757_ _04247_ _04332_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__o221a_1
XFILLER_57_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13722_ _06427_ _06457_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16510_ _08995_ _08997_ vssd1 vssd1 vccd1 vccd1 _09154_ sky130_fd_sc_hd__nor2_1
XFILLER_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10934_ rbzero.tex_b1\[24\] rbzero.tex_b1\[25\] _03806_ vssd1 vssd1 vccd1 vccd1 _03814_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17490_ _08335_ _09703_ vssd1 vssd1 vccd1 vccd1 _10056_ sky130_fd_sc_hd__and2_1
XFILLER_186_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13653_ _06283_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__and2_1
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16441_ rbzero.wall_tracer.texu\[0\] _09085_ vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__or2_1
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ rbzero.tex_b1\[57\] rbzero.tex_b1\[58\] _03773_ vssd1 vssd1 vccd1 vccd1 _03778_
+ sky130_fd_sc_hd__mux2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _05289_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__nand2_1
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _09013_ _09015_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__and2_1
X_19160_ _05189_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__buf_6
X_13584_ _06308_ _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _03740_ vssd1 vssd1 vccd1 vccd1 _03742_
+ sky130_fd_sc_hd__mux2_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _07959_ _07967_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__nor2_1
X_18111_ _01807_ _01810_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__or2_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12535_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or2_2
XFILLER_200_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19091_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.spi_buffer\[0\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15254_ rbzero.debug_overlay.playerX\[-6\] _07897_ vssd1 vssd1 vccd1 vccd1 _07899_
+ sky130_fd_sc_hd__nand2_1
X_18042_ _09668_ _09693_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nor2_1
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ rbzero.wall_tracer.trackDistY\[7\] _05218_ _05220_ rbzero.wall_tracer.trackDistX\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14205_ _06664_ _06940_ _06941_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__a21oi_1
X_11417_ _04022_ _04187_ _04186_ gpout0.hpos\[5\] _04196_ vssd1 vssd1 vccd1 vccd1
+ _04197_ sky130_fd_sc_hd__o221a_1
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15185_ _07837_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__xnor2_1
X_12397_ _05157_ _05160_ _05163_ net34 net35 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a32o_1
XFILLER_158_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14136_ _06861_ _06871_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__nand2_1
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11348_ _04088_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nand2_2
XFILLER_158_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19993_ rbzero.pov.ready_buffer\[19\] _03252_ _03253_ _07730_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01034_ sky130_fd_sc_hd__o221a_1
XFILLER_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14067_ _06769_ _06707_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__or2_1
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18944_ _02601_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__clkbuf_1
X_11279_ _04057_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__nand2_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13018_ _05743_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__or2_1
X_18875_ _02546_ _02547_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17826_ _01523_ _01529_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17757_ _01459_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ _07654_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16708_ rbzero.wall_tracer.visualWallDist\[9\] _04015_ vssd1 vssd1 vccd1 vccd1 _09350_
+ sky130_fd_sc_hd__nand2_2
X_17688_ _10236_ _10252_ vssd1 vssd1 vccd1 vccd1 _10253_ sky130_fd_sc_hd__xor2_1
XFILLER_90_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19427_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.debug_overlay.vplaneY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__nor2_1
X_16639_ _09277_ _09281_ vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__xor2_1
X_20221__243 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__inv_2
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19358_ _07703_ _02846_ _02847_ _07706_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__a31o_1
XFILLER_128_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18309_ _02006_ _02008_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19289_ rbzero.spi_registers.got_new_leak _02730_ _02728_ _02799_ vssd1 vssd1 vccd1
+ vccd1 _00785_ sky130_fd_sc_hd__a31o_1
XFILLER_202_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21320_ net241 _01089_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21251_ clknet_leaf_79_i_clk _01020_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21182_ clknet_leaf_70_i_clk _00951_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20304__318 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__inv_2
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ clknet_leaf_68_i_clk _00735_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20897_ clknet_leaf_84_i_clk _00666_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_201_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10650_ rbzero.tex_g1\[31\] rbzero.tex_g1\[32\] _03658_ vssd1 vssd1 vccd1 vccd1 _03665_
+ sky130_fd_sc_hd__mux2_1
X_20196__220 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__inv_2
XFILLER_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10581_ _03628_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _05087_ _04666_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__nand2_1
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21518_ net439 _01287_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12251_ _04325_ _04965_ _04976_ _05020_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__o2bb2a_2
XFILLER_107_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21449_ net370 _01218_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ _03924_ _03925_ rbzero.map_rom.a6 rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1
+ _03991_ sky130_fd_sc_hd__o22a_1
XFILLER_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _04948_ _04952_ net12 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__o21ai_1
XFILLER_107_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11133_ rbzero.debug_overlay.playerX\[0\] _03919_ _03921_ rbzero.debug_overlay.playerY\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16990_ _09628_ _09629_ vssd1 vssd1 vccd1 vccd1 _09630_ sky130_fd_sc_hd__and2b_1
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ _08535_ _08536_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__xnor2_1
X_11064_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _03876_ vssd1 vssd1 vccd1 vccd1 _03882_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18660_ _01498_ _01860_ _09027_ _09350_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__or4_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _08448_ _08516_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__xor2_4
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _10031_ _10033_ _10174_ _10175_ vssd1 vssd1 vccd1 vccd1 _10177_ sky130_fd_sc_hd__o211ai_2
XFILLER_92_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ rbzero.wall_tracer.stepDistY\[-2\] _07461_ vssd1 vssd1 vccd1 vccd1 _07550_
+ sky130_fd_sc_hd__nor2_1
XFILLER_188_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _02250_ _02287_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__xor2_1
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17542_ _10092_ _10107_ vssd1 vssd1 vccd1 vccd1 _10108_ sky130_fd_sc_hd__xor2_1
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14754_ _05794_ _07104_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__nor2_1
X_11966_ _04739_ _04740_ _04329_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__mux2_1
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13705_ _06402_ _06403_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__xnor2_1
X_10917_ rbzero.tex_b1\[32\] rbzero.tex_b1\[33\] _03795_ vssd1 vssd1 vccd1 vccd1 _03805_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14685_ _07394_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nand2_1
X_17473_ _09908_ _09917_ _09915_ vssd1 vssd1 vccd1 vccd1 _10039_ sky130_fd_sc_hd__a21o_1
XFILLER_205_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ rbzero.tex_b0\[10\] _04213_ _04329_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a21o_1
XFILLER_204_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19212_ rbzero.color_floor\[1\] _02751_ _02754_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__a21o_1
X_13636_ _06349_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__xnor2_2
XFILLER_189_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16424_ _08951_ _08953_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__xor2_4
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10848_ rbzero.tex_g0\[2\] rbzero.tex_g0\[1\] _03762_ vssd1 vssd1 vccd1 vccd1 _03769_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19143_ _02709_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__buf_2
X_13567_ _06111_ _06128_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__xnor2_2
X_16355_ _08358_ _08365_ _08999_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__a21o_1
XFILLER_73_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10779_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _03729_ vssd1 vssd1 vccd1 vccd1 _03733_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12518_ _05272_ _05253_ _05261_ _05262_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a211o_1
X_15306_ _07904_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__buf_4
XFILLER_185_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19074_ _02669_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__clkbuf_1
X_16286_ _08909_ _08853_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__or2b_1
X_13498_ _06168_ _06208_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a21o_1
XFILLER_173_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18025_ _01724_ _01725_ _01716_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15237_ _07881_ _07868_ _07872_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__and3b_1
X_12449_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__buf_6
XFILLER_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15168_ _07818_ _07819_ _07822_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__and3_1
XFILLER_119_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14119_ _06855_ _06699_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__and2b_1
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15099_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__nand2_1
X_19976_ rbzero.pov.ready_buffer\[27\] _03240_ _03243_ rbzero.debug_overlay.facingY\[-4\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__o221a_1
XFILLER_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18927_ _02591_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18858_ _02530_ _02531_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17809_ _01494_ _01512_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__xor2_2
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18789_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__and2_1
XFILLER_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20820_ clknet_leaf_6_i_clk _00589_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20751_ clknet_leaf_39_i_clk _00520_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_211_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20682_ clknet_leaf_2_i_clk _00466_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[11\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_195_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21303_ net224 _01072_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21234_ clknet_leaf_69_i_clk _01003_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21165_ clknet_leaf_63_i_clk _00934_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20116_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__buf_1
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21096_ net186 _00865_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20047_ _04990_ _04322_ _03275_ _03911_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a31o_1
XFILLER_74_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20228__249 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__inv_2
XFILLER_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11820_ _04595_ _04596_ _04345_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__mux2_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ rbzero.tex_g0\[10\] _04212_ _04217_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a21o_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ clknet_leaf_58_i_clk _00718_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _03692_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14470_ _07131_ _07205_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__and2_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ rbzero.debug_overlay.vplaneX\[0\] _04459_ _04460_ rbzero.debug_overlay.vplaneX\[-2\]
+ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a221o_1
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13421_ _06002_ _05976_ _06004_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a21bo_1
X_10633_ rbzero.tex_g1\[39\] rbzero.tex_g1\[40\] _03647_ vssd1 vssd1 vccd1 vccd1 _03656_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ _08674_ _08112_ _08747_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__or3_1
X_13352_ _06077_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10564_ _03619_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12303_ net23 net22 _05071_ net24 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a31o_1
X_16071_ _08696_ _08714_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__nor2_1
X_13283_ _06006_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__xnor2_1
X_10495_ _03583_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15022_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_1
X_12234_ net17 net16 _05003_ net18 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a31o_1
XFILLER_170_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19830_ rbzero.pov.ready_buffer\[61\] _07999_ _03146_ vssd1 vssd1 vccd1 vccd1 _03150_
+ sky130_fd_sc_hd__mux2_1
X_12165_ net48 _04903_ _04922_ net40 _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_1
XFILLER_64_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11116_ rbzero.tex_b0\[2\] rbzero.tex_b0\[1\] _03557_ vssd1 vssd1 vccd1 vccd1 _03909_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19761_ rbzero.pov.spi_buffer\[54\] rbzero.pov.spi_buffer\[55\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
X_12096_ _04867_ _04837_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__and2_1
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16973_ _09609_ _09612_ vssd1 vssd1 vccd1 vccd1 _09613_ sky130_fd_sc_hd__xnor2_2
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18712_ _02398_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__clkbuf_4
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _03865_ vssd1 vssd1 vccd1 vccd1 _03873_
+ sky130_fd_sc_hd__mux2_1
X_15924_ _08497_ _08501_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__xnor2_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19692_ rbzero.pov.spi_buffer\[21\] rbzero.pov.spi_buffer\[22\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 i_gpout1_sel[1] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_6
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03292_ _03292_ vssd1 vssd1 vccd1 vccd1 clknet_0__03292_ sky130_fd_sc_hd__clkbuf_16
X_18643_ _08418_ _02336_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _08109_ _08042_ _08125_ _08084_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__o22ai_1
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14806_ _07487_ _07456_ _07533_ _07535_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__a211oi_4
XFILLER_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18574_ _02188_ _02190_ _02187_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a21bo_1
XFILLER_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _08330_ _08415_ _08429_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__a21oi_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _05721_ _05734_ _05707_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__or3_1
XFILLER_75_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17525_ _09979_ _09984_ vssd1 vssd1 vccd1 vccd1 _10091_ sky130_fd_sc_hd__and2_1
X_14737_ _05844_ _07471_ _06239_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__a21o_1
X_11949_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _04356_ vssd1 vssd1 vccd1 vccd1 _04725_
+ sky130_fd_sc_hd__mux2_1
XFILLER_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17456_ _09614_ _10022_ vssd1 vssd1 vccd1 vccd1 _10023_ sky130_fd_sc_hd__xnor2_4
XFILLER_178_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14668_ _07394_ _07399_ _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__or3b_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16407_ _08412_ _08438_ _09051_ vssd1 vssd1 vccd1 vccd1 _09052_ sky130_fd_sc_hd__a21oi_2
XFILLER_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13619_ _05823_ _05920_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__or2_1
X_17387_ _09952_ _09953_ vssd1 vssd1 vccd1 vccd1 _09954_ sky130_fd_sc_hd__nand2_1
X_14599_ _07218_ _07323_ _07331_ _07216_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a211o_1
XFILLER_192_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19126_ net41 rbzero.spi_registers.ss_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02698_ sky130_fd_sc_hd__mux2_1
XFILLER_203_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16338_ _07566_ _07568_ _07571_ _08220_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__or4_2
XFILLER_173_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19057_ rbzero.pov.spi_buffer\[59\] rbzero.pov.ready_buffer\[59\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
X_16269_ _08250_ _08331_ _08862_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__a21oi_1
X_20333__344 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__inv_2
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18008_ _01708_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__nand2_1
XFILLER_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19959_ _03246_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__buf_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20803_ clknet_leaf_17_i_clk _00572_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20734_ clknet_leaf_91_i_clk _00503_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_81_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20665_ clknet_leaf_25_i_clk _00449_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20596_ rbzero.wall_tracer.rayAddendY\[-7\] _03443_ _07756_ _03461_ vssd1 vssd1 vccd1
+ vccd1 _01430_ sky130_fd_sc_hd__a22o_1
XFILLER_104_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21217_ clknet_leaf_71_i_clk _00986_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21148_ clknet_leaf_83_i_clk _00917_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20058__96 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__inv_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13970_ _06614_ _06706_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__nand2_2
X_21079_ net169 _00848_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12921_ _05567_ _05576_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__nor2_1
XFILLER_98_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15640_ _08282_ _08283_ _08284_ _07996_ vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__o22ai_2
XFILLER_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ rbzero.wall_tracer.rayAddendX\[-2\] _05588_ _05560_ vssd1 vssd1 vccd1 vccd1
+ _05589_ sky130_fd_sc_hd__mux2_2
X_19620__73 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _04341_ vssd1 vssd1 vccd1 vccd1 _04581_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _08214_ _08215_ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__nor2_1
X_12783_ _05513_ _05519_ _05520_ _05512_ rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1
+ vccd1 _05527_ sky130_fd_sc_hd__a32o_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09880_ sky130_fd_sc_hd__or2_1
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14522_ _07258_ _07053_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__xnor2_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ rbzero.debug_overlay.playerX\[-8\] _04466_ _04499_ rbzero.debug_overlay.playerX\[4\]
+ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__a221o_1
XFILLER_199_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18290_ _01988_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_49_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17241_ _08940_ _08943_ _09818_ vssd1 vssd1 vccd1 vccd1 _09819_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14453_ _07188_ _07189_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__and2b_1
X_11665_ gpout0.hpos\[8\] _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and2_1
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13404_ _06139_ _06140_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10616_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__clkbuf_4
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14384_ _06696_ _06740_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__or2_1
X_17172_ rbzero.traced_texa\[1\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a22o_1
X_11596_ rbzero.tex_r1\[63\] rbzero.tex_r1\[62\] _04338_ vssd1 vssd1 vccd1 vccd1 _04375_
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13335_ _06059_ _06060_ _06045_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16123_ _08008_ _08128_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__or2_1
X_10547_ _03610_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13266_ _06002_ _05976_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16054_ _08676_ _08677_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__xor2_1
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10478_ _03574_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12217_ _04883_ _04884_ _04966_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__mux2_1
X_15005_ rbzero.wall_tracer.stepDistX\[9\] _07582_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07673_ sky130_fd_sc_hd__mux2_1
XFILLER_68_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13197_ _05867_ _05688_ _05801_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__mux2_1
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19813_ _03135_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ net49 _04903_ _04918_ net52 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a22o_1
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03313_ clknet_0__03313_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03313_
+ sky130_fd_sc_hd__clkbuf_16
X_19744_ rbzero.pov.spi_buffer\[46\] rbzero.pov.spi_buffer\[47\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
X_12079_ net5 _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nor2_1
X_16956_ _09594_ _09596_ vssd1 vssd1 vccd1 vccd1 _09597_ sky130_fd_sc_hd__xor2_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15907_ _08551_ _08481_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__xor2_1
X_19675_ rbzero.pov.spi_buffer\[13\] rbzero.pov.spi_buffer\[14\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16887_ _09525_ _09527_ vssd1 vssd1 vccd1 vccd1 _09528_ sky130_fd_sc_hd__and2_1
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18626_ _02316_ _02322_ rbzero.wall_tracer.trackDistX\[10\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00599_ sky130_fd_sc_hd__o2bb2a_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _07923_ _07967_ _08482_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__or3_1
XFILLER_53_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18557_ _02144_ _02158_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a21bo_1
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15769_ _08408_ _08402_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__or2b_1
XFILLER_178_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17508_ _07974_ _08158_ vssd1 vssd1 vccd1 vccd1 _10074_ sky130_fd_sc_hd__or2_1
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18488_ _02039_ _02042_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__nand2_1
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17439_ _10003_ _10005_ vssd1 vssd1 vccd1 vccd1 _10006_ sky130_fd_sc_hd__xnor2_2
XANTENNA_14 _08008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_25 _09859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_36 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_47 _10027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20450_ _03353_ _03355_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19109_ rbzero.spi_registers.spi_buffer\[10\] rbzero.spi_registers.spi_buffer\[9\]
+ _02676_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21002_ clknet_leaf_51_i_clk _00771_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_sky
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20717_ clknet_leaf_16_i_clk _00007_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11450_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__buf_4
XFILLER_149_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20648_ clknet_leaf_5_i_clk _00432_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10401_ rbzero.tex_r1\[19\] rbzero.tex_r1\[20\] _03527_ vssd1 vssd1 vccd1 vccd1 _03532_
+ sky130_fd_sc_hd__mux2_1
X_11381_ rbzero.row_render.size\[4\] vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__inv_2
X_20579_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__or2_1
XFILLER_137_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _05690_ _05801_ _05817_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__o21ai_1
XFILLER_139_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ rbzero.tex_r1\[52\] rbzero.tex_r1\[53\] _03494_ vssd1 vssd1 vccd1 vccd1 _03496_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13051_ _05780_ _05746_ _05782_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nand4_2
XFILLER_106_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12002_ _04775_ _04776_ _04218_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__mux2_1
XFILLER_191_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16810_ _09318_ _09320_ vssd1 vssd1 vccd1 vccd1 _09452_ sky130_fd_sc_hd__or2_1
XFILLER_121_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17790_ _10243_ _10251_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__a21o_1
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16741_ _09251_ _09261_ _09259_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__a21o_1
XFILLER_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13953_ _06610_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__buf_2
XFILLER_207_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12904_ _05562_ _05566_ _05619_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__and3_1
XFILLER_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19460_ _02940_ _02941_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__nor2_1
XFILLER_207_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20362__370 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__inv_2
X_16672_ _09311_ _09312_ _09314_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__and3_1
X_13884_ _06201_ _06052_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__nor2_1
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18411_ _01946_ _01949_ _02108_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__and3_1
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15623_ _08191_ _08265_ _08267_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__a21bo_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _07728_ _02872_ _02877_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__a21o_1
X_12835_ _04031_ _05327_ _05371_ _04001_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a31o_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _02039_ _02040_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__nand2_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _08196_ _08198_ _07951_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__a21o_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _05496_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__buf_2
XFILLER_203_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _07238_ _07241_ _07239_ _07075_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__a22o_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18273_ _01646_ _01972_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__xnor2_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ rbzero.debug_overlay.facingX\[10\] _04453_ _04493_ _04495_ vssd1 vssd1 vccd1
+ vccd1 _04496_ sky130_fd_sc_hd__a211o_1
X_15485_ _08047_ _08124_ _08128_ _08129_ vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__o22a_1
X_12697_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__xnor2_2
XFILLER_203_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ _08939_ _08851_ vssd1 vssd1 vccd1 vccd1 _09803_ sky130_fd_sc_hd__and2_1
XFILLER_187_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14436_ _06689_ _06760_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__nor2_1
X_11648_ gpout0.hpos\[5\] _04424_ _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__or3_1
XFILLER_128_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 i_gpout1_sel[4] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_4
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 i_gpout3_sel[3] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_6
Xinput34 i_gpout5_sel[2] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_8
Xinput45 i_reset_lock_b vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_4
X_17155_ rbzero.row_render.texu\[5\] _09766_ _07728_ rbzero.wall_tracer.texu\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__a22o_1
X_11579_ rbzero.tex_r1\[17\] rbzero.tex_r1\[16\] _04290_ vssd1 vssd1 vccd1 vccd1 _04358_
+ sky130_fd_sc_hd__mux2_1
X_14367_ _05779_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__or2_1
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16106_ _08744_ _08749_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__nor2_1
X_13318_ _05973_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__inv_2
XFILLER_183_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14298_ _06882_ _07034_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__and2_1
X_17086_ _09657_ _09725_ vssd1 vssd1 vccd1 vccd1 _09726_ sky130_fd_sc_hd__xnor2_2
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16037_ _08680_ _08681_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__or2_1
X_13249_ _05962_ _05976_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a21o_1
XFILLER_171_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17988_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__inv_2
XFILLER_81_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19727_ rbzero.pov.spi_buffer\[38\] rbzero.pov.spi_buffer\[39\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16939_ _09442_ _09443_ vssd1 vssd1 vccd1 vccd1 _09580_ sky130_fd_sc_hd__nor2_1
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19658_ rbzero.pov.spi_buffer\[5\] rbzero.pov.spi_buffer\[6\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_129_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ _02109_ _02213_ _02211_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21620_ clknet_leaf_33_i_clk _01389_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21551_ net472 _01320_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20502_ _03395_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__a21o_1
XFILLER_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21482_ net403 _01251_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20433_ _03340_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__xnor2_1
X_20190__215 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__inv_2
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10950_ _03822_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10881_ _03786_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__buf_2
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__and2_1
XFILLER_106_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11502_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _04273_ vssd1 vssd1 vccd1 vccd1 _04282_
+ sky130_fd_sc_hd__mux2_1
XFILLER_169_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12482_ rbzero.wall_tracer.trackDistX\[-6\] vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__inv_2
X_15270_ rbzero.debug_overlay.playerX\[-5\] _05495_ vssd1 vssd1 vccd1 vccd1 _07915_
+ sky130_fd_sc_hd__nand2_1
XFILLER_196_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03316_ clknet_0__03316_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03316_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14221_ _06955_ _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__nor2_1
X_11433_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__buf_4
XFILLER_138_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _05825_ _06740_ _06678_ _06704_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__o22ai_1
X_11364_ _03476_ _04025_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o21ba_4
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13103_ _05838_ _05839_ _05811_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__mux2_1
XFILLER_152_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10315_ rbzero.tex_r1\[60\] rbzero.tex_r1\[61\] _03483_ vssd1 vssd1 vccd1 vccd1 _03487_
+ sky130_fd_sc_hd__mux2_1
X_14083_ _06703_ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__nor2_1
X_18960_ rbzero.pov.spi_buffer\[13\] rbzero.pov.ready_buffer\[13\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XFILLER_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11295_ _04071_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nor2_1
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13034_ _05701_ _05702_ _05683_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__or4_1
X_17911_ _01517_ _01521_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__and2_1
XFILLER_152_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18891_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] vssd1
+ vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__or2_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17842_ _01543_ _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17773_ _01474_ _08202_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__or4_1
X_14985_ rbzero.wall_tracer.stepDistX\[-1\] _07650_ vssd1 vssd1 vccd1 vccd1 _07663_
+ sky130_fd_sc_hd__nor2_1
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19512_ _02973_ _02979_ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a21oi_1
X_16724_ _08821_ _08159_ _08151_ _09243_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__o22ai_1
X_13936_ _06245_ _06672_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__nor2_1
XFILLER_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19443_ _02923_ _02924_ _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__o211a_1
XFILLER_90_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16655_ _09291_ _09293_ _09296_ vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__a21o_1
X_13867_ _06464_ _06552_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__nand2_1
XFILLER_35_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03043_ _03043_ vssd1 vssd1 vccd1 vccd1 clknet_0__03043_ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15606_ _08217_ _08225_ _08250_ vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__o21a_1
X_19374_ _02860_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__nand2_1
X_12818_ _05533_ _05555_ _05556_ _05284_ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1
+ vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
XFILLER_90_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16586_ _09227_ _09228_ vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__xor2_1
X_13798_ _05877_ _05888_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nor2_1
XFILLER_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18325_ _01801_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__and2_1
XFILLER_176_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _07560_ _08171_ _07562_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__o21ai_1
XFILLER_163_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12749_ _03924_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18256_ _01954_ _01955_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__nand2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15468_ _08084_ _08112_ _08103_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__or3_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ _09783_ _09787_ _09788_ vssd1 vssd1 vccd1 vccd1 _09790_ sky130_fd_sc_hd__o21ai_1
X_14419_ _07154_ _07155_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__or2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18187_ _01885_ _01886_ _01876_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a21o_1
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15399_ rbzero.wall_tracer.visualWallDist\[1\] _07925_ vssd1 vssd1 vccd1 vccd1 _08044_
+ sky130_fd_sc_hd__nand2_8
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17138_ _07524_ _09763_ rbzero.row_render.size\[1\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00529_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17069_ _09707_ _09708_ vssd1 vssd1 vccd1 vccd1 _09709_ sky130_fd_sc_hd__xnor2_2
XFILLER_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20982_ clknet_leaf_52_i_clk _00751_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21603_ net144 _01372_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21534_ net455 _01303_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21465_ net386 _01234_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20416_ _03272_ _03325_ _03326_ _03327_ rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1
+ _01384_ sky130_fd_sc_hd__a32o_1
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21396_ net317 _01165_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ _03890_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ _07503_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _04291_ vssd1 vssd1 vccd1 vccd1 _04757_
+ sky130_fd_sc_hd__mux2_1
XFILLER_112_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13721_ _06427_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__or2b_1
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10933_ _03813_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16440_ _07970_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__buf_4
X_13652_ _05824_ _06080_ _06282_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__o21ai_1
X_10864_ _03777_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__nand2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _09013_ _09015_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__nor2_1
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13583_ _06316_ _06318_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a21o_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10795_ _03741_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18110_ _01807_ _01810_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__nand2_1
XFILLER_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _07966_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _02678_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__clkbuf_1
X_12534_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] _05286_
+ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a31o_1
XFILLER_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _01741_ _01742_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__xnor2_2
X_15253_ rbzero.debug_overlay.playerX\[-6\] _07897_ vssd1 vssd1 vccd1 vccd1 _07898_
+ sky130_fd_sc_hd__or2_1
X_12465_ rbzero.wall_tracer.trackDistY\[6\] vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__inv_2
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_90 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_90/HI zeros[0] sky130_fd_sc_hd__conb_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14204_ _06704_ _06690_ _06663_ _05825_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__o22a_1
X_11416_ gpout0.hpos\[3\] _04189_ _04187_ _04022_ _04195_ vssd1 vssd1 vccd1 vccd1
+ _04196_ sky130_fd_sc_hd__a221o_1
XFILLER_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12396_ net68 _05142_ _05161_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a211o_1
XFILLER_125_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15184_ _07800_ _07812_ _07814_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__a21o_1
XFILLER_153_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14135_ _06861_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__nor2_1
XFILLER_158_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11347_ _04084_ _04087_ _04114_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19992_ rbzero.pov.ready_buffer\[18\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-2\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__a221o_1
XFILLER_125_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14066_ _06787_ _06791_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__xnor2_1
X_11278_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _04058_ sky130_fd_sc_hd__or2_1
X_18943_ rbzero.pov.spi_buffer\[5\] rbzero.pov.ready_buffer\[5\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
X_13017_ _05700_ _05731_ _05746_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__and4bb_2
XFILLER_67_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18874_ _02537_ _02539_ _02538_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a21boi_1
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17825_ _10126_ _01528_ _10271_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a21oi_1
Xhold1 rbzero.tex_r1\[40\] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17756_ _09368_ _09703_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__nand2_1
X_14968_ rbzero.wall_tracer.stepDistX\[-9\] _07502_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07654_ sky130_fd_sc_hd__mux2_1
XFILLER_81_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16707_ _09265_ _09240_ vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__or2b_1
X_13919_ _06639_ _06654_ _06655_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17687_ _10243_ _10251_ vssd1 vssd1 vccd1 vccd1 _10252_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14899_ _07591_ _07606_ _07607_ _04039_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__o211a_1
X_19426_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.debug_overlay.vplaneY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__and2_1
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16638_ _09278_ _09280_ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__xor2_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19357_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__or2_1
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16569_ _08160_ _09165_ _09211_ vssd1 vssd1 vccd1 vccd1 _09212_ sky130_fd_sc_hd__or3b_1
XFILLER_149_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18308_ _01817_ _01896_ _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a21oi_1
X_19288_ _02792_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__inv_2
X_18239_ _10239_ _09027_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__nor2_1
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21250_ clknet_leaf_81_i_clk _01019_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21181_ clknet_leaf_70_i_clk _00950_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20965_ clknet_leaf_68_i_clk _00734_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ clknet_leaf_83_i_clk _00665_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _03624_ vssd1 vssd1 vccd1 vccd1 _03628_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21517_ net438 _01286_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ _04984_ _04995_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__or3b_2
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21448_ net369 _01217_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ rbzero.map_rom.f1 _03942_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2_1
X_12181_ _04907_ _04949_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a21oi_1
X_21379_ net300 _01148_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11132_ rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__inv_2
XFILLER_122_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19627__79 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__inv_2
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15940_ _08539_ _08541_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__xnor2_1
X_11063_ _03881_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15871_ _08199_ _08201_ _08515_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__and3_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17610_ _10174_ _10175_ _10031_ _10033_ vssd1 vssd1 vccd1 vccd1 _10176_ sky130_fd_sc_hd__a211o_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _07486_ _07455_ _07548_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__a21oi_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _02252_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__xor2_1
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17541_ _10098_ _10106_ vssd1 vssd1 vccd1 vccd1 _10107_ sky130_fd_sc_hd__xnor2_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _07486_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__buf_4
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _04356_ vssd1 vssd1 vccd1 vccd1 _04740_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ _06405_ _06410_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__xor2_1
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _03804_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17472_ _09614_ _10022_ vssd1 vssd1 vccd1 vccd1 _10038_ sky130_fd_sc_hd__nand2_1
X_14684_ _07419_ _07420_ _05741_ _07106_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__a211o_1
XFILLER_189_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ rbzero.tex_b0\[11\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and3_1
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19211_ rbzero.spi_registers.new_floor\[1\] rbzero.spi_registers.got_new_floor _02711_
+ _03911_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a31o_1
X_16423_ _09067_ _08955_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__xnor2_4
XFILLER_204_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13635_ _06350_ _06370_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__o21a_1
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _03768_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19142_ rbzero.spi_registers.got_new_other _02708_ vssd1 vssd1 vccd1 vccd1 _02709_
+ sky130_fd_sc_hd__and2_1
X_16354_ _08363_ _08364_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__nor2_1
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13566_ _06131_ _06142_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__xnor2_1
XFILLER_197_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _03732_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15305_ _07948_ _07949_ _05496_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__mux2_1
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19073_ rbzero.pov.spi_buffer\[67\] rbzero.pov.ready_buffer\[67\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
X_12517_ _05263_ rbzero.wall_tracer.trackDistY\[-4\] _05252_ rbzero.wall_tracer.trackDistX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16285_ _08922_ _08927_ _08928_ _08929_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__o211a_1
X_13497_ _06209_ _06223_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and2b_1
XFILLER_173_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18024_ _01716_ _01724_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__or3_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15236_ rbzero.wall_tracer.rayAddendX\[8\] rbzero.wall_tracer.rayAddendX\[7\] _05448_
+ _07821_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__or4b_1
X_12448_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__buf_4
XFILLER_173_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ rbzero.wall_tracer.rayAddendX\[4\] rbzero.wall_tracer.rayAddendX\[3\] _07821_
+ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__o21ai_1
X_12379_ _05143_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__buf_2
XFILLER_113_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ _06848_ _06850_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15098_ _07742_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _07757_
+ sky130_fd_sc_hd__or2_1
X_19975_ rbzero.pov.ready_buffer\[26\] _03247_ _03249_ rbzero.debug_overlay.facingY\[-5\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__a221o_1
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14049_ _06742_ _06785_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__xnor2_1
X_18926_ _02589_ _02557_ _02590_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__and3b_1
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _02524_ _02526_ _02525_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a21boi_1
XFILLER_94_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17808_ _01496_ _01511_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__xor2_2
X_18788_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__nor2_1
XFILLER_94_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17739_ _10199_ _10231_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__nand2_1
X_20400__25 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
XFILLER_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20145__175 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__inv_2
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20750_ clknet_3_7_0_i_clk _00519_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__or2_1
XFILLER_211_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20681_ clknet_leaf_1_i_clk _00465_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_189_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21302_ net223 _01071_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21233_ clknet_leaf_68_i_clk _01002_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20310__323 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__inv_2
X_21164_ clknet_leaf_80_i_clk _00933_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21095_ net185 _00864_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20046_ _03283_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11750_ rbzero.tex_g0\[11\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__and3_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ clknet_leaf_66_i_clk _00717_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ rbzero.tex_g1\[7\] rbzero.tex_g1\[8\] _03691_ vssd1 vssd1 vccd1 vccd1 _03692_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _04004_ _04419_ _04450_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__and3_2
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20879_ clknet_leaf_60_i_clk _00648_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_186_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ _05978_ _05942_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__nor2_1
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10632_ _03655_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13351_ _06082_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__xor2_1
X_10563_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _03613_ vssd1 vssd1 vccd1 vccd1 _03619_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _03473_ _05044_ _05046_ _04317_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a221o_1
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16070_ _08696_ _08714_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__nand2_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10494_ rbzero.tex_r0\[42\] rbzero.tex_r0\[41\] _03580_ vssd1 vssd1 vccd1 vccd1 _03583_
+ sky130_fd_sc_hd__mux2_1
X_13282_ _06010_ _06012_ _06014_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a22o_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15021_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__or2_1
X_12233_ _03473_ _04814_ _04317_ _04809_ _04961_ _04960_ vssd1 vssd1 vccd1 vccd1 _05003_
+ sky130_fd_sc_hd__mux4_1
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ net38 _04907_ net8 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__and3_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11115_ _03908_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__clkbuf_1
X_20285__300 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__inv_2
X_12095_ net51 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16972_ _08162_ _09611_ vssd1 vssd1 vccd1 vccd1 _09612_ sky130_fd_sc_hd__and2_1
X_19760_ _03108_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11046_ _03872_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__clkbuf_1
X_15923_ _08566_ _08567_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__nand2_1
X_18711_ _05532_ _02403_ _02404_ _02399_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__o31a_1
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19691_ _03072_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03291_ _03291_ vssd1 vssd1 vccd1 vccd1 clknet_0__03291_ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18642_ _01620_ _09292_ _02239_ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__o31a_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _08084_ _08041_ _08498_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__or3_1
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _07511_ _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__nor2_1
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _02192_ _02185_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__or2b_1
XFILLER_40_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _08330_ _08415_ _08429_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__and3_1
X_12997_ _05589_ _05704_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__xor2_2
XFILLER_188_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17524_ _09963_ _09969_ _10089_ vssd1 vssd1 vccd1 vccd1 _10090_ sky130_fd_sc_hd__a21o_1
X_14736_ _07469_ _07470_ _05952_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__mux2_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11948_ _04254_ _04719_ _04723_ _04371_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a211o_1
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17455_ _10019_ _10021_ vssd1 vssd1 vccd1 vccd1 _10022_ sky130_fd_sc_hd__xor2_4
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _07375_ _07403_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__nand2_1
X_11879_ rbzero.tex_g1\[29\] rbzero.tex_g1\[28\] _04336_ vssd1 vssd1 vccd1 vccd1 _04656_
+ sky130_fd_sc_hd__mux2_1
X_16406_ _08371_ _08411_ vssd1 vssd1 vccd1 vccd1 _09051_ sky130_fd_sc_hd__nor2_1
X_13618_ _06311_ _06314_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17386_ _09920_ _09921_ _09951_ vssd1 vssd1 vccd1 vccd1 _09953_ sky130_fd_sc_hd__nand3_1
X_14598_ _07218_ _07323_ _07334_ _07332_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__a31o_1
XFILLER_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19125_ _02697_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__clkbuf_1
X_16337_ _08218_ _08232_ _08208_ _08981_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__a31o_1
X_13549_ _05975_ _06285_ _05921_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__and3b_1
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19056_ _02593_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__clkbuf_4
X_16268_ _08215_ _08335_ _08856_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__a21o_1
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18007_ _01462_ _09359_ _01707_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__o21ai_1
X_15219_ _07820_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _07870_
+ sky130_fd_sc_hd__nand2_1
XFILLER_99_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16199_ _08836_ _08842_ _08843_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__a21oi_1
XFILLER_142_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19958_ _03245_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18909_ rbzero.spi_registers.spi_counter\[1\] _02576_ vssd1 vssd1 vccd1 vccd1 _02578_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19889_ _03194_ _03193_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__nand2_1
XFILLER_68_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20802_ clknet_leaf_17_i_clk _00571_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20733_ clknet_leaf_91_i_clk _00502_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20664_ clknet_leaf_25_i_clk _00448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20595_ _02833_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21216_ clknet_leaf_72_i_clk _00985_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21147_ clknet_leaf_82_i_clk _00916_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21078_ net168 _00847_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20029_ _09749_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__clkbuf_4
X_12920_ _05567_ _05575_ _05576_ _05656_ _05563_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__o2111a_1
XFILLER_115_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12851_ rbzero.wall_tracer.visualWallDist\[-10\] rbzero.wall_tracer.rayAddendY\[-2\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__mux2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _04253_ _04575_ _04579_ _04119_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a211o_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ rbzero.wall_tracer.visualWallDist\[-10\] _04012_ vssd1 vssd1 vccd1 vccd1
+ _08215_ sky130_fd_sc_hd__nand2_4
X_20280__296 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__inv_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ rbzero.wall_tracer.mapX\[5\] _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__xnor2_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _07254_ _07257_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__xnor2_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ rbzero.debug_overlay.playerX\[5\] _04444_ _04439_ _04452_ rbzero.debug_overlay.playerX\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__a32o_1
XFILLER_187_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _08940_ _08943_ _05204_ vssd1 vssd1 vccd1 vccd1 _09818_ sky130_fd_sc_hd__a21oi_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _07175_ _07180_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__xor2_1
XFILLER_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ _04441_ _04442_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__nor2_1
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ _06069_ _06074_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__xor2_1
X_10615_ _03481_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__buf_4
X_17171_ rbzero.traced_texa\[0\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22o_1
X_14383_ _07115_ _07119_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__xnor2_1
X_20317__329 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__inv_2
X_11595_ _04140_ _04355_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or3_1
XFILLER_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16122_ _08284_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__buf_4
X_13334_ _06053_ _06056_ _06061_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__a21o_1
XFILLER_70_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10546_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _03602_ vssd1 vssd1 vccd1 vccd1 _03610_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ _08640_ _08648_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__xnor2_1
X_13265_ _05945_ _05949_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_4
XFILLER_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10477_ rbzero.tex_r0\[50\] rbzero.tex_r0\[49\] _03569_ vssd1 vssd1 vccd1 vccd1 _03574_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15004_ _07672_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__clkbuf_1
X_12216_ net18 _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nand2_1
X_13196_ _05591_ _05740_ _05931_ _05893_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a41o_1
XFILLER_68_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19812_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] _05189_ vssd1 vssd1
+ vccd1 vccd1 _03135_ sky130_fd_sc_hd__mux2_1
X_12147_ _04907_ net8 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nor2_2
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03312_ clknet_0__03312_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03312_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19743_ _03099_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12078_ net4 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__inv_2
X_16955_ _09207_ _09330_ _09457_ _09595_ vssd1 vssd1 vccd1 vccd1 _09596_ sky130_fd_sc_hd__a31o_2
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11029_ _03863_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__clkbuf_1
X_15906_ _08483_ _08480_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__nand2_1
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19674_ _03063_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__clkbuf_1
X_16886_ _09526_ _08356_ _09524_ vssd1 vssd1 vccd1 vccd1 _09527_ sky130_fd_sc_hd__o21ai_1
X_15837_ _07912_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__or3_1
X_18625_ _09889_ _02321_ _09780_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a21oi_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15768_ _08154_ _08167_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__or2b_1
X_18556_ _02159_ _02143_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__or2b_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14719_ _07455_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__buf_4
X_17507_ _09522_ _08159_ _08151_ _09661_ vssd1 vssd1 vccd1 vccd1 _10073_ sky130_fd_sc_hd__o22ai_1
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18487_ _02088_ _02090_ _02087_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a21bo_1
X_15699_ _08340_ _08341_ _08342_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17438_ _09702_ _09713_ _10004_ vssd1 vssd1 vccd1 vccd1 _10005_ sky130_fd_sc_hd__a21o_1
XFILLER_166_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 _08096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_26 _10171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17369_ _09926_ _09935_ vssd1 vssd1 vccd1 vccd1 _09936_ sky130_fd_sc_hd__nand2_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19108_ _02687_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__clkbuf_1
X_20257__276 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__inv_2
XFILLER_203_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _02651_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21001_ clknet_leaf_52_i_clk _00770_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20716_ clknet_leaf_12_i_clk _00006_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20647_ clknet_leaf_9_i_clk _00431_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10400_ _03531_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11380_ rbzero.row_render.size\[5\] vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__inv_2
XFILLER_109_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20578_ _03450_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _03495_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ _05695_ _05702_ _05785_ _05786_ _05766_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__o311a_1
XFILLER_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _04212_ vssd1 vssd1 vccd1 vccd1 _04776_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16740_ _09348_ _09381_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__xnor2_1
X_13952_ _06245_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12903_ _05615_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__xor2_2
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16671_ _09113_ _09152_ _09313_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__a21o_1
XFILLER_98_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13883_ _06239_ _06245_ _06202_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__or3_1
XFILLER_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18410_ _01946_ _01949_ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a21oi_2
X_15622_ _07981_ _08177_ _08266_ _08264_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19390_ rbzero.wall_tracer.rayAddendY\[-1\] _07706_ _02876_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _02877_ sky130_fd_sc_hd__a22o_1
X_12834_ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__buf_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _10238_ _09294_ _09977_ _01737_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__o22ai_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _08171_ _08197_ _05193_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__o21ai_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _03936_ _05503_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__nor2_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14504_ _06239_ _07071_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__nor2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18272_ _01968_ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__xnor2_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ rbzero.debug_overlay.facingX\[-5\] _04454_ _04455_ rbzero.debug_overlay.facingX\[-7\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a221o_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _08035_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__buf_4
X_12696_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nor2_1
XFILLER_187_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ rbzero.wall_tracer.mapX\[11\] _09781_ _09779_ _09802_ vssd1 vssd1 vccd1 vccd1
+ _00576_ sky130_fd_sc_hd__a22o_1
X_14435_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__dlymetal6s2s_1
X_11647_ _04005_ _04023_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a21o_1
Xinput13 i_gpout1_sel[5] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_4
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17154_ rbzero.row_render.texu\[4\] _09766_ _07728_ rbzero.wall_tracer.texu\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a22o_1
Xinput24 i_gpout3_sel[4] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_4
Xinput35 i_gpout5_sel[3] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_2
X_14366_ _05793_ _07041_ _07102_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a21oi_2
XFILLER_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput46 i_tex_in[0] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_4
X_11578_ rbzero.tex_r1\[19\] rbzero.tex_r1\[18\] _04356_ vssd1 vssd1 vccd1 vccd1 _04357_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16105_ _08744_ _08749_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__xor2_1
X_13317_ _05939_ _05961_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__nor2_1
X_10529_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _03591_ vssd1 vssd1 vccd1 vccd1 _03601_
+ sky130_fd_sc_hd__mux2_1
X_17085_ _09722_ _09724_ vssd1 vssd1 vccd1 vccd1 _09725_ sky130_fd_sc_hd__xor2_2
X_14297_ _07031_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__xor2_2
XFILLER_170_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16036_ _08624_ _08628_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__xnor2_1
X_13248_ _05983_ _05975_ _05984_ _05974_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__o22a_1
XFILLER_131_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ _05695_ _05677_ _05801_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__mux2_1
XFILLER_112_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17987_ _09249_ _01576_ _01579_ _01577_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__o22a_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19726_ _03090_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__clkbuf_1
X_16938_ _09538_ _09578_ vssd1 vssd1 vccd1 vccd1 _09579_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19657_ _03054_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__clkbuf_1
X_19596__51 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
X_16869_ _09507_ _09509_ vssd1 vssd1 vccd1 vccd1 _09510_ sky130_fd_sc_hd__nor2_1
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ _02303_ _02304_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__or2_1
XFILLER_77_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18539_ _02149_ _02156_ _02155_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__o21bai_1
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21550_ net471 _01319_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20501_ _03398_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__inv_2
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21481_ net402 _01250_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20432_ _03333_ _03334_ _03335_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20294_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__buf_1
XFILLER_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ rbzero.tex_b1\[50\] rbzero.tex_b1\[51\] _03784_ vssd1 vssd1 vccd1 vccd1 _03786_
+ sky130_fd_sc_hd__mux2_1
XFILLER_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__nor2_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11501_ _04230_ _04276_ _04280_ _04232_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a211o_1
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ rbzero.wall_tracer.trackDistX\[-5\] vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__inv_2
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03315_ clknet_0__03315_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03315_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14220_ _06923_ _06931_ _06956_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21boi_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__buf_4
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _05825_ _06678_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nor2_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ _04100_ _04114_ _04120_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__nor3_4
XFILLER_180_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13102_ _05710_ _05713_ _05715_ _05687_ _05791_ _05826_ vssd1 vssd1 vccd1 vccd1 _05839_
+ sky130_fd_sc_hd__mux4_1
XFILLER_125_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10314_ _03486_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14082_ _06685_ _06695_ _06702_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__and3_1
XFILLER_152_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11294_ rbzero.texV\[4\] _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__a21boi_1
X_13033_ _05719_ _05721_ _05734_ _05708_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__or4_1
X_17910_ _01502_ _01510_ _01612_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a21o_1
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18890_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\] vssd1
+ vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nor2_1
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17841_ _10195_ _10284_ _01544_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17772_ _08149_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__buf_2
X_14984_ _00008_ _07549_ _07662_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__a21oi_1
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19511_ _02905_ rbzero.wall_tracer.rayAddendY\[8\] vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__xnor2_1
X_13935_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__clkbuf_4
X_16723_ _09243_ _08821_ _08419_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__or3_1
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19442_ _02921_ _02922_ _02923_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a211oi_2
X_16654_ _09291_ _09293_ _09296_ vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__nand3_1
X_13866_ _06602_ _06557_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__xor2_4
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03042_ _03042_ vssd1 vssd1 vccd1 vccd1 clknet_0__03042_ sky130_fd_sc_hd__clkbuf_16
X_15605_ _07945_ _08238_ vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__nor2_2
XFILLER_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12817_ _05548_ _05552_ _05554_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__or3_1
XFILLER_34_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19373_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__nand2_1
X_16585_ _08329_ _08427_ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__nor2_1
X_13797_ _06529_ _06533_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__nand2_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18324_ _01902_ _02012_ _02011_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a21o_1
X_15536_ _07560_ _07562_ _08171_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__or3_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__buf_4
XFILLER_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18255_ _08257_ _01475_ _01476_ _01739_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__o22ai_1
XFILLER_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15467_ _08102_ vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__buf_2
XFILLER_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12679_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__nand2_1
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ _09783_ _09787_ _09788_ vssd1 vssd1 vccd1 vccd1 _09789_ sky130_fd_sc_hd__or3_1
X_14418_ _07146_ _07153_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__nor2_1
XFILLER_128_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18186_ _01876_ _01885_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__nand3_1
X_15398_ _08035_ _08042_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__or2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17137_ _07514_ _09763_ rbzero.row_render.size\[0\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00528_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14349_ _07084_ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__nand2_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17068_ _08519_ _09565_ vssd1 vssd1 vccd1 vccd1 _09708_ sky130_fd_sc_hd__or2_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16019_ _08622_ _08653_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__nor2_1
XFILLER_83_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20369__377 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__inv_2
XFILLER_170_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20068__105 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__inv_2
XFILLER_131_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19709_ rbzero.pov.spi_buffer\[29\] rbzero.pov.spi_buffer\[30\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20981_ clknet_leaf_49_i_clk _00750_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03309_ _03309_ vssd1 vssd1 vccd1 vccd1 clknet_0__03309_ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21602_ net143 _01371_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21533_ net454 _01302_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21464_ net385 _01233_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20415_ _02695_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_146_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21395_ net316 _01164_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ rbzero.tex_b1\[15\] _04221_ _04222_ _04218_ vssd1 vssd1 vccd1 vccd1 _04756_
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13720_ _06438_ _06455_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__o21ai_1
XFILLER_112_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10932_ rbzero.tex_b1\[25\] rbzero.tex_b1\[26\] _03806_ vssd1 vssd1 vccd1 vccd1 _03813_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19575__32 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
XFILLER_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ _05988_ _06380_ _06387_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__o21bai_1
XFILLER_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10863_ rbzero.tex_b1\[58\] rbzero.tex_b1\[59\] _03773_ vssd1 vssd1 vccd1 vccd1 _03777_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12602_ rbzero.wall_tracer.rayAddendY\[-4\] rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\]
+ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__or4_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _08361_ _07967_ _08097_ _09014_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__o31a_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _06309_ _06315_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__nor2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ rbzero.tex_g0\[28\] rbzero.tex_g0\[27\] _03740_ vssd1 vssd1 vccd1 vccd1 _03741_
+ sky130_fd_sc_hd__mux2_1
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19590__46 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__or2_1
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and2_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18040_ _08257_ _01620_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__nor2_1
X_15252_ rbzero.debug_overlay.playerX\[-7\] rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__or3_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12464_ _05217_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.trackDistY\[7\]
+ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a22o_1
Xtop_ew_algofoogle_80 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_80/HI o_rgb[10] sky130_fd_sc_hd__conb_1
X_14203_ _05825_ _06690_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__nor2_1
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_91 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_91/HI zeros[1] sky130_fd_sc_hd__conb_1
X_11415_ gpout0.hpos\[3\] _04189_ _04191_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_
+ sky130_fd_sc_hd__o211a_1
X_15183_ _07835_ _07836_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__nand2_1
X_12395_ net47 _05145_ _05143_ _05149_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a31o_1
XFILLER_126_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _06862_ _06869_ _06870_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__a21boi_1
XFILLER_153_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__buf_4
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19991_ rbzero.pov.ready_buffer\[17\] _03252_ _03253_ _04462_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01032_ sky130_fd_sc_hd__o221a_1
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ _06713_ _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__and2_1
XFILLER_140_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18942_ _02600_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11277_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _04057_ sky130_fd_sc_hd__nand2_1
X_13016_ _05747_ _05684_ _05749_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__o211a_1
XFILLER_140_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18873_ _02544_ _02545_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nand2_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17824_ _01526_ _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__xor2_1
XFILLER_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2 rbzero.spi_registers.ss_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14967_ _07653_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__clkbuf_1
X_17755_ _09249_ _10200_ _01458_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__o21ba_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ _09222_ _09236_ _09234_ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__a21o_1
X_13918_ _06617_ _06638_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__and2_1
X_12063__1 clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__inv_2
X_14898_ rbzero.wall_tracer.visualWallDist\[-8\] _07595_ vssd1 vssd1 vccd1 vccd1 _07607_
+ sky130_fd_sc_hd__or2_1
X_17686_ _10247_ _10250_ vssd1 vssd1 vccd1 vccd1 _10251_ sky130_fd_sc_hd__xor2_1
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19425_ _02893_ _02896_ _02907_ _07676_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a31o_1
X_13849_ _06574_ _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__nand2_1
X_16637_ _08237_ _09279_ _08170_ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nand2_1
XFILLER_188_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16568_ _08054_ _09029_ vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__nor2_1
XFILLER_204_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18307_ _01892_ _01893_ _01895_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__and3_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15519_ _08161_ _08163_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__nor2_1
X_19287_ _02798_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__clkbuf_1
X_16499_ _08979_ _08239_ _09141_ _09142_ vssd1 vssd1 vccd1 vccd1 _09143_ sky130_fd_sc_hd__o31a_1
XFILLER_148_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18238_ _01936_ _01937_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__xor2_1
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18169_ _01868_ _01869_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21180_ clknet_leaf_70_i_clk _00949_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20964_ clknet_leaf_68_i_clk _00733_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20895_ clknet_leaf_83_i_clk _00664_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20122__154 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__inv_2
XFILLER_179_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21516_ net437 _01285_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21447_ net368 _01216_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11200_ _03936_ _03982_ rbzero.map_rom.a6 rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1
+ _03989_ sky130_fd_sc_hd__a22o_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12180_ net9 _04950_ net11 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21378_ net299 _01147_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11131_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__inv_2
XFILLER_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11062_ rbzero.tex_b0\[28\] rbzero.tex_b0\[27\] _03876_ vssd1 vssd1 vccd1 vccd1 _03881_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15870_ rbzero.wall_tracer.visualWallDist\[-12\] _07925_ vssd1 vssd1 vccd1 vccd1
+ _08515_ sky130_fd_sc_hd__and2_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _05834_ _07392_ _07472_ _07527_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__a22o_1
XFILLER_97_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _05834_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__buf_4
X_17540_ _10103_ _10105_ vssd1 vssd1 vccd1 vccd1 _10106_ sky130_fd_sc_hd__xor2_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _04356_ vssd1 vssd1 vccd1 vccd1 _04739_
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ _06431_ _06433_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__xor2_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ rbzero.tex_b1\[33\] rbzero.tex_b1\[34\] _03795_ vssd1 vssd1 vccd1 vccd1 _03804_
+ sky130_fd_sc_hd__mux2_1
X_17471_ _10019_ _10021_ vssd1 vssd1 vccd1 vccd1 _10037_ sky130_fd_sc_hd__or2_1
X_14683_ _07107_ _07413_ _07414_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__or3_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11895_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _04272_ vssd1 vssd1 vccd1 vccd1 _04671_
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19210_ _02753_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13634_ _06351_ _06369_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__nand2_1
X_16422_ _08617_ _08672_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__xor2_2
XFILLER_189_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10846_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _03762_ vssd1 vssd1 vccd1 vccd1 _03768_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16353_ _08995_ _08997_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__xor2_2
X_19141_ _02707_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__buf_4
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13565_ _06281_ _06283_ _06301_ _06300_ _06284_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__o32a_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ rbzero.tex_g0\[36\] rbzero.tex_g0\[35\] _03729_ vssd1 vssd1 vccd1 vccd1 _03732_
+ sky130_fd_sc_hd__mux2_1
X_20097__131 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__inv_2
XFILLER_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15304_ rbzero.debug_overlay.playerX\[-4\] vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__inv_2
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19072_ _02668_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
X_12516_ _05261_ _05262_ _05266_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or4b_1
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16284_ _08870_ _08887_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__xnor2_1
X_13496_ _06229_ _06227_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__or2b_1
XFILLER_185_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18023_ _01717_ _01619_ _01723_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__and3_1
X_15235_ rbzero.wall_tracer.rayAddendX\[10\] _07855_ _07880_ _07884_ vssd1 vssd1 vccd1
+ vccd1 _00506_ sky130_fd_sc_hd__a211o_1
XFILLER_157_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12447_ _05202_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15166_ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__clkbuf_4
X_12378_ net33 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__buf_2
XFILLER_125_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _06851_ _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__and2b_1
X_11329_ _04048_ _04051_ _04053_ _04056_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a221o_1
XFILLER_140_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19974_ rbzero.pov.ready_buffer\[25\] _03247_ _03249_ rbzero.debug_overlay.facingY\[-6\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__a221o_1
X_15097_ _07678_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__buf_6
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14048_ _06666_ _06708_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__nor2_1
XFILLER_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18925_ rbzero.spi_registers.spi_counter\[4\] rbzero.spi_registers.spi_counter\[3\]
+ _02580_ rbzero.spi_registers.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a31o_1
XFILLER_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18856_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__and2_1
XFILLER_132_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17807_ _01502_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__xnor2_2
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20397__22 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18787_ rbzero.wall_tracer.trackDistY\[-2\] _02406_ _02471_ vssd1 vssd1 vccd1 vccd1
+ _00611_ sky130_fd_sc_hd__o21ba_1
X_15999_ _08642_ _08643_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17738_ _10042_ _10194_ _10192_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a21o_1
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17669_ _10103_ _10105_ vssd1 vssd1 vccd1 vccd1 _10234_ sky130_fd_sc_hd__nor2_1
XFILLER_78_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19408_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__nand2_1
XFILLER_211_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20680_ clknet_leaf_1_i_clk _00464_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19339_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nand2_1
XFILLER_176_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21301_ net222 _01070_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21232_ clknet_leaf_70_i_clk _01001_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_117_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21163_ clknet_leaf_81_i_clk _00932_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21094_ net184 _00863_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20045_ _03281_ _05190_ _03282_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__and3b_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ clknet_leaf_66_i_clk _00716_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _03646_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__buf_4
XFILLER_202_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _04436_ _04448_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nor2_4
X_20878_ clknet_leaf_61_i_clk _00647_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ rbzero.tex_g1\[40\] rbzero.tex_g1\[41\] _03647_ vssd1 vssd1 vccd1 vccd1 _03655_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13350_ _06083_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ _03618_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12301_ _04163_ _05043_ _05049_ _04809_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a22o_1
XFILLER_127_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13281_ _06010_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__nor2_1
X_10493_ _03582_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15020_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__nand2_1
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ _04996_ _04998_ _05000_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__o211a_2
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12163_ _04809_ _04907_ _04909_ net10 _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__o311a_1
XFILLER_64_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11114_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _03898_ vssd1 vssd1 vccd1 vccd1 _03908_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12094_ _04851_ _04863_ _04864_ _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a22o_1
X_16971_ _05211_ _09610_ vssd1 vssd1 vccd1 vccd1 _09611_ sky130_fd_sc_hd__nor2_2
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18710_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _02401_ _02402_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22oi_1
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ rbzero.tex_b0\[36\] rbzero.tex_b0\[35\] _03865_ vssd1 vssd1 vccd1 vccd1 _03872_
+ sky130_fd_sc_hd__mux2_1
X_15922_ _08557_ _08563_ _08565_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__nand3_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ rbzero.pov.spi_buffer\[20\] rbzero.pov.spi_buffer\[21\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
XFILLER_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03290_ _03290_ vssd1 vssd1 vccd1 vccd1 clknet_0__03290_ sky130_fd_sc_hd__clkbuf_16
X_18641_ _02237_ _02238_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__nand2_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _08074_ _08125_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__or2_1
XFILLER_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14804_ _07104_ _07450_ _05742_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__mux2_1
XFILLER_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18572_ _02039_ _02042_ _02191_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a21o_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _05721_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__inv_2
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15784_ _08426_ _08428_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__nand2_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _09967_ _09968_ vssd1 vssd1 vccd1 vccd1 _10089_ sky130_fd_sc_hd__nor2_1
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14735_ _07380_ _07427_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__nand2_1
X_11947_ _04225_ _04720_ _04721_ _04722_ _04208_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o221a_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _07400_ _07402_ _05892_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__mux2_1
XFILLER_33_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17454_ _09616_ _09729_ _10020_ vssd1 vssd1 vccd1 vccd1 _10021_ sky130_fd_sc_hd__a21oi_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11878_ _04653_ _04654_ _04265_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__mux2_1
X_13617_ _06353_ _06318_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__xnor2_1
X_16405_ _09025_ _09049_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__xnor2_2
X_10829_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _03751_ vssd1 vssd1 vccd1 vccd1 _03759_
+ sky130_fd_sc_hd__mux2_1
X_14597_ _07332_ _07333_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__nor2_1
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17385_ _09920_ _09921_ _09951_ vssd1 vssd1 vccd1 vccd1 _09952_ sky130_fd_sc_hd__a21o_1
XFILLER_186_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19124_ rbzero.spi_registers.mosi rbzero.spi_registers.mosi_buffer\[0\] _05189_ vssd1
+ vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13548_ _05945_ _05949_ _05990_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16336_ _07571_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__inv_2
XFILLER_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19055_ _02659_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
X_16267_ _08226_ _08816_ _08162_ _08160_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__or4_1
X_13479_ _05990_ _06080_ _06084_ _05991_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__o22a_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15218_ rbzero.wall_tracer.rayAddendX\[8\] rbzero.wall_tracer.rayAddendX\[7\] _07821_
+ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__o21a_1
X_18006_ _09522_ _09217_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__or3_1
XFILLER_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16198_ _08815_ _08835_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__nor2_1
XFILLER_142_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__and2_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19957_ rbzero.pov.ready _02707_ _02820_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and3_1
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20151__180 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__inv_2
XFILLER_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18908_ _02577_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19888_ _03194_ rbzero.pov.ready_buffer\[44\] _02822_ vssd1 vssd1 vccd1 vccd1 _03195_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _02516_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20801_ clknet_leaf_15_i_clk _00570_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20732_ clknet_leaf_90_i_clk _00501_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20663_ clknet_leaf_24_i_clk _00447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20594_ _02828_ _02834_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__and2b_1
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_178_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20234__255 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__inv_2
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21215_ clknet_leaf_72_i_clk _00984_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21146_ clknet_leaf_82_i_clk _00915_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21077_ net167 _00846_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20028_ _02704_ _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__nor2_1
XFILLER_150_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12850_ _04000_ _05472_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__and2_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _04224_ _04576_ _04577_ _04578_ _04141_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o221a_1
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _05512_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _07256_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__inv_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11732_ rbzero.debug_overlay.playerX\[1\] _04449_ _04464_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a22o_1
X_20391__17 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _06704_ _06761_ _07060_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__o21ba_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _04011_ _04421_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__nor2_1
XFILLER_187_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13402_ _06121_ _06125_ _06124_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__a21bo_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17170_ rbzero.traced_texa\[-1\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a22o_1
X_10614_ _03645_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__clkbuf_1
X_14382_ _07117_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__or2_1
XFILLER_168_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ _04242_ _04363_ _04372_ _04207_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o211a_1
XFILLER_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16121_ _08765_ _08758_ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__xnor2_1
X_13333_ _06057_ _06067_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nor2_1
XFILLER_128_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10545_ _03609_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _08688_ _08683_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__xnor2_1
X_13264_ _05943_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__xnor2_1
X_10476_ _03573_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15003_ rbzero.wall_tracer.stepDistX\[8\] _07579_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07672_ sky130_fd_sc_hd__mux2_1
X_12215_ _04960_ net16 net17 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a21o_1
X_13195_ _05928_ _05901_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__or2_1
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19811_ _03134_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__clkbuf_1
X_12146_ net11 _04912_ _04914_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__o211ai_1
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03311_ clknet_0__03311_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03311_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19742_ rbzero.pov.spi_buffer\[45\] rbzero.pov.spi_buffer\[46\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
X_12077_ net7 _04848_ net3 net4 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__and4b_1
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16954_ _09342_ _09328_ _09456_ vssd1 vssd1 vccd1 vccd1 _09595_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15905_ _08509_ _08544_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__xnor2_4
X_11028_ rbzero.tex_b0\[44\] rbzero.tex_b0\[43\] _03854_ vssd1 vssd1 vccd1 vccd1 _03863_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19673_ rbzero.pov.spi_buffer\[12\] rbzero.pov.spi_buffer\[13\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16885_ _08705_ vssd1 vssd1 vccd1 vccd1 _09526_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18624_ _02319_ _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__xor2_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _07958_ _08104_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__nor2_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18555_ _02184_ _02196_ _02251_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a21o_1
X_15767_ _08371_ _08411_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__xor2_1
X_12979_ _05710_ _05713_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__or3_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17506_ _10071_ _09961_ vssd1 vssd1 vccd1 vccd1 _10072_ sky130_fd_sc_hd__nand2_1
X_14718_ _07406_ _07432_ _07434_ _07454_ _05929_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__a32o_4
XFILLER_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18486_ _02182_ _02183_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__and2_1
X_15698_ _08340_ _08341_ _08342_ vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__and3_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17437_ _09709_ _09712_ vssd1 vssd1 vccd1 vccd1 _10004_ sky130_fd_sc_hd__nor2_1
XFILLER_162_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _07384_ _07385_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
XANTENNA_16 _08096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_27 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17368_ _09933_ _09934_ vssd1 vssd1 vccd1 vccd1 _09935_ sky130_fd_sc_hd__and2_1
XANTENNA_49 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19107_ rbzero.spi_registers.spi_buffer\[9\] rbzero.spi_registers.spi_buffer\[8\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16319_ _08962_ _08963_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__xnor2_1
X_17299_ rbzero.wall_tracer.trackDistX\[-5\] _09870_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09871_ sky130_fd_sc_hd__mux2_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19038_ rbzero.pov.spi_buffer\[50\] rbzero.pov.ready_buffer\[50\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21000_ clknet_leaf_52_i_clk _00769_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20715_ clknet_leaf_15_i_clk _00016_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20646_ clknet_leaf_9_i_clk _00430_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20577_ _02721_ _03448_ _03449_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__and3_1
XFILLER_137_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10330_ rbzero.tex_r1\[53\] rbzero.tex_r1\[54\] _03494_ vssd1 vssd1 vccd1 vccd1 _03495_
+ sky130_fd_sc_hd__mux2_1
XFILLER_192_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12000_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _04250_ vssd1 vssd1 vccd1 vccd1 _04775_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21129_ clknet_leaf_59_i_clk _00898_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13951_ _06675_ _06672_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__nor2_1
XFILLER_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12902_ _05562_ _05566_ _05601_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and3_1
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13882_ _06568_ _06586_ _06587_ _06618_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__a31o_1
X_16670_ _09149_ _09151_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__and2b_1
XFILLER_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__inv_2
X_15621_ _07988_ vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__inv_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _01737_ _10238_ _09294_ _09977_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__or4_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _07549_ _07552_ _07555_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__and3_1
X_12764_ _05510_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _06239_ _07071_ _07238_ _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__or4bb_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11715_ rbzero.debug_overlay.facingX\[-6\] _04475_ _04458_ rbzero.debug_overlay.facingX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__a22o_1
XFILLER_72_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15483_ _08125_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18271_ _01756_ _01970_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__xnor2_4
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__nand2_1
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17222_ _09800_ _09801_ vssd1 vssd1 vccd1 vccd1 _09802_ sky130_fd_sc_hd__xnor2_1
X_14434_ _06153_ _06705_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__and2_1
X_11646_ gpout0.hpos\[4\] _04024_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__nor2_1
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput14 i_gpout2_sel[0] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
Xinput25 i_gpout3_sel[5] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_2
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14365_ _05793_ _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__nor2_1
XFILLER_156_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17153_ rbzero.row_render.texu\[3\] _09766_ _07728_ rbzero.wall_tracer.texu\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__a22o_1
Xinput36 i_gpout5_sel[4] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_2
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ _04341_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__clkbuf_8
XFILLER_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput47 i_tex_in[1] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_16
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13316_ _05939_ _06052_ _05922_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__or3b_2
XFILLER_155_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16104_ _08745_ _08746_ _08748_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__a21boi_1
X_10528_ _03600_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17084_ _09538_ _09578_ _09723_ vssd1 vssd1 vccd1 vccd1 _09724_ sky130_fd_sc_hd__a21boi_2
X_14296_ _06703_ _06841_ _07032_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__a21oi_2
XFILLER_157_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _05945_ _05949_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__and2_2
X_16035_ _08631_ _08675_ _08678_ _08679_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__o22a_1
X_10459_ _03564_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13178_ _05880_ _05882_ _05811_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__mux2_1
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12129_ _04871_ _04881_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or3_2
XFILLER_112_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17986_ _01580_ _01590_ _01588_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a21o_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19725_ rbzero.pov.spi_buffer\[37\] rbzero.pov.spi_buffer\[38\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
X_16937_ _09575_ _09577_ vssd1 vssd1 vccd1 vccd1 _09578_ sky130_fd_sc_hd__xnor2_2
XFILLER_111_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19656_ rbzero.pov.spi_buffer\[4\] rbzero.pov.spi_buffer\[5\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16868_ _09363_ _09371_ _09508_ vssd1 vssd1 vccd1 vccd1 _09509_ sky130_fd_sc_hd__a21oi_1
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18607_ _02301_ _02302_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__and2_1
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ _08440_ _08463_ vssd1 vssd1 vccd1 vccd1 _08464_ sky130_fd_sc_hd__nand2_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20263__281 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__inv_2
XFILLER_129_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16799_ _09439_ _09440_ vssd1 vssd1 vccd1 vccd1 _09441_ sky130_fd_sc_hd__xor2_2
X_18538_ _02141_ _02160_ _02140_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a21bo_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18469_ _10094_ _09350_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__nor2_1
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20500_ _03395_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__and3_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21480_ net401 _01249_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20431_ _03338_ _03339_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__nand2_1
XFILLER_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20346__356 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__inv_2
XFILLER_84_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11500_ _04277_ _04278_ _04279_ _04226_ _04210_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__o221a_1
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12480_ _05214_ rbzero.wall_tracer.trackDistX\[10\] _05224_ rbzero.wall_tracer.trackDistY\[4\]
+ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__a221o_1
Xclkbuf_1_0__f__03314_ clknet_0__03314_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03314_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _04128_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__clkbuf_8
XFILLER_184_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20629_ clknet_leaf_76_i_clk _00413_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _06862_ _06869_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11362_ _04097_ _04114_ _04117_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__nor3_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20091__126 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__inv_2
X_13101_ _05836_ _05837_ _05807_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__mux2_1
X_10313_ rbzero.tex_r1\[61\] rbzero.tex_r1\[62\] _03483_ vssd1 vssd1 vccd1 vccd1 _03486_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1_0_i_clk clknet_1_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14081_ _06737_ _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11293_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _04073_ sky130_fd_sc_hd__nand2_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _05691_ _05673_ _05683_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__or4_1
XFILLER_191_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17840_ _10281_ _10283_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__nor2_1
XFILLER_65_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17771_ _08157_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__buf_2
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14983_ rbzero.wall_tracer.stepDistX\[-2\] _07650_ vssd1 vssd1 vccd1 vccd1 _07662_
+ sky130_fd_sc_hd__nor2_1
X_19510_ _07679_ _02978_ _02979_ _02988_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a31o_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16722_ _09244_ _09248_ vssd1 vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__nand2_1
X_13934_ _06607_ _06610_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__xor2_4
XFILLER_75_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19441_ _02904_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02924_
+ sky130_fd_sc_hd__nor2_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _08239_ _09135_ _09294_ _09295_ vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__o31ai_1
X_13865_ _06425_ _06555_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__nand2_2
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03041_ _03041_ vssd1 vssd1 vccd1 vccd1 clknet_0__03041_ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15604_ _08206_ _08248_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__xnor2_2
X_19372_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__or2_1
X_12816_ _05548_ _05552_ _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__o21ai_1
X_16584_ _09225_ _09226_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__nand2_1
X_13796_ _05855_ _05877_ _06061_ _06078_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__a41o_1
XFILLER_128_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18323_ _02016_ _02022_ rbzero.wall_tracer.trackDistX\[7\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00596_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15535_ _07989_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__clkbuf_4
XFILLER_163_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12747_ _05454_ _05456_ _05491_ _05494_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a31o_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18254_ _08257_ _08242_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__or4_1
XFILLER_147_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15466_ _08109_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__buf_4
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12678_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__nand2_1
XFILLER_129_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17205_ rbzero.wall_tracer.mapX\[8\] _05525_ vssd1 vssd1 vccd1 vccd1 _09788_ sky130_fd_sc_hd__xor2_1
X_14417_ _07146_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__and2_1
X_11629_ _04402_ _04404_ _04407_ _04306_ _04241_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a221o_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18185_ _10271_ _01766_ _01884_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__or3b_1
X_15397_ _08041_ vssd1 vssd1 vccd1 vccd1 _08042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17136_ _07855_ vssd1 vssd1 vccd1 vccd1 _09764_ sky130_fd_sc_hd__clkbuf_4
X_14348_ _07059_ _07083_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__or2_1
XFILLER_144_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14279_ _06666_ _06760_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__nor2_1
XFILLER_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17067_ _09704_ _09705_ _09706_ vssd1 vssd1 vccd1 vccd1 _09707_ sky130_fd_sc_hd__a21bo_1
XFILLER_100_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16018_ _08658_ _08662_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__xor2_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _10292_ _01671_ _01549_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__a21o_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19708_ _03047_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__clkbuf_4
X_20980_ clknet_leaf_49_i_clk _00749_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03308_ _03308_ vssd1 vssd1 vccd1 vccd1 clknet_0__03308_ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21601_ net142 _01370_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21532_ net453 _01301_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21463_ net384 _01232_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20414_ rbzero.traced_texa\[-12\] rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1 _03326_
+ sky130_fd_sc_hd__or2_1
XFILLER_135_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21394_ net315 _01163_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19639__89 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__inv_2
XFILLER_89_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ rbzero.tex_b1\[14\] _04338_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and2_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10931_ _03812_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13650_ _06381_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__and2b_1
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ _03776_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _05352_ _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and2_1
X_13581_ _06288_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nor2_1
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _03717_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__clkbuf_4
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15320_ _05196_ rbzero.wall_tracer.stepDistX\[-6\] vssd1 vssd1 vccd1 vccd1 _07965_
+ sky130_fd_sc_hd__nor2_1
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__or2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15251_ _07895_ _07595_ _07896_ _07642_ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__o211a_1
X_12463_ rbzero.wall_tracer.trackDistX\[7\] vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__inv_2
XFILLER_71_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_81 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_81/HI o_rgb[11] sky130_fd_sc_hd__conb_1
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14202_ _06926_ _06935_ _06938_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__a21boi_1
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ rbzero.row_render.size\[1\] _04192_ _04193_ _04148_ vssd1 vssd1 vccd1 vccd1
+ _04194_ sky130_fd_sc_hd__a211o_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_92 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_92/HI zeros[2] sky130_fd_sc_hd__conb_1
X_15182_ _07820_ _04462_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1
+ _07836_ sky130_fd_sc_hd__or3b_1
X_12394_ net46 _05144_ _05139_ _04323_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a22o_1
XFILLER_181_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14133_ _06863_ _06868_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__or2b_1
XFILLER_137_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11345_ _04089_ _04114_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__or3b_4
X_19990_ rbzero.pov.ready_buffer\[16\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-4\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__a221o_1
XFILLER_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ _06666_ _06663_ _06712_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__o21ai_1
X_18941_ rbzero.pov.spi_buffer\[4\] rbzero.pov.ready_buffer\[4\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
X_11276_ rbzero.texV\[8\] _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a21boi_1
XFILLER_152_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13015_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__buf_4
X_18872_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__nand2_1
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17823_ _09117_ _10266_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__nor2_1
X_20329__340 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__inv_2
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 rbzero.pov.spi_buffer\[37\] vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlygate4sd3_1
X_17754_ _09249_ _09480_ _09484_ _09096_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__o22a_1
XFILLER_94_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14966_ rbzero.wall_tracer.stepDistX\[-10\] _07484_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07653_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16705_ _09345_ _09346_ vssd1 vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__nor2_1
X_13917_ _06616_ _06595_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17685_ _09126_ _10248_ _10100_ _10249_ vssd1 vssd1 vccd1 vccd1 _10250_ sky130_fd_sc_hd__o31a_1
X_14897_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.trackDistX\[-8\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__mux2_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_32_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19424_ _02893_ _02896_ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16636_ _05209_ rbzero.wall_tracer.stepDistX\[5\] vssd1 vssd1 vccd1 vccd1 _09279_
+ sky130_fd_sc_hd__nand2_2
X_13848_ _06583_ _06584_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__nor2_1
XFILLER_165_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19355_ _02843_ _02844_ _07703_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__a21oi_1
X_16567_ _09090_ _09112_ _09110_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__a21o_1
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13779_ _05855_ _06153_ _06501_ _06502_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a22o_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18306_ _01928_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__xnor2_1
X_15518_ _08162_ _08159_ _08160_ _08151_ vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__o22a_1
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19286_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_leak\[5\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_i_clk clknet_opt_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16498_ _08977_ _08978_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__or2_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _09526_ _09703_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__nand2_1
X_20375__382 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__inv_2
X_15449_ _08093_ rbzero.debug_overlay.playerX\[-1\] _05496_ vssd1 vssd1 vccd1 vccd1
+ _08094_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20074__110 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__inv_2
XFILLER_117_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18168_ _09674_ _09693_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__nor2_1
XFILLER_191_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _09755_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__clkbuf_1
X_18099_ _01684_ _01685_ _01785_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a21o_1
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20061_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__buf_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20963_ clknet_leaf_68_i_clk _00732_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20894_ clknet_leaf_83_i_clk _00663_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21515_ net436 _01284_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21446_ net367 _01215_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21377_ net298 _01146_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__clkinv_2
XFILLER_135_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11061_ _03880_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__clkbuf_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _07547_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__clkbuf_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _07485_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__clkbuf_1
X_11963_ _04738_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13702_ _06396_ _06413_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__xor2_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10914_ _03803_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17470_ _10028_ _10035_ rbzero.wall_tracer.trackDistX\[0\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00589_ sky130_fd_sc_hd__o2bb2a_1
X_14682_ _07107_ _07413_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__nand2_2
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ _04667_ _04668_ _04669_ _04379_ _04332_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__o221a_1
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16421_ _09064_ _09065_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__or2b_1
X_13633_ _06351_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nor2_1
X_10845_ _03767_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19140_ _04890_ _04315_ _02703_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__nor4_4
XFILLER_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ _08281_ _08296_ _08996_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__a21oi_2
X_13564_ _06284_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10776_ _03731_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _07946_ _07947_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__nand2_1
XFILLER_200_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19071_ rbzero.pov.spi_buffer\[66\] rbzero.pov.ready_buffer\[66\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
X_12515_ rbzero.wall_tracer.trackDistY\[-3\] _05267_ _05263_ rbzero.wall_tracer.trackDistY\[-4\]
+ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__o221a_1
X_13495_ _06230_ _06196_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and2b_1
XFILLER_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16283_ _08924_ _08926_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__nand2_1
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18022_ _01717_ _01619_ _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15234_ _07882_ _07883_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__nor2_1
X_12446_ net71 rbzero.wall_tracer.state\[2\] _05190_ vssd1 vssd1 vccd1 vccd1 _05202_
+ sky130_fd_sc_hd__and3_1
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _05141_ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__nor2_1
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _07785_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__buf_2
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14116_ _06692_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__and2_1
XFILLER_158_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11328_ _04053_ _04056_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o21a_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ rbzero.wall_tracer.rayAddendX\[0\] _00013_ _07747_ _07755_ vssd1 vssd1 vccd1
+ vccd1 _00496_ sky130_fd_sc_hd__o22a_1
X_19973_ rbzero.pov.ready_buffer\[24\] _03247_ _03249_ rbzero.debug_overlay.facingY\[-7\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__a221o_1
XFILLER_180_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18924_ rbzero.spi_registers.spi_counter\[5\] rbzero.spi_registers.spi_counter\[4\]
+ _02583_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__and3_1
XFILLER_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14047_ _06768_ _06783_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__xnor2_1
X_11259_ rbzero.wall_tracer.state\[10\] _04038_ _04039_ vssd1 vssd1 vccd1 vccd1 _00014_
+ sky130_fd_sc_hd__o21a_1
XFILLER_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18855_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__nor2_1
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17806_ _01507_ _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__xor2_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18786_ _02464_ _02398_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__and3_1
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15998_ _07601_ _04014_ _07990_ _07936_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__and4_1
XFILLER_208_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17737_ _10186_ _10288_ _01440_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__a21o_1
X_14949_ _07621_ _07640_ _07641_ _07642_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__o211a_1
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17668_ _10197_ _10232_ vssd1 vssd1 vccd1 vccd1 _10233_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20106__139 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__inv_2
X_19407_ rbzero.wall_tracer.rayAddendY\[0\] _00013_ _02892_ vssd1 vssd1 vccd1 vccd1
+ _00810_ sky130_fd_sc_hd__o21a_1
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16619_ _09251_ _09261_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17599_ _10037_ _10038_ _10164_ vssd1 vssd1 vccd1 vccd1 _10165_ sky130_fd_sc_hd__and3_1
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19338_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nand2_1
X_19269_ _02788_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21300_ net221 _01069_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21231_ clknet_leaf_74_i_clk _01000_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_145_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21162_ clknet_leaf_81_i_clk _00931_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21093_ net183 _00862_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19617__70 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
X_20044_ _04886_ _03278_ _04887_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__a21o_1
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19632__84 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__inv_2
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_0_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ clknet_leaf_65_i_clk _00715_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ clknet_leaf_61_i_clk _00646_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ _03654_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10561_ rbzero.tex_r0\[10\] rbzero.tex_r0\[9\] _03613_ vssd1 vssd1 vccd1 vccd1 _03618_
+ sky130_fd_sc_hd__mux2_1
X_12300_ _05066_ _05067_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__or3b_2
XFILLER_195_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _06015_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__or2_1
X_10492_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _03580_ vssd1 vssd1 vccd1 vccd1 _03582_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12231_ net125 _04960_ _04966_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a2111o_2
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21429_ net350 _01198_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12162_ _04317_ _04931_ _04932_ net9 net11 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__o221a_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _03907_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ net5 net4 vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nor2_1
XFILLER_151_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16970_ rbzero.wall_tracer.visualWallDist\[11\] _04015_ vssd1 vssd1 vccd1 vccd1 _09610_
+ sky130_fd_sc_hd__nand2_1
X_20211__234 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__inv_2
XFILLER_104_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ _03871_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__clkbuf_1
X_15921_ _08557_ _08563_ _08565_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__a21o_1
XFILLER_118_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _09284_ _09287_ _08151_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a21o_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _08097_ _08491_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__nor2_1
XFILLER_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _07473_ _07499_ _07532_ _07527_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__o211a_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18571_ _02259_ _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__xor2_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _08135_ _08427_ _08422_ vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__o21ai_1
XFILLER_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _05703_ _05722_ _05727_ _05731_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a211o_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _10050_ _10087_ vssd1 vssd1 vccd1 vccd1 _10088_ sky130_fd_sc_hd__xnor2_1
X_14734_ _07378_ _07413_ _07415_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__a21o_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11946_ rbzero.tex_b0\[47\] _04347_ _04348_ _04217_ vssd1 vssd1 vccd1 vccd1 _04722_
+ sky130_fd_sc_hd__a31o_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _09726_ _09728_ vssd1 vssd1 vccd1 vccd1 _10020_ sky130_fd_sc_hd__nor2_1
X_14665_ _07386_ _07401_ _05779_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__mux2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ rbzero.tex_g1\[25\] rbzero.tex_g1\[24\] _04336_ vssd1 vssd1 vccd1 vccd1 _04654_
+ sky130_fd_sc_hd__mux2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16404_ _09047_ _09048_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__xnor2_2
X_13616_ _06319_ _06316_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__or2b_1
X_10828_ _03758_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
X_17384_ _09938_ _09950_ vssd1 vssd1 vccd1 vccd1 _09951_ sky130_fd_sc_hd__xnor2_1
X_14596_ _07216_ _07331_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nor2_1
XFILLER_164_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19123_ _02696_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__clkbuf_1
X_16335_ _08230_ rbzero.wall_tracer.stepDistY\[6\] vssd1 vssd1 vccd1 vccd1 _08980_
+ sky130_fd_sc_hd__nand2_1
X_13547_ _06136_ _06137_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__xor2_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10759_ _03722_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19054_ rbzero.pov.spi_buffer\[58\] rbzero.pov.ready_buffer\[58\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16266_ _08853_ _08910_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13478_ _05990_ _06134_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__nor2_1
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18005_ _01582_ _01706_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__xnor2_1
X_15217_ _07845_ _07864_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__nor2_1
X_12429_ _05191_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__clkbuf_1
X_16197_ _08840_ _08841_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__nor2_1
XFILLER_126_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15148_ _07802_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__nor2_1
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15079_ rbzero.wall_tracer.rayAddendX\[-1\] _07706_ _07739_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _07740_ sky130_fd_sc_hd__a22o_1
X_19956_ rbzero.pov.ready_buffer\[36\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-6\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__o221a_1
XFILLER_136_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18907_ _02574_ _02575_ _02576_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__and3_1
XFILLER_68_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20186__211 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__inv_2
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19887_ rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__inv_2
XFILLER_132_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18838_ rbzero.wall_tracer.trackDistY\[5\] _02515_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_110_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18769_ rbzero.wall_tracer.trackDistY\[-4\] _02455_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20800_ clknet_leaf_15_i_clk _00569_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20731_ clknet_leaf_85_i_clk _00500_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20662_ clknet_leaf_24_i_clk _00446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20593_ _07679_ _02832_ _03459_ _07855_ rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__a32o_1
XFILLER_143_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21214_ clknet_leaf_72_i_clk _00983_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21145_ clknet_leaf_61_i_clk _00914_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21076_ net166 _00845_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20027_ _04892_ _04992_ _04883_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ rbzero.tex_g0\[47\] _04135_ _04136_ _04126_ vssd1 vssd1 vccd1 vccd1 _04578_
+ sky130_fd_sc_hd__a31o_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _05524_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ rbzero.debug_overlay.playerX\[-7\] _04455_ _04458_ rbzero.debug_overlay.playerX\[-9\]
+ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a221o_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ clknet_leaf_13_i_clk _00698_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _06153_ _07072_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21o_1
XFILLER_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11662_ gpout0.hpos\[7\] _04414_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__nor2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13401_ _06136_ _06137_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__or2b_1
XFILLER_211_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ rbzero.tex_g1\[48\] rbzero.tex_g1\[49\] _03635_ vssd1 vssd1 vccd1 vccd1 _03645_
+ sky130_fd_sc_hd__mux2_1
XFILLER_211_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14381_ _06696_ _06760_ _07116_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__o21ba_1
X_11593_ _04254_ _04366_ _04370_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__a211o_1
XFILLER_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _08759_ _08756_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__and2b_1
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13332_ _06058_ _06063_ _06064_ _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a2bb2o_1
X_10544_ rbzero.tex_r0\[18\] rbzero.tex_r0\[17\] _03602_ vssd1 vssd1 vccd1 vccd1 _03609_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16051_ _08638_ _08651_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10475_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _03569_ vssd1 vssd1 vccd1 vccd1 _03573_
+ sky130_fd_sc_hd__mux2_1
X_13263_ _05998_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__nor2_1
XFILLER_108_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ _07671_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12214_ net18 net19 _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__and3b_1
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13194_ _05826_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12145_ _04910_ net66 _04915_ net12 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a211o_1
X_19810_ rbzero.pov.sclk_buffer\[1\] rbzero.pov.sclk_buffer\[0\] _05189_ vssd1 vssd1
+ vccd1 vccd1 _03134_ sky130_fd_sc_hd__mux2_1
XFILLER_97_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03310_ clknet_0__03310_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03310_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ _04840_ net64 _04846_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a211o_1
X_16953_ _09592_ _09593_ vssd1 vssd1 vccd1 vccd1 _09594_ sky130_fd_sc_hd__nor2_4
X_19741_ _03098_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15904_ _08547_ _08548_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__nor2_4
X_11027_ _03862_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__clkbuf_1
X_19672_ _03062_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__clkbuf_1
X_16884_ _08705_ _08059_ _09524_ vssd1 vssd1 vccd1 vccd1 _09525_ sky130_fd_sc_hd__or3_1
XFILLER_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20406__7 clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
X_18623_ _02229_ _02231_ _02230_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a21boi_1
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _07913_ _07967_ _08022_ _07923_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__o22ai_1
XFILLER_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19611__65 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
XFILLER_46_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18554_ _02193_ _02195_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__nor2_1
X_15766_ _08400_ _08409_ _08410_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__a21oi_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _05584_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__xor2_2
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17505_ _09663_ _09959_ vssd1 vssd1 vccd1 vccd1 _10071_ sky130_fd_sc_hd__or2_1
XFILLER_75_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _07439_ _07444_ _07449_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__nand4_1
X_11929_ rbzero.tex_b0\[56\] _04338_ _04225_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a21o_1
X_18485_ _02171_ _02181_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or2_1
X_15697_ _08097_ _08022_ vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__nor2_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ _09994_ _10002_ vssd1 vssd1 vccd1 vccd1 _10003_ sky130_fd_sc_hd__xnor2_1
X_14648_ _05893_ _07365_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__and2_1
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _08158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_39 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _09931_ _09932_ vssd1 vssd1 vccd1 vccd1 _09934_ sky130_fd_sc_hd__nand2_1
XFILLER_174_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14579_ _07285_ _07293_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__nand2_1
X_19106_ _02686_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16318_ _07913_ _08264_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__and2b_1
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17298_ _09863_ _09867_ _09868_ _09869_ vssd1 vssd1 vccd1 vccd1 _09870_ sky130_fd_sc_hd__o31ai_1
XFILLER_174_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19037_ _02650_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__clkbuf_1
X_16249_ _08877_ _08878_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__or2b_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19939_ _02820_ _03232_ _03197_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__o21a_1
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20240__260 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__inv_2
X_20714_ clknet_leaf_11_i_clk _00005_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20645_ clknet_leaf_8_i_clk _00429_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__or2_1
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20158__187 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__inv_2
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21128_ clknet_leaf_59_i_clk _00897_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _06685_ _06686_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__nand2_1
X_21059_ clknet_leaf_56_i_clk _00828_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12901_ _05632_ _05634_ _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__or4b_4
XFILLER_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13881_ _06591_ _06589_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__and2b_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _08263_ _08264_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__and2_1
X_20323__335 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__inv_2
X_12832_ _04031_ _05372_ _05568_ _04001_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a211o_1
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _07894_ _05459_ _08195_ _05193_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__a211o_1
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12763_ rbzero.map_rom.f2 _05509_ _05414_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__mux2_1
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14502_ _06002_ _06770_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__nand2_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _01969_ _10110_ _01879_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ rbzero.debug_overlay.facingX\[-3\] _04463_ _04466_ rbzero.debug_overlay.facingX\[-8\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__a221o_1
XFILLER_202_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15482_ _08126_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__inv_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _05418_ _05439_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__nand3b_1
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ rbzero.wall_tracer.mapX\[11\] _05525_ vssd1 vssd1 vccd1 vccd1 _09801_ sky130_fd_sc_hd__xnor2_1
X_14433_ _07142_ _07169_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__or2_1
XFILLER_202_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11645_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__inv_2
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17152_ rbzero.row_render.texu\[2\] _09766_ _07728_ rbzero.wall_tracer.texu\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__a22o_1
X_14364_ _07099_ _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__or2_2
Xinput15 i_gpout2_sel[1] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11576_ _04232_ _04333_ _04340_ _04354_ _04244_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o311a_1
Xinput26 i_gpout4_sel[0] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_4
Xinput37 i_gpout5_sel[5] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
Xinput48 i_tex_in[2] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
X_16103_ _07964_ _08674_ _08747_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__or3_1
X_13315_ _05973_ _05961_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__or2_1
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10527_ rbzero.tex_r0\[26\] rbzero.tex_r0\[25\] _03591_ vssd1 vssd1 vccd1 vccd1 _03600_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17083_ _09575_ _09577_ vssd1 vssd1 vccd1 vccd1 _09723_ sky130_fd_sc_hd__or2b_1
X_14295_ _06818_ _06840_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__nor2_1
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ _08008_ _08104_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__or2_1
X_10458_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _03558_ vssd1 vssd1 vccd1 vccd1 _03564_
+ sky130_fd_sc_hd__mux2_1
X_13246_ _05961_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__buf_2
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _03525_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
X_13177_ _05902_ _05879_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__or2_1
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ net7 _04882_ _04894_ _04899_ _04837_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a32o_2
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17985_ _01575_ _01607_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__or2_1
XFILLER_97_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12059_ _03474_ _04815_ _04005_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__o21ai_1
X_19724_ _03089_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
X_16936_ _09415_ _09441_ _09576_ vssd1 vssd1 vccd1 vccd1 _09577_ sky130_fd_sc_hd__a21o_1
XFILLER_133_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19655_ _03053_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__clkbuf_1
X_16867_ _09244_ _09248_ _09370_ vssd1 vssd1 vccd1 vccd1 _09508_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15818_ _08460_ _08461_ _08462_ vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__a21oi_1
X_18606_ _02301_ _02302_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__nor2_1
XFILLER_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16798_ _09297_ _09299_ vssd1 vssd1 vccd1 vccd1 _09440_ sky130_fd_sc_hd__and2_1
X_20298__312 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__inv_2
X_18537_ _02228_ _02234_ rbzero.wall_tracer.trackDistX\[9\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00598_ sky130_fd_sc_hd__o2bb2a_1
X_15749_ _08316_ _08314_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__nand2_1
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18468_ _02038_ _02053_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a21bo_1
XFILLER_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17419_ _09975_ _09985_ vssd1 vssd1 vccd1 vccd1 _09986_ sky130_fd_sc_hd__xor2_2
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18399_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__and2b_1
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20430_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03339_
+ sky130_fd_sc_hd__nand2_1
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20164__191 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__inv_2
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03313_ clknet_0__03313_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03313_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11430_ _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__buf_4
X_20628_ clknet_leaf_18_i_clk _00412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11361_ _04093_ _04114_ _04122_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__nor3_4
XFILLER_138_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20559_ _09763_ _09194_ rbzero.traced_texVinit\[3\] _09762_ vssd1 vssd1 vccd1 vccd1
+ _01411_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13100_ _05642_ _05645_ _05796_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__mux2_1
X_10312_ _03485_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14080_ _06798_ _06816_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _04072_ sky130_fd_sc_hd__or2_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13031_ _05642_ _05744_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nand2_1
XFILLER_191_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17770_ _05198_ _08445_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__nand2_2
X_14982_ _07661_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16721_ _09226_ _09228_ _09225_ vssd1 vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__a21bo_1
X_13933_ _06666_ _06668_ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__or3_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19440_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__and2_1
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ _09133_ _09134_ vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__or2_1
X_13864_ _06559_ _06378_ _06558_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__nand3_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03040_ _03040_ vssd1 vssd1 vccd1 vccd1 clknet_0__03040_ sky130_fd_sc_hd__clkbuf_16
X_15603_ _08241_ _08247_ vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__xor2_2
X_19371_ _02859_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__clkbuf_1
X_12815_ rbzero.wall_tracer.mapY\[10\] _05404_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__xor2_1
XFILLER_90_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16583_ _08823_ _08159_ _08151_ _09096_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__o22ai_1
X_13795_ _06057_ _06530_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__o21ba_1
XFILLER_15_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18322_ _02020_ _02021_ _09817_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__o21a_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15534_ _08170_ _08178_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__nor2_1
X_12746_ _05492_ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__or2_1
XFILLER_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _01859_ _01863_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__nand2_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15465_ _08109_ _08085_ _08104_ vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__or3_1
XFILLER_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__nor2_1
XFILLER_163_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17204_ rbzero.wall_tracer.mapX\[7\] _05512_ _09782_ vssd1 vssd1 vccd1 vccd1 _09787_
+ sky130_fd_sc_hd__o21a_1
X_14416_ _07147_ _07152_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11628_ _04405_ _04406_ _04218_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
X_18184_ _10271_ _01766_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__o21bai_1
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15396_ _08039_ _08040_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__nand2_1
XFILLER_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17135_ _07831_ vssd1 vssd1 vccd1 vccd1 _09763_ sky130_fd_sc_hd__buf_2
X_14347_ _07059_ _07083_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__nand2_1
X_11559_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__buf_4
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17066_ _03953_ _09283_ _08377_ _09433_ vssd1 vssd1 vccd1 vccd1 _09706_ sky130_fd_sc_hd__or4_1
X_14278_ _07013_ _07014_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__xor2_2
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16017_ _08659_ _08661_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__nand2_2
XFILLER_171_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13229_ _05648_ _05792_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__nor2_1
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _01441_ _01547_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__or2_1
XFILLER_78_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19707_ _03080_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16919_ _07602_ _09283_ _05209_ _09287_ vssd1 vssd1 vccd1 vccd1 _09560_ sky130_fd_sc_hd__or4_1
XFILLER_168_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17899_ _01592_ _01601_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__03307_ _03307_ vssd1 vssd1 vccd1 vccd1 clknet_0__03307_ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19638_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__buf_1
XFILLER_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19569_ rbzero.pov.spi_counter\[6\] _03034_ _03036_ vssd1 vssd1 vccd1 vccd1 _00828_
+ sky130_fd_sc_hd__o21a_1
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21600_ net141 _01369_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21531_ net452 _01300_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21462_ net383 _01231_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20413_ rbzero.traced_texa\[-12\] rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1 _03325_
+ sky130_fd_sc_hd__nand2_1
XFILLER_175_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21393_ net314 _01162_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20352__361 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__inv_2
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10930_ rbzero.tex_b1\[26\] rbzero.tex_b1\[27\] _03806_ vssd1 vssd1 vccd1 vccd1 _03812_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ rbzero.tex_b1\[59\] rbzero.tex_b1\[60\] _03773_ vssd1 vssd1 vccd1 vccd1 _03776_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12600_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__or2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13580_ _06287_ _06286_ _05988_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__o21a_1
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _03739_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12531_ _05285_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _07595_ _07592_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__nand2_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ rbzero.wall_tracer.trackDistX\[8\] vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__inv_2
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14201_ _06805_ _06678_ _06937_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__or3b_1
XFILLER_138_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ rbzero.row_render.size\[2\] gpout0.hpos\[2\] _04163_ gpout0.hpos\[0\] vssd1
+ vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__a22o_1
Xtop_ew_algofoogle_82 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_82/HI o_rgb[12] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_93 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_93/HI zeros[3] sky130_fd_sc_hd__conb_1
X_15181_ _07820_ _04462_ _07833_ _07834_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__o22ai_1
X_12393_ _05145_ _05143_ _04021_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a31o_1
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14132_ _06863_ _06868_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11344_ _04082_ _04088_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nand2_1
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _06786_ _06794_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__xor2_1
XFILLER_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18940_ _02599_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__clkbuf_1
X_11275_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _04055_ sky130_fd_sc_hd__nand2_1
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13014_ _05750_ _05702_ _05683_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__or3_1
X_18871_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__or2_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17822_ _01524_ _01525_ _10131_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__or3b_1
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 rbzero.spi_registers.mosi vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14965_ _07652_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__clkbuf_1
X_17753_ _10235_ _10253_ _01456_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a21o_1
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13916_ _06644_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20180__206 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__inv_2
X_16704_ _09220_ _09344_ vssd1 vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__and2_1
X_17684_ _09670_ _10099_ vssd1 vssd1 vccd1 vccd1 _10249_ sky130_fd_sc_hd__nand2_1
X_14896_ _07591_ _07604_ _07605_ _04039_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__o211a_1
XFILLER_78_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19423_ _02906_ rbzero.wall_tracer.rayAddendY\[2\] vssd1 vssd1 vccd1 vccd1 _02907_
+ sky130_fd_sc_hd__xnor2_1
X_16635_ _08242_ _09129_ _08180_ vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__a21oi_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _06263_ _06582_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__and2_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19354_ _02840_ _02841_ _02842_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__o21ai_1
X_16566_ _09175_ _09176_ _09178_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__o21ai_1
X_13778_ _06513_ _06514_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__and2b_1
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18305_ _02003_ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__and2b_1
X_15517_ _08135_ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__clkbuf_4
XFILLER_176_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12729_ _05424_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__and2_2
X_19285_ _02797_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__clkbuf_1
X_16497_ _08985_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18236_ _01933_ _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__nand2_1
XFILLER_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15448_ _08028_ _08092_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__and2_1
XFILLER_176_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18167_ _01866_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__xnor2_2
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15379_ _07913_ _07924_ _07941_ _07967_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__or4_1
XFILLER_128_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _09753_ _04319_ _09754_ vssd1 vssd1 vccd1 vccd1 _09755_ sky130_fd_sc_hd__and3_1
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18098_ _01670_ _01673_ _01789_ _01669_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a211o_1
XFILLER_144_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17049_ _09683_ _09688_ vssd1 vssd1 vccd1 vccd1 _09689_ sky130_fd_sc_hd__and2_1
XFILLER_104_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ clknet_leaf_68_i_clk _00731_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ clknet_leaf_83_i_clk _00662_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21514_ net435 _01283_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20276__292 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__inv_2
XFILLER_148_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21445_ net366 _01214_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21376_ net297 _01145_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20327_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__buf_1
XFILLER_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _03876_ vssd1 vssd1 vccd1 vccd1 _03880_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ rbzero.wall_tracer.stepDistY\[-10\] _07484_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07485_ sky130_fd_sc_hd__mux2_1
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _04735_ _04737_ _04324_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__o21bai_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _06436_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__nand2_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ rbzero.tex_b1\[34\] rbzero.tex_b1\[35\] _03795_ vssd1 vssd1 vccd1 vccd1 _03803_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14681_ _07106_ _07415_ _07416_ _07417_ _05892_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__o311a_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _04272_ vssd1 vssd1 vccd1 vccd1 _04669_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16420_ _09061_ _09062_ _09063_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__a21o_1
X_13632_ _06352_ _06367_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__a21o_1
X_10844_ rbzero.tex_g0\[4\] rbzero.tex_g0\[3\] _03762_ vssd1 vssd1 vccd1 vccd1 _03767_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16351_ _08249_ _08280_ vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__nor2_1
X_13563_ _06291_ _06298_ _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__o21a_1
XFILLER_125_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10775_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _03729_ vssd1 vssd1 vccd1 vccd1 _03731_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15302_ rbzero.debug_overlay.playerX\[-5\] _07898_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__o21ai_1
XFILLER_201_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ rbzero.wall_tracer.trackDistY\[3\] _05264_ rbzero.wall_tracer.trackDistY\[2\]
+ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__o22a_1
X_19070_ _02667_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16282_ _08924_ _08926_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__nor2_1
X_13494_ _06196_ _06230_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18021_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__inv_2
X_15233_ _07870_ _07873_ _07881_ _07830_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__a31o_1
XFILLER_201_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ _05201_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15164_ _07788_ _07797_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__nand2_1
X_12376_ net32 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__clkbuf_4
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14115_ _06675_ _06690_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__nor2_1
XFILLER_158_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ _04101_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15095_ _07703_ _07753_ _07754_ _07706_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__a31o_1
X_19972_ rbzero.pov.ready_buffer\[23\] _03240_ _03243_ rbzero.debug_overlay.facingY\[-8\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__o221a_1
XFILLER_125_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14046_ _06781_ _06782_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__or2b_1
XFILLER_141_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18923_ _02588_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11258_ _04035_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18854_ _02529_ _02016_ rbzero.wall_tracer.trackDistY\[7\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00620_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11189_ _03977_ _03936_ _03919_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__and3b_1
XFILLER_68_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17805_ _09276_ _09674_ _10245_ _01508_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__o31a_1
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18785_ _02468_ _05531_ _02469_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__or3b_1
X_15997_ _07598_ _07951_ _05207_ _07927_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__or4b_1
XFILLER_76_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14948_ _04035_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__buf_4
X_17736_ _10285_ _10287_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__nor2_1
XFILLER_208_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17667_ _10199_ _10231_ vssd1 vssd1 vccd1 vccd1 _10232_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14879_ _05278_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__buf_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19406_ _04035_ _02882_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a21o_1
XFILLER_78_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ _09259_ _09260_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__nor2_1
XFILLER_211_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17598_ _10039_ _10163_ vssd1 vssd1 vccd1 vccd1 _10164_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16549_ _09089_ _09192_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__xnor2_2
X_19337_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__nor2_1
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19268_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_floor\[4\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_163_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18219_ _01854_ _01819_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__or2b_1
XFILLER_176_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19199_ rbzero.spi_registers.new_sky\[3\] rbzero.color_sky\[3\] _02740_ vssd1 vssd1
+ vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_102_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21230_ clknet_leaf_70_i_clk _00999_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21161_ clknet_leaf_84_i_clk _00930_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21092_ net182 _00861_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20043_ _04887_ _04886_ _03278_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__and3_1
XFILLER_113_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ clknet_leaf_65_i_clk _00714_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20876_ clknet_leaf_61_i_clk _00645_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _03617_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10491_ _03581_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12230_ gpout2.clk_div\[1\] _04981_ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21428_ net349 _01197_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12161_ gpout0.hpos\[0\] _04163_ _04910_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21359_ net280 _01128_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11112_ rbzero.tex_b0\[4\] rbzero.tex_b0\[3\] _03898_ vssd1 vssd1 vccd1 vccd1 _03907_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12092_ _04021_ _04855_ _04853_ net42 vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a22o_1
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _03865_ vssd1 vssd1 vccd1 vccd1 _03871_
+ sky130_fd_sc_hd__mux2_1
X_15920_ _08564_ _08503_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__xor2_1
XFILLER_110_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_i_clk clknet_opt_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _08495_ _08141_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__xnor2_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _07473_ _07492_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__nand2_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18570_ _02265_ _02266_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__xnor2_1
X_15782_ _08425_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__buf_4
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _05702_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__nor3_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__clkbuf_4
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17521_ _10085_ _10086_ vssd1 vssd1 vccd1 vccd1 _10087_ sky130_fd_sc_hd__nand2_1
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ rbzero.tex_b0\[46\] _04337_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__and2_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17452_ _09918_ _10018_ vssd1 vssd1 vccd1 vccd1 _10019_ sky130_fd_sc_hd__xnor2_4
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _05893_ _07041_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__and2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ rbzero.tex_g1\[27\] rbzero.tex_g1\[26\] _04271_ vssd1 vssd1 vccd1 vccd1 _04653_
+ sky130_fd_sc_hd__mux2_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16403_ _08165_ _08432_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__and2_1
X_13615_ _06338_ _06343_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10827_ rbzero.tex_g0\[12\] rbzero.tex_g0\[11\] _03751_ vssd1 vssd1 vccd1 vccd1 _03758_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17383_ _09947_ _09949_ vssd1 vssd1 vccd1 vccd1 _09950_ sky130_fd_sc_hd__xor2_1
X_14595_ _07216_ _07331_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__and2_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19122_ net42 rbzero.spi_registers.mosi_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02696_ sky130_fd_sc_hd__mux2_1
X_16334_ _08977_ _08978_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__xnor2_2
XFILLER_201_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13546_ _05824_ _06080_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__or3_2
X_20292__307 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__inv_2
XFILLER_119_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10758_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _03718_ vssd1 vssd1 vccd1 vccd1 _03722_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19053_ _02658_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
X_16265_ _08901_ _08908_ _08909_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__a21oi_1
X_13477_ _06041_ _06067_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__or2_1
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10689_ _03685_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ _07863_ _07867_ _00013_ rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1
+ vccd1 _00504_ sky130_fd_sc_hd__o2bb2a_1
X_18004_ _08445_ _09353_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__nand2_1
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12428_ net71 rbzero.wall_tracer.state\[12\] _05190_ vssd1 vssd1 vccd1 vccd1 _05191_
+ sky130_fd_sc_hd__and3_1
XFILLER_161_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16196_ _08831_ _08837_ _08839_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__and3_1
XFILLER_126_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _07730_ rbzero.debug_overlay.vplaneX\[-5\] _07800_ _07801_ vssd1 vssd1 vccd1
+ vccd1 _07803_ sky130_fd_sc_hd__nor4_1
X_12359_ gpout4.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__inv_2
XFILLER_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ rbzero.debug_overlay.vplaneX\[-6\] _07735_ _07738_ vssd1 vssd1 vccd1 vccd1
+ _07739_ sky130_fd_sc_hd__o21ai_1
X_19955_ _02721_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14029_ _06762_ _06764_ _06765_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__nand3_1
X_18906_ rbzero.spi_registers.spi_counter\[0\] _02558_ vssd1 vssd1 vccd1 vccd1 _02576_
+ sky130_fd_sc_hd__nand2_1
XFILLER_136_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19886_ _03192_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18837_ _02513_ _02514_ _01792_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18768_ _09812_ _02454_ _09877_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o21ai_1
X_17719_ _10281_ _10283_ vssd1 vssd1 vccd1 vccd1 _10284_ sky130_fd_sc_hd__xor2_1
XFILLER_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18699_ _02390_ _02394_ rbzero.wall_tracer.trackDistX\[11\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00600_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_208_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20730_ clknet_leaf_86_i_clk _00499_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20661_ clknet_leaf_9_i_clk _00445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20592_ _02829_ _02831_ _02830_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__a21bo_1
XFILLER_176_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21213_ clknet_leaf_72_i_clk _00982_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21144_ clknet_leaf_61_i_clk _00913_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21075_ net165 _00844_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20026_ _03259_ _03268_ _03269_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__a21oi_1
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ rbzero.debug_overlay.playerX\[-6\] _04475_ _04454_ rbzero.debug_overlay.playerX\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a22o_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ clknet_leaf_76_i_clk _00697_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _04418_ _04430_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__and2_1
XFILLER_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20859_ clknet_leaf_55_i_clk _00628_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ _06068_ _06064_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__xor2_1
XFILLER_168_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ _03644_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__clkbuf_1
X_14380_ _06176_ _07116_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__and2_1
XFILLER_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11592_ _04119_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__buf_4
XFILLER_161_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _06065_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__nor2_1
XFILLER_195_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10543_ _03608_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16050_ _08692_ _08694_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__nor2_1
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13262_ _05977_ _05987_ _05997_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and3_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _03572_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15001_ rbzero.wall_tracer.stepDistX\[7\] _07575_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07671_ sky130_fd_sc_hd__mux2_1
X_12213_ _04977_ net16 _04979_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a31o_1
XFILLER_109_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _05901_ _05891_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20135__166 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__inv_2
XFILLER_159_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12144_ _04910_ _04325_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__nor2_1
XFILLER_151_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19740_ rbzero.pov.spi_buffer\[44\] rbzero.pov.spi_buffer\[45\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03098_ sky130_fd_sc_hd__mux2_1
X_12075_ _04840_ _04738_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__nor2_1
XFILLER_150_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16952_ _09454_ _09591_ vssd1 vssd1 vccd1 vccd1 _09593_ sky130_fd_sc_hd__nor2_1
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15903_ _08470_ _08546_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__and2_1
X_11026_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _03854_ vssd1 vssd1 vccd1 vccd1 _03862_
+ sky130_fd_sc_hd__mux2_1
X_19671_ rbzero.pov.spi_buffer\[11\] rbzero.pov.spi_buffer\[12\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XFILLER_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16883_ _09521_ _09523_ vssd1 vssd1 vccd1 vccd1 _09524_ sky130_fd_sc_hd__nand2_1
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18622_ _02317_ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__nand2_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _08477_ _08472_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__xor2_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _02235_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__xnor2_1
X_15765_ _08372_ _08399_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__nor2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _05567_ _05599_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
XFILLER_46_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _09391_ _08427_ _09941_ _09942_ vssd1 vssd1 vccd1 vccd1 _10070_ sky130_fd_sc_hd__o31ai_2
X_11928_ rbzero.tex_b0\[57\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__and3_1
X_14716_ _07104_ _07450_ _07451_ _07452_ _05742_ _07375_ vssd1 vssd1 vccd1 vccd1 _07453_
+ sky130_fd_sc_hd__mux4_2
X_15696_ _08338_ _08339_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__nand2_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18484_ _02171_ _02181_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__nand2_1
XFILLER_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20300__314 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__inv_2
XFILLER_127_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14647_ _05893_ _07101_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__nor2_1
X_17435_ _10000_ _10001_ vssd1 vssd1 vccd1 vccd1 _10002_ sky130_fd_sc_hd__xnor2_2
XFILLER_166_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11859_ _04379_ _04633_ _04634_ _04635_ _04229_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__o221a_1
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_18 _08215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _07311_ _07313_ _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__a21o_1
XFILLER_159_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17366_ _09931_ _09932_ vssd1 vssd1 vccd1 vccd1 _09933_ sky130_fd_sc_hd__or2_1
XFILLER_186_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19105_ rbzero.spi_registers.spi_buffer\[8\] rbzero.spi_registers.spi_buffer\[7\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
X_13529_ _06255_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16317_ _07924_ _08276_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__nor2_1
X_17297_ _09807_ _09194_ vssd1 vssd1 vccd1 vccd1 _09869_ sky130_fd_sc_hd__or2_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19036_ rbzero.pov.spi_buffer\[49\] rbzero.pov.ready_buffer\[49\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
X_16248_ _08872_ _08128_ _08868_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__or3_1
XFILLER_51_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ _08519_ _08823_ _08329_ _08377_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__o22ai_1
XFILLER_86_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19938_ _03920_ _03227_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__and2_1
X_19869_ rbzero.debug_overlay.playerX\[2\] _03155_ _03179_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00985_ sky130_fd_sc_hd__o211a_1
XFILLER_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20713_ clknet_leaf_9_i_clk _00004_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20644_ clknet_leaf_7_i_clk _00428_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20575_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__nand2_1
XFILLER_192_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21127_ clknet_leaf_66_i_clk _00896_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21058_ clknet_leaf_56_i_clk _00827_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _05628_ _05626_ _05633_ _05631_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a211o_1
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20009_ _03256_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
X_13880_ _06592_ _06567_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and2b_1
XFILLER_207_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ rbzero.wall_tracer.visualWallDist\[8\] _04031_ vssd1 vssd1 vccd1 vccd1 _05568_
+ sky130_fd_sc_hd__nor2_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _07893_ _05369_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__nor2_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ rbzero.debug_overlay.playerX\[2\] _05508_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05509_ sky130_fd_sc_hd__mux2_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _06002_ _07072_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__nand2_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ rbzero.debug_overlay.facingX\[0\] _04459_ _04460_ rbzero.debug_overlay.facingX\[-2\]
+ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a221o_1
XFILLER_199_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15481_ _08034_ _08046_ _08124_ _08125_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__or4_1
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _05436_ _05440_ _05434_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__o21a_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _07141_ _07140_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__and2b_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ rbzero.wall_tracer.mapX\[10\] _05525_ _09799_ vssd1 vssd1 vccd1 vccd1 _09800_
+ sky130_fd_sc_hd__a21bo_1
X_11644_ _04415_ _04417_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__and2b_1
XFILLER_202_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17151_ rbzero.row_render.texu\[1\] _09766_ _07728_ rbzero.wall_tracer.texu\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__a22o_1
X_14363_ _07043_ _07098_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__nor2_1
X_11575_ _04306_ _04346_ _04353_ _04241_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a211o_1
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 i_gpout2_sel[2] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_16
XFILLER_155_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 i_gpout4_sel[1] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_6
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16102_ _07601_ _08227_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__nand2_2
X_13314_ _06021_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 i_mode[0] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_8
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10526_ _03599_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
Xinput49 i_tex_in[3] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_6
X_17082_ _09680_ _09721_ vssd1 vssd1 vccd1 vccd1 _09722_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14294_ _06735_ _07030_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__xnor2_2
XFILLER_156_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ _08676_ _08677_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__and2_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13245_ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__clkbuf_4
X_10457_ _03563_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _05778_ _05829_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a21o_1
XFILLER_124_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10388_ rbzero.tex_r1\[25\] rbzero.tex_r1\[26\] _03516_ vssd1 vssd1 vccd1 vccd1 _03525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _04851_ _04896_ _04898_ _04865_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a22o_2
X_17984_ _01445_ _01447_ _01571_ _01569_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a31o_1
XFILLER_96_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19723_ rbzero.pov.spi_buffer\[36\] rbzero.pov.spi_buffer\[37\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
X_12058_ _04812_ _04817_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__or3b_1
XFILLER_133_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16935_ _09439_ _09440_ vssd1 vssd1 vccd1 vccd1 _09576_ sky130_fd_sc_hd__nor2_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11009_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _03843_ vssd1 vssd1 vccd1 vccd1 _03853_
+ sky130_fd_sc_hd__mux2_1
X_19654_ rbzero.pov.spi_buffer\[3\] rbzero.pov.spi_buffer\[4\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03053_ sky130_fd_sc_hd__mux2_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16866_ _09499_ _09506_ vssd1 vssd1 vccd1 vccd1 _09507_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18605_ _02204_ _02214_ _02202_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15817_ _08441_ _08459_ vssd1 vssd1 vccd1 vccd1 _08462_ sky130_fd_sc_hd__nor2_1
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16797_ _09425_ _09438_ vssd1 vssd1 vccd1 vccd1 _09439_ sky130_fd_sc_hd__xnor2_2
XFILLER_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18536_ _02232_ _02233_ _09817_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__o21a_1
XFILLER_206_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _07996_ _08194_ _08386_ _08385_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__o31a_1
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _02054_ _02035_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__or2b_1
X_15679_ _08317_ _08323_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17418_ _09979_ _09984_ vssd1 vssd1 vccd1 vccd1 _09985_ sky130_fd_sc_hd__xor2_2
XFILLER_166_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18398_ _02093_ _02095_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__nand2_1
XFILLER_140_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17349_ _09654_ _09909_ _09914_ vssd1 vssd1 vccd1 vccd1 _09916_ sky130_fd_sc_hd__and3_1
XFILLER_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20360_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__buf_1
XFILLER_101_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ rbzero.pov.spi_buffer\[41\] rbzero.pov.ready_buffer\[41\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
X_20118__150 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__inv_2
XFILLER_115_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19587__43 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_83_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03312_ clknet_0__03312_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03312_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20627_ clknet_leaf_51_i_clk _00411_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_col\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_137_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _04116_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__clkinv_4
XFILLER_153_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20558_ _09763_ _09859_ rbzero.traced_texVinit\[2\] _09762_ vssd1 vssd1 vccd1 vccd1
+ _01410_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_192_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10311_ rbzero.tex_r1\[62\] rbzero.tex_r1\[63\] _03483_ vssd1 vssd1 vccd1 vccd1 _03485_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11291_ rbzero.texV\[5\] _04070_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__xor2_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20489_ _03272_ _03386_ _03388_ _03250_ rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1
+ _01396_ sky130_fd_sc_hd__a32o_1
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13030_ _05725_ _05764_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a21bo_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14981_ rbzero.wall_tracer.stepDistX\[-3\] _07545_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07661_ sky130_fd_sc_hd__mux2_1
XFILLER_208_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16720_ _09352_ _09361_ vssd1 vssd1 vccd1 vccd1 _09362_ sky130_fd_sc_hd__xnor2_1
X_13932_ _06659_ _06664_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20247__267 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__inv_2
XFILLER_208_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13863_ _06335_ _06560_ _06562_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__and3_1
X_16651_ _05211_ _09138_ vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__or2_2
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12814_ _05533_ _05551_ _05553_ _05284_ rbzero.wall_tracer.mapY\[9\] vssd1 vssd1
+ vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
X_15602_ _08242_ _08239_ _08245_ _08246_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__o31a_1
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19370_ rbzero.wall_tracer.rayAddendY\[-3\] _02858_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _02859_ sky130_fd_sc_hd__mux2_1
X_13794_ _06511_ _06512_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__nand2_1
XFILLER_76_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16582_ _08821_ _08823_ _08419_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__or3_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18321_ _02017_ _02018_ _02019_ _05531_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a31o_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _05446_ _05447_ _05451_ _05449_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__o211a_1
X_15533_ _08177_ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__buf_4
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _08074_ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__buf_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18252_ _01841_ _01842_ _01844_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a21bo_1
XFILLER_203_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__nand2_2
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _07132_ _07151_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__xnor2_1
X_17203_ rbzero.wall_tracer.mapX\[7\] _09781_ _09779_ _09786_ vssd1 vssd1 vccd1 vccd1
+ _00572_ sky130_fd_sc_hd__a22o_1
XFILLER_175_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11627_ rbzero.tex_r1\[37\] rbzero.tex_r1\[36\] _04250_ vssd1 vssd1 vccd1 vccd1 _04406_
+ sky130_fd_sc_hd__mux2_1
XFILLER_187_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15395_ _05197_ rbzero.wall_tracer.stepDistX\[-9\] vssd1 vssd1 vccd1 vccd1 _08040_
+ sky130_fd_sc_hd__or2_2
X_18183_ _01646_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14346_ _07080_ _07082_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__xor2_1
X_17134_ rbzero.row_render.side _09762_ _07728_ _07895_ vssd1 vssd1 vccd1 vccd1 _00527_
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__buf_4
X_10509_ _03590_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17065_ _07602_ _09283_ _05210_ _09433_ vssd1 vssd1 vccd1 vccd1 _09705_ sky130_fd_sc_hd__or4_1
X_14277_ _06689_ _06668_ _06750_ _06748_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__o31a_1
XFILLER_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11489_ _04244_ _04256_ _04268_ _04116_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a31o_1
XFILLER_100_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16016_ _08574_ _08660_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__and2_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _05697_ _05792_ _05778_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__a21o_1
XFILLER_98_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _05802_ _05815_ _05884_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__mux2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17967_ _10183_ _09906_ _10294_ _01550_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__or4bb_4
XFILLER_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19706_ rbzero.pov.spi_buffer\[28\] rbzero.pov.spi_buffer\[29\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16918_ _09553_ _09558_ vssd1 vssd1 vccd1 vccd1 _09559_ sky130_fd_sc_hd__xnor2_2
XFILLER_66_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17898_ _01599_ _01600_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__and2b_1
XFILLER_77_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03306_ _03306_ vssd1 vssd1 vccd1 vccd1 clknet_0__03306_ sky130_fd_sc_hd__clkbuf_16
X_19637_ clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__buf_1
X_16849_ _08823_ _09164_ _09354_ vssd1 vssd1 vccd1 vccd1 _09490_ sky130_fd_sc_hd__or3_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19568_ rbzero.pov.spi_counter\[6\] _03034_ _03026_ vssd1 vssd1 vccd1 vccd1 _03036_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18519_ _02105_ _02115_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a21oi_1
X_19499_ _02952_ _02975_ _02976_ _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__nand4_1
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21530_ net451 _01299_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21461_ net382 _01230_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[40\] sky130_fd_sc_hd__dfxtp_1
X_20412_ _03324_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21392_ net313 _01161_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ _03775_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10791_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _03729_ vssd1 vssd1 vccd1 vccd1 _03739_
+ sky130_fd_sc_hd__mux2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _05205_ rbzero.map_rom.d6 _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__mux2_1
XFILLER_158_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _05214_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.trackDistY\[9\]
+ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a2bb2o_1
X_21659_ clknet_leaf_78_i_clk _01428_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14200_ _06926_ _06935_ _06936_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11412_ rbzero.row_render.size\[0\] gpout0.hpos\[0\] _04163_ vssd1 vssd1 vccd1 vccd1
+ _04192_ sky130_fd_sc_hd__a21o_1
Xtop_ew_algofoogle_72 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_72/HI o_rgb[0] sky130_fd_sc_hd__conb_1
X_15180_ _07785_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _07834_
+ sky130_fd_sc_hd__and2_1
X_12392_ net43 _05142_ _05144_ net42 _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
Xtop_ew_algofoogle_83 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_83/HI o_rgb[13] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_94 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_94/HI zeros[4] sky130_fd_sc_hd__conb_1
XFILLER_138_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _06828_ _06864_ _06865_ _06867_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_125_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ _04093_ _04114_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__or3_4
XFILLER_193_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14062_ _06722_ _06720_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__xnor2_1
X_11274_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _04054_ sky130_fd_sc_hd__or2_1
XFILLER_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13013_ _05601_ _05638_ _05649_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__or3_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18870_ _02543_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
X_17821_ _08263_ _08266_ _10134_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__and3_1
XFILLER_121_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5 rbzero.pov.spi_buffer\[32\] vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17752_ _10236_ _10252_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__nor2_1
XFILLER_208_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14964_ rbzero.wall_tracer.stepDistX\[-11\] _07465_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07652_ sky130_fd_sc_hd__mux2_1
XFILLER_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16703_ _09220_ _09344_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__nor2_1
X_13915_ _06645_ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17683_ _09674_ vssd1 vssd1 vccd1 vccd1 _10248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ rbzero.wall_tracer.visualWallDist\[-9\] _07595_ vssd1 vssd1 vccd1 vccd1 _07605_
+ sky130_fd_sc_hd__or2_1
XFILLER_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19422_ _02905_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__buf_4
XFILLER_78_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16634_ _09117_ _09276_ vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__nor2_1
XFILLER_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13846_ _06263_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__nor2_1
XFILLER_204_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19353_ _02840_ _02841_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or3_1
X_13777_ _06477_ _06479_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__xor2_1
X_16565_ _09188_ _09191_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__nor2_1
X_10989_ _03842_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18304_ _02001_ _02002_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__nand2_1
X_19581__38 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
XFILLER_128_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15516_ _08159_ _08160_ _08152_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__nor3_2
XFILLER_149_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12728_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__or2_1
X_19284_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_leak\[4\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
X_16496_ _09135_ _09139_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18235_ _01462_ _09480_ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__or3_1
XFILLER_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12659_ _05408_ rbzero.wall_tracer.mapY\[5\] _05283_ vssd1 vssd1 vccd1 vccd1 _05409_
+ sky130_fd_sc_hd__mux2_1
X_15447_ rbzero.debug_overlay.playerX\[-2\] _08027_ rbzero.debug_overlay.playerX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__o21ai_1
XFILLER_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18166_ _09434_ _09988_ _08802_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15378_ _07958_ _08022_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__nor2_1
XFILLER_184_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _04814_ _03474_ _04317_ vssd1 vssd1 vccd1 vccd1 _09754_ sky130_fd_sc_hd__a21o_1
X_14329_ _07062_ _07065_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18097_ _01792_ _01798_ rbzero.wall_tracer.trackDistX\[5\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00594_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17048_ _09684_ _09687_ vssd1 vssd1 vccd1 vccd1 _09688_ sky130_fd_sc_hd__xor2_1
XFILLER_104_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18999_ _02630_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20961_ clknet_leaf_69_i_clk _00730_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ clknet_leaf_82_i_clk _00661_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21513_ net434 _01282_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21444_ net365 _01213_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21375_ net296 _01144_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _04206_ _04736_ _04314_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a21o_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13700_ _06428_ _06435_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__nand2_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _03802_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__clkbuf_1
X_14680_ _07378_ _07413_ _06239_ _05779_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a211o_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11892_ rbzero.tex_b0\[15\] _04327_ _04328_ _04329_ vssd1 vssd1 vccd1 vccd1 _04668_
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ _06366_ _06354_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__and2b_1
X_10843_ _03766_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13562_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nand2_1
X_16350_ _08970_ _08994_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__xnor2_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10774_ _03730_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20359__368 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__inv_2
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12513_ rbzero.wall_tracer.trackDistX\[2\] vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__inv_2
X_15301_ rbzero.debug_overlay.playerX\[-4\] rbzero.debug_overlay.playerX\[-5\] _07898_
+ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__or3_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16281_ _08915_ _08925_ _08921_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__o21a_1
X_13493_ _06227_ _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__xor2_1
XFILLER_201_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18020_ _01720_ _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15232_ _07870_ _07873_ _07881_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__a21oi_1
X_12444_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__buf_2
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15163_ _07816_ _07817_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__nand2_1
X_12375_ _05141_ net32 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and2_1
XFILLER_154_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14114_ _06848_ _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__xnor2_1
X_11326_ _04103_ _04104_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__nor2_1
X_15094_ _07738_ _07752_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__nand2_1
X_19971_ rbzero.pov.ready_buffer\[22\] _03240_ _03243_ rbzero.debug_overlay.facingY\[-9\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__o221a_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14045_ _06774_ _06775_ _06780_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__a21o_1
X_18922_ _02574_ _02586_ _02587_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__and3_1
X_11257_ _04037_ rbzero.wall_tracer.state\[14\] vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__and2b_1
XFILLER_45_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18853_ _02527_ _02528_ _02406_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__o21a_1
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ rbzero.map_rom.f3 rbzero.map_rom.f2 rbzero.map_rom.i_col\[4\] vssd1 vssd1
+ vccd1 vccd1 _03977_ sky130_fd_sc_hd__or3_1
XFILLER_132_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17804_ _10099_ _10244_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__nand2_1
X_18784_ _02465_ _02466_ _02467_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__or3_1
XFILLER_209_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15996_ _08593_ _08595_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17735_ _05268_ _09781_ _01439_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__a21oi_1
X_14947_ rbzero.wall_tracer.visualWallDist\[7\] _07594_ vssd1 vssd1 vccd1 vccd1 _07641_
+ sky130_fd_sc_hd__or2_1
XFILLER_209_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17666_ _10214_ _10230_ vssd1 vssd1 vccd1 vccd1 _10231_ sky130_fd_sc_hd__xor2_1
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14878_ _04019_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19405_ _03913_ _02889_ _02890_ _07695_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a31o_1
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16617_ _09256_ _09258_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__and2_1
X_13829_ _06271_ _06269_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__or2b_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17597_ _10160_ _10162_ vssd1 vssd1 vccd1 vccd1 _10163_ sky130_fd_sc_hd__xor2_1
XFILLER_91_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19336_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__or2_1
X_16548_ _09188_ _09191_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__xor2_2
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19267_ _02787_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16479_ _09121_ _09122_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__xnor2_1
X_18218_ _01821_ _01853_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__or2_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19198_ rbzero.color_sky\[2\] _02740_ _02745_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__a21o_1
XFILLER_191_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18149_ _01848_ _01849_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__nor2_1
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21160_ clknet_leaf_84_i_clk _00929_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21091_ net181 _00860_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[31\] sky130_fd_sc_hd__dfxtp_1
X_20042_ _04886_ _03278_ _03280_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__o21ba_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20388__14 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20944_ clknet_leaf_67_i_clk _00713_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20875_ clknet_leaf_62_i_clk _00644_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10490_ rbzero.tex_r0\[44\] rbzero.tex_r0\[43\] _03580_ vssd1 vssd1 vccd1 vccd1 _03581_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21427_ net348 _01196_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12160_ _04918_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__inv_2
XFILLER_163_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21358_ net279 _01127_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11111_ _03906_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12091_ net68 _04857_ _04838_ _04323_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a22o_1
X_21289_ clknet_leaf_42_i_clk _01058_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _03870_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15850_ _08113_ _08139_ _08140_ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__o21bai_1
XFILLER_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _00004_ _07530_ _07531_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a21oi_1
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _08135_ _08422_ _08425_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__or3_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _05638_ _05695_ _05677_ _05681_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or4_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17520_ _10051_ _10052_ _10084_ vssd1 vssd1 vccd1 vccd1 _10086_ sky130_fd_sc_hd__nand3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _05834_ _07455_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__and2_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _04356_ vssd1 vssd1 vccd1 vccd1 _04720_
+ sky130_fd_sc_hd__mux2_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17451_ _10015_ _10017_ vssd1 vssd1 vccd1 vccd1 _10018_ sky130_fd_sc_hd__xnor2_2
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14663_ _07388_ _07381_ _05931_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__mux2_1
X_11875_ _04648_ _04651_ _04209_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__mux2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _09045_ _09046_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__nand2_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13614_ _06305_ _06321_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__xor2_2
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10826_ _03757_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17382_ _09639_ _09646_ _09948_ vssd1 vssd1 vccd1 vccd1 _09949_ sky130_fd_sc_hd__a21oi_2
X_14594_ _07329_ _07330_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__and2b_1
XFILLER_186_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19121_ _03555_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__buf_6
X_16333_ _07598_ _08230_ _08147_ _08236_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__or4_1
X_13545_ _06065_ _06134_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__or2_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10757_ _03721_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19052_ rbzero.pov.spi_buffer\[57\] rbzero.pov.ready_buffer\[57\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
X_13476_ _06179_ _06181_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__and2b_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16264_ _08897_ _08906_ _08905_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__a21o_1
X_10688_ rbzero.tex_g1\[13\] rbzero.tex_g1\[14\] _03680_ vssd1 vssd1 vccd1 vccd1 _03685_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18003_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15215_ _07865_ _07866_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__or2_1
X_12427_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__clkbuf_8
XFILLER_154_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16195_ _08831_ _08837_ _08839_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__a21oi_1
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12358_ net52 _05103_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a21oi_1
X_15146_ _07730_ rbzero.debug_overlay.vplaneX\[-5\] _07800_ _07801_ vssd1 vssd1 vccd1
+ vccd1 _07802_ sky130_fd_sc_hd__o22a_1
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _04082_ _04088_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nor2_2
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15077_ rbzero.debug_overlay.vplaneX\[-6\] _07708_ _07736_ _07737_ vssd1 vssd1 vccd1
+ vccd1 _07738_ sky130_fd_sc_hd__a2bb2o_1
X_19954_ rbzero.pov.ready_buffer\[35\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-7\]
+ _03209_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__o221a_1
X_12289_ net43 _05043_ _05044_ net41 net23 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a221o_1
X_14028_ _05982_ _06740_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nor2_1
X_18905_ rbzero.spi_registers.spi_counter\[0\] _02558_ vssd1 vssd1 vccd1 vccd1 _02575_
+ sky130_fd_sc_hd__or2_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19885_ net39 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__o21ai_2
X_20112__145 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__inv_2
XFILLER_110_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18836_ _02510_ _02511_ _02512_ _04016_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a31o_1
XFILLER_209_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18767_ _02452_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__xnor2_1
X_15979_ _07958_ _08128_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__nor2_1
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17718_ _10088_ _10155_ _10282_ vssd1 vssd1 vccd1 vccd1 _10283_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18698_ _05532_ _02393_ _09817_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__o21a_1
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _10204_ _10213_ vssd1 vssd1 vccd1 vccd1 _10214_ sky130_fd_sc_hd__xor2_1
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20660_ clknet_leaf_10_i_clk _00444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-11\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_211_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19319_ rbzero.spi_registers.new_vshift\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20591_ _07679_ _02830_ _03458_ _07855_ rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__a32o_1
XFILLER_91_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21212_ clknet_leaf_18_i_clk _00981_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21143_ clknet_leaf_61_i_clk _00912_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21074_ net164 _00843_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20025_ _04892_ _04992_ _04037_ _03911_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a31o_1
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20087__122 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__inv_2
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ clknet_leaf_13_i_clk _00696_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11660_ _04004_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__and2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ clknet_leaf_55_i_clk _00627_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10611_ rbzero.tex_g1\[49\] rbzero.tex_g1\[50\] _03635_ vssd1 vssd1 vccd1 vccd1 _03644_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11591_ _04225_ _04367_ _04368_ _04369_ _04208_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o221a_1
XFILLER_161_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20789_ clknet_leaf_21_i_clk _00558_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13330_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__buf_2
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10542_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _03602_ vssd1 vssd1 vccd1 vccd1 _03608_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13261_ _05977_ _05987_ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ rbzero.tex_r0\[52\] rbzero.tex_r0\[51\] _03569_ vssd1 vssd1 vccd1 vccd1 _03572_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12212_ net42 _04963_ _04980_ _04981_ _04021_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a32o_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15000_ _07670_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13192_ _05703_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nor2_2
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12143_ _04910_ net64 _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a21bo_1
XFILLER_194_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12074_ net5 net6 vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nand2_1
X_16951_ _09454_ _09591_ vssd1 vssd1 vccd1 vccd1 _09592_ sky130_fd_sc_hd__and2_1
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _03861_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__clkbuf_1
X_15902_ _08470_ _08546_ vssd1 vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__nor2_2
XFILLER_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19670_ _03061_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16882_ _08282_ _08129_ _08047_ _09522_ vssd1 vssd1 vccd1 vccd1 _09523_ sky130_fd_sc_hd__o22ai_1
X_18621_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__nand2_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _08472_ _08477_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__or2b_1
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18552_ _02141_ _02248_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__xor2_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _08402_ _08408_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__xnor2_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__xor2_2
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _10067_ _10068_ vssd1 vssd1 vccd1 vccd1 _10069_ sky130_fd_sc_hd__and2_1
XFILLER_73_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14715_ _07419_ _07420_ _07106_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__a21o_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _04701_ _04702_ _04266_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__mux2_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _02179_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__and2_1
X_15695_ _08338_ _08339_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__or2_1
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _09707_ _09708_ _09706_ vssd1 vssd1 vccd1 vccd1 _10001_ sky130_fd_sc_hd__o21a_1
X_14646_ _07106_ _07379_ _07380_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__a31o_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11858_ rbzero.tex_g1\[10\] _04291_ _04329_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a21o_1
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 _09194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _03748_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
X_17365_ _09368_ _09165_ _09628_ _09629_ vssd1 vssd1 vccd1 vccd1 _09932_ sky130_fd_sc_hd__o31a_1
X_14577_ _07295_ _07306_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__nor2_1
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11789_ _04565_ _04566_ _04345_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__mux2_1
X_19104_ _02685_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16316_ _08192_ _08960_ _08179_ _08190_ vssd1 vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_201_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13528_ _06263_ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__and2_1
XFILLER_186_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17296_ _09864_ _09865_ _09866_ vssd1 vssd1 vccd1 vccd1 _09868_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19035_ _02593_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__clkbuf_4
X_16247_ _08889_ _08891_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__xor2_1
X_13459_ _06194_ _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__nand2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16178_ _08112_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15129_ _07785_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _07786_
+ sky130_fd_sc_hd__nand2_1
XFILLER_141_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_92_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19937_ _03193_ _03230_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1
+ _03231_ sky130_fd_sc_hd__o21a_1
X_19868_ rbzero.pov.ready_buffer\[70\] _02823_ _03138_ _03178_ vssd1 vssd1 vccd1 vccd1
+ _03179_ sky130_fd_sc_hd__a211o_1
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18819_ _02497_ _02498_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__nand2_1
X_19799_ _03128_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03299_ clknet_0__03299_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03299_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20712_ clknet_leaf_15_i_clk _00003_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20643_ clknet_leaf_8_i_clk _00427_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20574_ gpout1.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__nor2_1
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21126_ clknet_leaf_66_i_clk _00895_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21057_ clknet_leaf_56_i_clk _00826_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20008_ _02595_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__and2_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _05563_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__nand2_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__xor2_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14500_ _07222_ _07224_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__xnor2_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ rbzero.debug_overlay.facingX\[-4\] _04464_ _04465_ rbzero.debug_overlay.facingX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a22o_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _05196_ rbzero.wall_tracer.stepDistX\[-10\] _08053_ vssd1 vssd1 vccd1 vccd1
+ _08125_ sky130_fd_sc_hd__o21bai_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12692_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__or2_1
XFILLER_188_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14431_ _07164_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__or2_1
X_11643_ _04045_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nand2_2
X_20141__171 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__inv_2
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17150_ _07706_ vssd1 vssd1 vccd1 vccd1 _09766_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14362_ _07043_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__and2_1
X_11574_ _04349_ _04351_ _04352_ _04225_ _04253_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o221a_1
XFILLER_195_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 i_gpout2_sel[3] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_8
Xinput28 i_gpout4_sel[2] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_6
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16101_ _08594_ _07938_ vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__nor2_1
X_13313_ _06039_ _06048_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__o21ai_1
X_10525_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _03591_ vssd1 vssd1 vccd1 vccd1 _03599_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 i_mode[1] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_16
X_14293_ _07027_ _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__xor2_2
XFILLER_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17081_ _09718_ _09720_ vssd1 vssd1 vccd1 vccd1 _09721_ sky130_fd_sc_hd__xor2_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13244_ _05941_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__and2_1
X_16032_ _07988_ _08674_ _08020_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__or3_1
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10456_ rbzero.tex_r0\[60\] rbzero.tex_r0\[59\] _03558_ vssd1 vssd1 vccd1 vccd1 _03563_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13175_ _05826_ _05911_ _05755_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a21o_1
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10387_ _03524_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _03555_ _04857_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a21o_2
X_17983_ _01663_ _01560_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__or2b_1
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19722_ _03088_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
X_12057_ _03474_ _04809_ _04810_ _04818_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a41o_1
X_16934_ _09550_ _09574_ vssd1 vssd1 vccd1 vccd1 _09575_ sky130_fd_sc_hd__xnor2_2
XFILLER_78_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11008_ _03852_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19653_ _03052_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16865_ _09500_ _09505_ vssd1 vssd1 vccd1 vccd1 _09506_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18604_ _02291_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__xor2_1
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15816_ _08145_ _08122_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16796_ _09436_ _09437_ vssd1 vssd1 vccd1 vccd1 _09438_ sky130_fd_sc_hd__xnor2_2
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ _02229_ _02230_ _02231_ _05531_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a31o_1
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15747_ _07943_ _07968_ _07942_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__a21bo_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20224__246 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__inv_2
XFILLER_92_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12959_ _05638_ _05682_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__or2_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18466_ _02083_ _02097_ _02096_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a21o_1
X_15678_ _08320_ _08322_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17417_ _09982_ _09983_ vssd1 vssd1 vccd1 vccd1 _09984_ sky130_fd_sc_hd__xnor2_2
X_14629_ _05793_ _07365_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__nand2_1
XFILLER_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18397_ _02093_ _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__nor2_1
XFILLER_193_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17348_ _09654_ _09909_ _09914_ vssd1 vssd1 vccd1 vccd1 _09915_ sky130_fd_sc_hd__a21oi_1
XFILLER_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17279_ rbzero.wall_tracer.trackDistX\[-7\] _09852_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09853_ sky130_fd_sc_hd__mux2_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19018_ _02640_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20270__288 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__inv_2
XFILLER_138_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_opt_5_0_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_5_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20199__223 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__inv_2
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03311_ clknet_0__03311_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03311_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20626_ clknet_leaf_51_i_clk _00410_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f1 sky130_fd_sc_hd__dfxtp_1
XFILLER_196_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20557_ rbzero.traced_texVinit\[1\] _03443_ _09771_ _09076_ vssd1 vssd1 vccd1 vccd1
+ _01409_ sky130_fd_sc_hd__a22o_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10310_ _03484_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ _04067_ _04066_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__nand2_1
XFILLER_180_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20488_ _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__inv_2
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21109_ net199 _00878_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[49\] sky130_fd_sc_hd__dfxtp_1
X_14980_ _05201_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__buf_4
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13931_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16650_ _08239_ _09292_ _09289_ _09290_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__a2bb2o_1
X_13862_ _06277_ _06563_ _06597_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__or3b_1
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15601_ _08243_ _08244_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__or2_1
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ _05548_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__or2b_1
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16581_ _09092_ _09095_ vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__nand2_1
X_13793_ _05855_ _06061_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__nand2_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18320_ _02017_ _02018_ _02019_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a21oi_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _08147_ rbzero.wall_tracer.stepDistX\[1\] _08175_ _08176_ vssd1 vssd1 vccd1
+ vccd1 _08177_ sky130_fd_sc_hd__a22oi_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and2_1
XFILLER_63_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _01949_ _01950_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__and2_1
XFILLER_43_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15463_ _08106_ _08107_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__or2_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__nor2_1
X_17202_ _09782_ _09785_ vssd1 vssd1 vccd1 vccd1 _09786_ sky130_fd_sc_hd__xnor2_1
X_14414_ _07072_ _07148_ _07150_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__and3b_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11626_ rbzero.tex_r1\[39\] rbzero.tex_r1\[38\] _04250_ vssd1 vssd1 vccd1 vccd1 _04405_
+ sky130_fd_sc_hd__mux2_1
X_18182_ _01877_ _01882_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__xnor2_1
X_15394_ _07925_ _08037_ _08038_ vssd1 vssd1 vccd1 vccd1 _08039_ sky130_fd_sc_hd__a21o_2
XFILLER_196_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _07706_ vssd1 vssd1 vccd1 vccd1 _09762_ sky130_fd_sc_hd__buf_4
X_14345_ _07015_ _07022_ _07081_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a21oi_1
XFILLER_200_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11557_ _04128_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__buf_4
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10508_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _03580_ vssd1 vssd1 vccd1 vccd1 _03590_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17064_ _05198_ _09703_ vssd1 vssd1 vccd1 vccd1 _09704_ sky130_fd_sc_hd__nand2_2
X_11488_ _04258_ _04260_ _04267_ _04210_ _04242_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__a221o_1
X_14276_ _07007_ _07012_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__xnor2_2
XFILLER_183_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16015_ _08111_ _08579_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__nor2_1
X_10439_ rbzero.tex_r1\[1\] rbzero.tex_r1\[2\] _03549_ vssd1 vssd1 vccd1 vccd1 _03552_
+ sky130_fd_sc_hd__mux2_1
X_13227_ _05743_ _05874_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__o21a_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _05891_ _05892_ _05591_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12109_ _04874_ _04876_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__and3_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13089_ _05795_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__clkbuf_4
X_17966_ _01667_ _01668_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__nand2_1
XFILLER_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19705_ _03079_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__clkbuf_1
X_16917_ _09556_ _09557_ vssd1 vssd1 vccd1 vccd1 _09558_ sky130_fd_sc_hd__nand2_1
X_17897_ _01593_ _01598_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__03305_ _03305_ vssd1 vssd1 vccd1 vccd1 clknet_0__03305_ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16848_ _08823_ _09028_ _09164_ _08329_ vssd1 vssd1 vccd1 vccd1 _09489_ sky130_fd_sc_hd__o22a_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19567_ _03034_ _03035_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__nor2_1
XFILLER_81_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16779_ _09141_ _09420_ _08170_ vssd1 vssd1 vccd1 vccd1 _09421_ sky130_fd_sc_hd__a21oi_1
XFILLER_209_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18518_ _02102_ _02104_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__nor2_1
XFILLER_94_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19498_ rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\] _02905_
+ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__o21ai_1
XFILLER_179_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18449_ _02145_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__nand2_1
XFILLER_179_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21460_ net381 _01229_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20411_ _02721_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__and3_1
XFILLER_146_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21391_ net312 _01160_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20207__230 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__inv_2
XFILLER_44_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _03738_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21658_ clknet_leaf_88_i_clk _01427_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12460_ rbzero.wall_tracer.trackDistX\[9\] vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__inv_2
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ gpout0.hpos\[2\] _04149_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nand3b_1
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20609_ _03469_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__clkbuf_1
X_12391_ net41 _05139_ net34 net35 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a211o_1
XFILLER_123_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_73 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_73/HI o_rgb[1] sky130_fd_sc_hd__conb_1
X_21589_ net130 _01358_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_84 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_84/HI o_rgb[16] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_95 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_95/HI zeros[5] sky130_fd_sc_hd__conb_1
XFILLER_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14130_ _06828_ _06864_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__a21o_1
X_11342_ _04092_ _04081_ _04089_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__nor3_2
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20253__272 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__inv_2
X_14061_ _06757_ _06797_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__xnor2_1
X_11273_ _04048_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nand2_1
XFILLER_181_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13012_ _05695_ _05702_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__or3_1
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17820_ _10129_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__buf_2
XFILLER_95_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _10214_ _10230_ _10228_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a21o_1
X_14963_ _07651_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16702_ _09210_ _09237_ _09343_ vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__a21boi_1
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13914_ _06572_ _06627_ _06629_ _06650_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__o211a_1
XFILLER_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17682_ _10245_ _10246_ vssd1 vssd1 vccd1 vccd1 _10247_ sky130_fd_sc_hd__xor2_1
XFILLER_75_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14894_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.trackDistX\[-9\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__mux2_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19421_ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__buf_2
X_16633_ _08971_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__buf_4
X_13845_ _06248_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19352_ _02824_ _02837_ _02825_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__o21ai_2
X_16564_ _08549_ _08957_ _09204_ _09206_ vssd1 vssd1 vccd1 vccd1 _09207_ sky130_fd_sc_hd__a31o_2
XFILLER_204_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13776_ _06406_ _06511_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__a21bo_1
XFILLER_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10988_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _03762_ vssd1 vssd1 vccd1 vccd1 _03842_
+ sky130_fd_sc_hd__mux2_1
XFILLER_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18303_ _02001_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__nor2_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15515_ _08124_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__clkbuf_4
X_12727_ _05473_ _05474_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__xnor2_4
X_19283_ _02796_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16495_ _08816_ _09138_ vssd1 vssd1 vccd1 vccd1 _09139_ sky130_fd_sc_hd__nor2_1
XFILLER_203_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18234_ _09661_ _09483_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__or2_1
XFILLER_188_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15446_ rbzero.wall_tracer.visualWallDist\[-1\] _08090_ _07951_ vssd1 vssd1 vccd1
+ vccd1 _08091_ sky130_fd_sc_hd__mux2_1
X_12658_ rbzero.debug_overlay.playerY\[5\] _05407_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05408_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20336__347 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__inv_2
X_11609_ rbzero.tex_r1\[55\] _04221_ _04222_ _04266_ vssd1 vssd1 vccd1 vccd1 _04388_
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18165_ _09292_ _09695_ _09668_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a21o_1
XFILLER_191_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15377_ _08021_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__clkbuf_2
X_12589_ _05289_ _05295_ _05303_ _05301_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a31o_1
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _05189_ vssd1 vssd1 vccd1 vccd1 _09753_ sky130_fd_sc_hd__clkbuf_4
X_14328_ _07063_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18096_ _01796_ _01797_ _09817_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__o21a_1
XFILLER_102_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _09685_ _09686_ vssd1 vssd1 vccd1 vccd1 _09687_ sky130_fd_sc_hd__xnor2_1
X_14259_ _06724_ _06672_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__nor2_1
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19629__81 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__inv_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ rbzero.pov.spi_buffer\[31\] rbzero.pov.ready_buffer\[31\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XFILLER_86_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17949_ _01650_ _01651_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__and2b_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20960_ clknet_leaf_68_i_clk _00729_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20081__117 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__inv_2
XFILLER_54_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20891_ clknet_leaf_82_i_clk _00660_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21512_ net433 _01281_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21443_ net364 _01212_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21374_ net295 _01143_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ rbzero.color_sky\[4\] rbzero.color_floor\[4\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04736_ sky130_fd_sc_hd__mux2_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ rbzero.tex_b1\[35\] rbzero.tex_b1\[36\] _03795_ vssd1 vssd1 vccd1 vccd1 _03802_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ rbzero.tex_b0\[14\] _04291_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and2_1
XFILLER_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ _06354_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10842_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _03762_ vssd1 vssd1 vccd1 vccd1 _03766_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13561_ _06078_ _06161_ _06292_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__o31a_1
XFILLER_164_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10773_ rbzero.tex_g0\[38\] rbzero.tex_g0\[37\] _03729_ vssd1 vssd1 vccd1 vccd1 _03730_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15300_ _05207_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__buf_6
XFILLER_160_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ rbzero.wall_tracer.trackDistX\[-3\] vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__inv_2
XFILLER_185_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16280_ _08918_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__inv_2
X_13492_ _06175_ _06185_ _06228_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ _07821_ rbzero.wall_tracer.rayAddendX\[10\] vssd1 vssd1 vccd1 vccd1 _07881_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_201_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12443_ net71 rbzero.wall_tracer.state\[4\] _03480_ vssd1 vssd1 vccd1 vccd1 _05200_
+ sky130_fd_sc_hd__and3_1
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15162_ _07785_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _07817_
+ sky130_fd_sc_hd__or2_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12374_ net33 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__inv_2
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14113_ _06691_ _06849_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _04103_ _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15093_ _07738_ _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__or2_1
X_19970_ rbzero.pov.ready_buffer\[43\] _03240_ _03243_ rbzero.debug_overlay.facingX\[10\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__o221a_1
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14044_ _06774_ _06775_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and3_1
XFILLER_158_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_141_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18921_ rbzero.spi_registers.spi_counter\[4\] _02583_ vssd1 vssd1 vccd1 vccd1 _02587_
+ sky130_fd_sc_hd__or2_1
XFILLER_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18852_ _02524_ _02525_ _02526_ _05531_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a31o_1
X_11187_ _03974_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__nand2_1
X_17803_ _01505_ _01506_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__xor2_2
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18783_ _02465_ _02466_ _02467_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__o21a_1
X_15995_ _08633_ _08632_ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__xor2_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17734_ _09812_ _10181_ _10182_ _05414_ _01438_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__o311a_1
XFILLER_48_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14946_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.trackDistX\[7\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__mux2_1
XFILLER_82_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _10228_ _10229_ vssd1 vssd1 vccd1 vccd1 _10230_ sky130_fd_sc_hd__nor2_1
X_14877_ _07590_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19404_ _02883_ _02888_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__nand2_1
X_16616_ _09256_ _09258_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__nor2_1
X_13828_ _06268_ _06235_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__or2b_1
X_17596_ _09918_ _10018_ _10161_ vssd1 vssd1 vccd1 vccd1 _10162_ sky130_fd_sc_hd__a21boi_1
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16547_ _09053_ _09189_ _09190_ vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__a21oi_2
X_19335_ _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__and2b_1
X_13759_ _06461_ _06458_ _06465_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__a211o_1
XFILLER_188_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19266_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_floor\[3\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_203_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16478_ _08383_ _07959_ vssd1 vssd1 vccd1 vccd1 _09122_ sky130_fd_sc_hd__nor2_1
XFILLER_188_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18217_ _01688_ _01690_ _01816_ _01814_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a31o_1
X_15429_ _05206_ _08068_ _08072_ _08073_ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__a22o_2
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19197_ rbzero.spi_registers.new_sky\[2\] rbzero.spi_registers.got_new_sky _02711_
+ _02741_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a31o_1
XFILLER_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18148_ _01716_ _01725_ _01724_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__o21ba_1
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18079_ _01697_ _01780_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21090_ net180 _00859_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20041_ _04886_ _04990_ _03275_ _03911_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__a31o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ clknet_leaf_67_i_clk _00712_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_187_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ clknet_leaf_62_i_clk _00643_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20319__331 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__inv_2
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21426_ net347 _01195_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21357_ net278 _01126_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11110_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _03898_ vssd1 vssd1 vccd1 vccd1 _03906_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12090_ _04851_ _04856_ _04861_ _04850_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a22o_1
XFILLER_155_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21288_ clknet_leaf_31_i_clk _01057_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11041_ rbzero.tex_b0\[38\] rbzero.tex_b0\[37\] _03865_ vssd1 vssd1 vccd1 vccd1 _03870_
+ sky130_fd_sc_hd__mux2_1
X_19608__62 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ rbzero.wall_tracer.stepDistY\[-6\] _07461_ vssd1 vssd1 vccd1 vccd1 _07531_
+ sky130_fd_sc_hd__nor2_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20365__373 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__inv_2
X_19623__76 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _08424_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__buf_2
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _05728_ _05645_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__nand2_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20064__101 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__inv_2
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _07466_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__clkbuf_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _04717_ _04718_ _04329_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__mux2_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17450_ _09657_ _09725_ _10016_ vssd1 vssd1 vccd1 vccd1 _10017_ sky130_fd_sc_hd__a21o_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _05892_ _07395_ _07398_ _07375_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__o211a_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11874_ _04649_ _04650_ _04224_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__mux2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16401_ _08367_ _09026_ _09044_ vssd1 vssd1 vccd1 vccd1 _09046_ sky130_fd_sc_hd__nand3_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _06345_ _06346_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__xnor2_1
X_10825_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _03751_ vssd1 vssd1 vccd1 vccd1 _03757_
+ sky130_fd_sc_hd__mux2_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _09521_ _09525_ _09645_ vssd1 vssd1 vccd1 vccd1 _09948_ sky130_fd_sc_hd__a21oi_1
X_14593_ _07213_ _07328_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__nand2_1
XFILLER_125_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19120_ _02694_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__clkbuf_1
X_16332_ _07602_ _08230_ _08147_ _08225_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__or4b_2
X_13544_ _06132_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__xor2_2
XFILLER_164_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10756_ rbzero.tex_g0\[46\] rbzero.tex_g0\[45\] _03718_ vssd1 vssd1 vccd1 vccd1 _03721_
+ sky130_fd_sc_hd__mux2_1
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _02657_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
X_16263_ _08897_ _08907_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__xor2_1
XFILLER_199_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13475_ _05910_ _06176_ _06085_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__and3_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ _03684_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18002_ _09249_ _09703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__and2_1
XFILLER_185_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15214_ _07843_ _07845_ _07864_ _07676_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__a31o_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ _03480_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__buf_4
XFILLER_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16194_ _08793_ _08838_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__or2_1
XFILLER_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15145_ _07742_ rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 _07801_
+ sky130_fd_sc_hd__and2_1
X_12357_ net49 _05084_ _05107_ net50 vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a22o_1
XFILLER_153_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _04084_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__or2_2
X_15076_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__nand2_1
X_19953_ rbzero.pov.ready_buffer\[34\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-8\]
+ _03209_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__o221a_1
X_12288_ net39 _05046_ _05049_ net40 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a22o_1
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14027_ _06704_ _06761_ _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__or3_1
X_18904_ _02557_ _02573_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__and2_1
X_11239_ gpout0.hpos\[2\] gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _04023_ sky130_fd_sc_hd__and3_2
X_19884_ _03189_ _03191_ _02714_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__o21a_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18835_ _02510_ _02511_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a21oi_1
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18766_ _02443_ _02445_ _02444_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a21boi_1
X_15978_ _07912_ _08328_ _08040_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__or3b_2
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17717_ _10152_ _10154_ vssd1 vssd1 vccd1 vccd1 _10282_ sky130_fd_sc_hd__nor2_1
X_14929_ rbzero.wall_tracer.visualWallDist\[1\] _07618_ vssd1 vssd1 vccd1 vccd1 _07629_
+ sky130_fd_sc_hd__or2_1
XFILLER_209_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18697_ _02391_ _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17648_ _10211_ _10212_ vssd1 vssd1 vccd1 vccd1 _10213_ sky130_fd_sc_hd__nor2_1
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17579_ _10127_ _10136_ _10142_ _10144_ vssd1 vssd1 vccd1 vccd1 _10145_ sky130_fd_sc_hd__o22a_1
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19318_ _02815_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20590_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__or2_1
XFILLER_56_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20193__218 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__inv_2
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _02777_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21211_ clknet_leaf_17_i_clk _00980_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21142_ clknet_leaf_61_i_clk _00911_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21073_ net163 _00842_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20024_ _04992_ _03267_ _03268_ _03209_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__o211a_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ clknet_leaf_13_i_clk _00695_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20857_ clknet_leaf_57_i_clk _00626_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _03643_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11590_ rbzero.tex_r1\[30\] _04350_ _04265_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__a21o_1
X_20788_ clknet_leaf_20_i_clk _00557_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _03607_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13260_ _05993_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__or2b_1
XFILLER_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10472_ _03571_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12211_ _04960_ _04961_ _04963_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__and3_1
XFILLER_109_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21409_ net330 _01178_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13191_ _05743_ _05754_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nor2_2
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _04910_ _04738_ net12 net11 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o211a_1
XFILLER_159_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12073_ _04840_ net66 _04844_ net6 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a211o_1
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16950_ _09345_ _09590_ vssd1 vssd1 vccd1 vccd1 _09591_ sky130_fd_sc_hd__xor2_1
X_15901_ _08509_ _08544_ _08545_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__a21oi_1
X_11024_ rbzero.tex_b0\[46\] rbzero.tex_b0\[45\] _03854_ vssd1 vssd1 vccd1 vccd1 _03861_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16881_ _07994_ vssd1 vssd1 vccd1 vccd1 _09522_ sky130_fd_sc_hd__buf_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15832_ _08473_ _08474_ _08476_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__a21bo_1
X_18620_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__or2_1
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15763_ _08406_ _08407_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__nand2_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _02236_ _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _05594_ _05596_ _05598_ _05584_ _05628_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__o41a_2
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _07348_ _07353_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__nand2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _10057_ _10066_ vssd1 vssd1 vccd1 vccd1 _10068_ sky130_fd_sc_hd__or2_1
X_11926_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _04263_ vssd1 vssd1 vccd1 vccd1 _04702_
+ sky130_fd_sc_hd__mux2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _02176_ _02178_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__nand2_1
XFILLER_166_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15694_ _08084_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__or3_1
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _09700_ _09997_ _09998_ _09999_ vssd1 vssd1 vccd1 vccd1 _10000_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _05931_ _07381_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nor2_1
XFILLER_33_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11857_ rbzero.tex_g1\[11\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__and3_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10808_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _03740_ vssd1 vssd1 vccd1 vccd1 _03748_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17364_ _09929_ _09930_ vssd1 vssd1 vccd1 vccd1 _09931_ sky130_fd_sc_hd__xor2_1
XFILLER_186_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14576_ _07095_ _07035_ _07043_ _07098_ _07312_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__a221o_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _04262_ vssd1 vssd1 vccd1 vccd1 _04566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19103_ rbzero.spi_registers.spi_buffer\[7\] rbzero.spi_registers.spi_buffer\[6\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
X_16315_ _08008_ _08204_ vssd1 vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__or2_1
X_13527_ _06256_ _06257_ _06262_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__or3_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17295_ _09864_ _09865_ _09866_ vssd1 vssd1 vccd1 vccd1 _09867_ sky130_fd_sc_hd__and3_1
X_10739_ _03711_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19034_ _02648_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__clkbuf_1
X_16246_ _08879_ _08883_ _08890_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__a21oi_1
X_13458_ _06191_ _06189_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__or2b_1
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ _05171_ _05175_ net36 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or3b_1
X_16177_ _08112_ _08328_ _08747_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__or3_1
X_13389_ _06121_ _06124_ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__and3_1
XFILLER_138_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15128_ rbzero.debug_overlay.vplaneX\[10\] vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15059_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__or2_1
X_19936_ _02820_ _03227_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__nor2_1
XFILLER_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19867_ _03176_ _03177_ _02822_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18818_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__or2_1
XFILLER_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19798_ rbzero.pov.spi_buffer\[72\] rbzero.pov.spi_buffer\[73\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
XFILLER_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19602__57 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
X_18749_ _02435_ _02436_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nor3_1
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03298_ clknet_0__03298_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03298_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_209_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20711_ clknet_leaf_11_i_clk _00002_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20201__225 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__inv_2
XFILLER_149_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20642_ clknet_leaf_26_i_clk _00426_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20573_ _03447_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_opt_1_0_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21125_ clknet_leaf_65_i_clk _00894_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21056_ clknet_leaf_57_i_clk _00825_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20007_ _03020_ _03019_ _03025_ rbzero.pov.spi_done vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__a31o_1
XFILLER_87_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _03924_ _05503_ _05499_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__o21ai_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _04481_ _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__nand2_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20909_ clknet_leaf_79_i_clk _00678_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_12691_ _05421_ _05430_ _05433_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a31o_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14430_ _07137_ _07045_ _07165_ _07166_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11642_ _04414_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__inv_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20176__202 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__inv_2
XFILLER_211_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14361_ _07095_ _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ rbzero.tex_r1\[1\] rbzero.tex_r1\[0\] _04342_ vssd1 vssd1 vccd1 vccd1 _04352_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 i_gpout2_sel[4] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_6
X_16100_ _08519_ _08075_ _08674_ _08377_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__o22ai_2
X_13312_ _06022_ _06038_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nand2_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10524_ _03598_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 i_gpout4_sel[3] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_8
X_17080_ _09550_ _09574_ _09719_ vssd1 vssd1 vccd1 vccd1 _09720_ sky130_fd_sc_hd__a21oi_2
XFILLER_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14292_ _06737_ _06817_ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__a21boi_2
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16031_ _07980_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__or3_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13243_ _05979_ _05899_ _05846_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__o21ai_2
XFILLER_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10455_ _03562_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ _05867_ _05783_ _05792_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__mux2_1
XFILLER_124_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ rbzero.tex_r1\[26\] rbzero.tex_r1\[27\] _03516_ vssd1 vssd1 vccd1 vccd1 _03524_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ _04852_ clknet_1_0__leaf__04835_ _04855_ gpout0.clk_div\[1\] _04838_ vssd1
+ vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a221o_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ _01660_ _01662_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__or2_1
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19721_ rbzero.pov.spi_buffer\[35\] rbzero.pov.spi_buffer\[36\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12056_ _04819_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__nor2_1
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16933_ _09571_ _09573_ vssd1 vssd1 vccd1 vccd1 _09574_ sky130_fd_sc_hd__xnor2_2
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03321_ _03321_ vssd1 vssd1 vccd1 vccd1 clknet_0__03321_ sky130_fd_sc_hd__clkbuf_16
X_11007_ rbzero.tex_b0\[54\] rbzero.tex_b0\[53\] _03843_ vssd1 vssd1 vccd1 vccd1 _03852_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19652_ rbzero.pov.spi_buffer\[2\] rbzero.pov.spi_buffer\[3\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03052_ sky130_fd_sc_hd__mux2_1
X_16864_ _09501_ _09504_ vssd1 vssd1 vccd1 vccd1 _09505_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18603_ _02208_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__xnor2_1
X_15815_ _08441_ _08459_ vssd1 vssd1 vccd1 vccd1 _08460_ sky130_fd_sc_hd__xor2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16795_ _09290_ _09291_ vssd1 vssd1 vccd1 vccd1 _09437_ sky130_fd_sc_hd__nand2_1
XFILLER_206_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15746_ _08373_ _08390_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__xnor2_1
X_18534_ _02229_ _02230_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a21oi_1
X_12958_ _05674_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__buf_2
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11909_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _04271_ vssd1 vssd1 vccd1 vccd1 _04685_
+ sky130_fd_sc_hd__mux2_1
XFILLER_206_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15677_ _08321_ _08286_ vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__xnor2_1
X_18465_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__xor2_1
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12889_ _04001_ _05456_ _05624_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a22oi_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14628_ _07363_ _07364_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__xnor2_2
X_17416_ _09114_ _09417_ vssd1 vssd1 vccd1 vccd1 _09983_ sky130_fd_sc_hd__nor2_1
X_18396_ _01952_ _01959_ _02094_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ _09912_ _09913_ vssd1 vssd1 vccd1 vccd1 _09914_ sky130_fd_sc_hd__or2_1
XFILLER_202_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14559_ _07289_ _07290_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__or2_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _09812_ _09849_ _09850_ _09851_ vssd1 vssd1 vccd1 vccd1 _09852_ sky130_fd_sc_hd__o31ai_1
XFILLER_88_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19017_ rbzero.pov.spi_buffer\[40\] rbzero.pov.ready_buffer\[40\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
X_16229_ _08872_ _08491_ _08579_ _08873_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__o22a_1
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19919_ rbzero.debug_overlay.playerY\[0\] _08030_ vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__nand2_1
XFILLER_151_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03310_ clknet_0__03310_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03310_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20625_ clknet_leaf_52_i_clk _00409_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f2 sky130_fd_sc_hd__dfxtp_2
XFILLER_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20556_ _07695_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__buf_4
XFILLER_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20487_ _03383_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and3_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20171__198 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__inv_2
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21108_ net198 _00877_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13930_ _06603_ _06612_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__xnor2_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21039_ clknet_leaf_2_i_clk _00808_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _06277_ _06563_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__o21bai_4
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15600_ _08243_ _08244_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__xnor2_2
X_12812_ rbzero.wall_tracer.mapY\[9\] _05404_ _05550_ vssd1 vssd1 vccd1 vccd1 _05552_
+ sky130_fd_sc_hd__o21a_1
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16580_ _09170_ _09172_ _09169_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__a21bo_1
X_13792_ _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15531_ _08148_ rbzero.wall_tracer.stepDistY\[1\] _07990_ vssd1 vssd1 vccd1 vccd1
+ _08176_ sky130_fd_sc_hd__o21a_1
XFILLER_188_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _05459_ _05484_ _05488_ _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__and4b_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _01938_ _01948_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_91_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ _08086_ _08087_ _08105_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__nor2_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _09783_ _09784_ vssd1 vssd1 vccd1 vccd1 _09785_ sky130_fd_sc_hd__or2_1
X_14413_ _06760_ _07117_ _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__or3b_1
X_11625_ _04266_ _04403_ _04229_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o21a_1
X_18181_ _01756_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__xnor2_1
X_15393_ _07904_ rbzero.wall_tracer.stepDistY\[-9\] _05206_ vssd1 vssd1 vccd1 vccd1
+ _08038_ sky130_fd_sc_hd__a21o_1
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17132_ _09760_ _09761_ _09748_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__a21oi_1
X_14344_ _07020_ _07021_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__and2_1
XFILLER_168_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ rbzero.tex_r1\[11\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__and3_1
XFILLER_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _03589_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17063_ _03953_ _09283_ vssd1 vssd1 vccd1 vccd1 _09703_ sky130_fd_sc_hd__nor2_4
X_14275_ _07008_ _07011_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11487_ _04261_ _04264_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16014_ _08573_ _08575_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__xnor2_1
X_13226_ _05928_ _05901_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__nor2_1
XFILLER_174_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _03551_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13157_ _05743_ _05826_ _05893_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__and3_1
XFILLER_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ rbzero.tex_r1\[34\] rbzero.tex_r1\[35\] _03505_ vssd1 vssd1 vccd1 vccd1 _03515_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20230__251 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__inv_2
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _04877_ _04878_ _04879_ _04869_ net7 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o221a_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13088_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__buf_4
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _01664_ _01666_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__nand2_1
X_19704_ rbzero.pov.spi_buffer\[27\] rbzero.pov.spi_buffer\[28\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
XFILLER_211_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12039_ _04022_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__buf_2
X_16916_ _08873_ _09540_ _09555_ _08872_ vssd1 vssd1 vccd1 vccd1 _09557_ sky130_fd_sc_hd__o22ai_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17896_ _01593_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__and2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03304_ _03304_ vssd1 vssd1 vccd1 vccd1 clknet_0__03304_ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16847_ _08054_ _09216_ vssd1 vssd1 vccd1 vccd1 _09488_ sky130_fd_sc_hd__nor2_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20148__178 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__inv_2
XFILLER_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19566_ rbzero.pov.spi_counter\[5\] _03031_ _03020_ vssd1 vssd1 vccd1 vccd1 _03035_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16778_ _05210_ rbzero.wall_tracer.stepDistX\[6\] vssd1 vssd1 vccd1 vccd1 _09420_
+ sky130_fd_sc_hd__nand2_1
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18517_ _02204_ _02214_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15729_ _08188_ _08238_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__nor2_1
XFILLER_34_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19497_ _02950_ _02951_ _02968_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_59_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18448_ _10238_ _09292_ _09991_ _01737_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__o22ai_1
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18379_ _02075_ _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__or2_1
X_20410_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__or2_1
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21390_ net311 _01159_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20313__326 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__inv_2
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20272_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__buf_1
XFILLER_150_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21657_ clknet_leaf_81_i_clk _01426_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11410_ _04147_ _04148_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or2_1
XFILLER_138_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20608_ _02721_ _03467_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__and3_1
XFILLER_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12390_ net39 _05144_ _05156_ _05153_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a211o_1
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21588_ net509 _01357_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_74 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_74/HI o_rgb[2] sky130_fd_sc_hd__conb_1
XFILLER_138_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_85 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_85/HI o_rgb[17] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_96 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_96/HI zeros[6] sky130_fd_sc_hd__conb_1
X_11341_ _04100_ _04114_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__or3_4
XFILLER_180_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20539_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03430_
+ sky130_fd_sc_hd__or2_1
XFILLER_158_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14060_ _06784_ _06796_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__xnor2_1
X_11272_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _04052_
+ sky130_fd_sc_hd__or2_1
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20288__303 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__inv_2
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _05691_ _05744_ _05682_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or3_1
XFILLER_152_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14962_ rbzero.wall_tracer.stepDistX\[-12\] _07460_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07651_ sky130_fd_sc_hd__mux2_1
X_17750_ _10189_ _01453_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701_ _09238_ _09209_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__or2b_1
X_13913_ _06632_ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17681_ _09276_ _09674_ vssd1 vssd1 vccd1 vccd1 _10246_ sky130_fd_sc_hd__nor2_1
X_14893_ _07591_ _07600_ _07603_ _04039_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__o211a_1
XFILLER_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19420_ rbzero.debug_overlay.vplaneY\[10\] vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__clkbuf_4
X_13844_ _06579_ _06580_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__and2_1
XFILLER_130_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16632_ _09268_ _09274_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19351_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__and2_1
X_13775_ _06061_ _06009_ _06510_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__o21bai_1
X_16563_ _09089_ _09205_ _09192_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__a21boi_1
X_10987_ _03841_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18302_ _01890_ _01892_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__and2_1
XFILLER_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _05423_ _05426_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__and2b_1
X_15514_ _08158_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__buf_4
X_16494_ _08230_ rbzero.wall_tracer.stepDistY\[7\] _08235_ _09137_ vssd1 vssd1 vccd1
+ vccd1 _09138_ sky130_fd_sc_hd__a22oi_4
X_19282_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_leak\[3\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XFILLER_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18233_ _09661_ _09480_ _09484_ _01462_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__o22ai_1
X_15445_ _08089_ rbzero.debug_overlay.playerY\[-1\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _08090_ sky130_fd_sc_hd__mux2_1
XFILLER_175_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12657_ _05405_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ rbzero.tex_r1\[54\] _04273_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__and2_1
XFILLER_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15376_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__or2_1
X_18164_ _01863_ _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__and2_1
XFILLER_128_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12588_ _05332_ _05341_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and2_1
X_14327_ _06680_ _06739_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__or2_1
X_17115_ _09752_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11539_ gpout0.hpos\[0\] _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__nand2_1
XFILLER_129_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18095_ _01793_ _01794_ _01795_ _09863_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__a31o_1
XFILLER_128_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17046_ _08237_ _09279_ _08283_ vssd1 vssd1 vccd1 vccd1 _09686_ sky130_fd_sc_hd__a21oi_2
X_14258_ _06882_ _06883_ _06994_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__nor3_4
XFILLER_171_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13209_ _05852_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a21oi_4
X_14189_ _05984_ _06671_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__nor2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _02629_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__clkbuf_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _01647_ _01648_ _01649_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a21o_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20403__28 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17879_ _07974_ _09164_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__or2_1
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20890_ clknet_leaf_83_i_clk _00659_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19549_ rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\] _03019_ vssd1 vssd1
+ vccd1 vccd1 _03022_ sky130_fd_sc_hd__and3_1
XFILLER_59_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19572__29 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
XFILLER_179_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21511_ net432 _01280_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21442_ net363 _01211_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21373_ net294 _01142_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _03801_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _04666_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkinv_4
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10841_ _03765_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _06293_ _06296_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nand2_1
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10772_ _03717_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__clkbuf_4
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12511_ _05263_ rbzero.wall_tracer.trackDistY\[-4\] _05265_ vssd1 vssd1 vccd1 vccd1
+ _05266_ sky130_fd_sc_hd__a21o_1
X_13491_ _06173_ _06186_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__nor2_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15230_ _07879_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__inv_2
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _05199_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15161_ _07785_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _07816_
+ sky130_fd_sc_hd__nand2_1
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ net34 net64 _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__nor3b_1
XFILLER_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14112_ _06681_ _06688_ _06693_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ rbzero.texV\[7\] _04058_ _04057_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a21boi_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15092_ _07750_ _07751_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__and2_1
XFILLER_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _06777_ _06778_ _06779_ _06773_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__a22o_1
XFILLER_181_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18920_ rbzero.spi_registers.spi_counter\[4\] _02583_ vssd1 vssd1 vccd1 vccd1 _02586_
+ sky130_fd_sc_hd__nand2_1
XFILLER_158_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11255_ _04020_ _04026_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__and2_1
XFILLER_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18851_ _02524_ _02525_ _02526_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a21oi_1
X_11186_ rbzero.map_rom.f2 _03933_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__or2_1
XFILLER_171_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17802_ _09674_ _09417_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__nor2_1
XFILLER_94_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18782_ _02457_ _02459_ _02458_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a21boi_1
X_15994_ _08589_ _08598_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17733_ _09812_ _10297_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__nand2_1
X_14945_ _07621_ _07638_ _07639_ _07620_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__o211a_1
XFILLER_48_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17664_ _10225_ _10227_ vssd1 vssd1 vccd1 vccd1 _10229_ sky130_fd_sc_hd__and2_1
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ rbzero.wall_tracer.stepDistY\[11\] _07589_ _05188_ vssd1 vssd1 vccd1 vccd1
+ _07590_ sky130_fd_sc_hd__mux2_1
XFILLER_91_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20342__352 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__inv_2
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19403_ _02883_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__or2_1
X_16615_ _07932_ _09103_ _09100_ _09257_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__o31a_1
X_13827_ _06232_ _06275_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__and2_1
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17595_ _10015_ _10017_ vssd1 vssd1 vccd1 vccd1 _10161_ sky130_fd_sc_hd__or2b_1
XFILLER_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19334_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__nand2_1
X_13758_ _06490_ _06493_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__o21ai_1
X_16546_ _09050_ _09052_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__nor2_1
XFILLER_91_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12709_ _05444_ _05443_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__or2b_1
X_19265_ _02786_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13689_ _06379_ _06421_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__xnor2_2
X_16477_ _08963_ _09119_ _09120_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__a21bo_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18216_ _01900_ _01804_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__or2b_1
XFILLER_129_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15428_ rbzero.wall_tracer.visualWallDist\[-3\] _04013_ _05206_ vssd1 vssd1 vccd1
+ vccd1 _08073_ sky130_fd_sc_hd__a21oi_1
X_19196_ _02744_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18147_ _01839_ _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__xnor2_1
X_15359_ _07905_ _08003_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__and2_1
XFILLER_176_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18078_ _01777_ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__xor2_1
XFILLER_132_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17029_ _08178_ _09668_ vssd1 vssd1 vccd1 vccd1 _09669_ sky130_fd_sc_hd__nor2_2
X_20040_ _04990_ _03275_ _03279_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__o21a_1
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20942_ clknet_leaf_67_i_clk _00711_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20873_ clknet_leaf_62_i_clk _00642_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21425_ net346 _01194_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21356_ net277 _01125_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21287_ clknet_leaf_42_i_clk _01056_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[5\] sky130_fd_sc_hd__dfxtp_4
XFILLER_150_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11040_ _03869_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20238_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__buf_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _05609_ _05641_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__xnor2_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _04342_ vssd1 vssd1 vccd1 vccd1 _04718_
+ sky130_fd_sc_hd__mux2_1
X_14730_ rbzero.wall_tracer.stepDistY\[-11\] _07465_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07466_ sky130_fd_sc_hd__mux2_1
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20394__19 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14661_ _05741_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__or2_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ rbzero.tex_g1\[23\] rbzero.tex_g1\[22\] _04211_ vssd1 vssd1 vccd1 vccd1 _04650_
+ sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _06348_ _06326_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__xnor2_1
X_16400_ _08367_ _09026_ _09044_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__a21o_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10824_ _03756_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _07213_ _07328_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__nor2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17380_ _09939_ _09946_ vssd1 vssd1 vccd1 vccd1 _09947_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13543_ _06135_ _06133_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nor2_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16331_ _08974_ _08975_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__xnor2_2
X_10755_ _03720_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19050_ rbzero.pov.spi_buffer\[56\] rbzero.pov.ready_buffer\[56\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
X_16262_ _08905_ _08906_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__and2b_1
X_13474_ _06157_ _06166_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a21bo_1
XFILLER_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10686_ rbzero.tex_g1\[14\] rbzero.tex_g1\[15\] _03680_ vssd1 vssd1 vccd1 vccd1 _03684_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _07843_ _07845_ _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__a21oi_1
X_18001_ _01701_ _01702_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__or2_1
X_12425_ _04032_ _03914_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor2_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16193_ _08284_ _08579_ _08727_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__o21a_1
XFILLER_138_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144_ _07742_ rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 _07800_
+ sky130_fd_sc_hd__nor2_1
X_12356_ net124 _05082_ _05087_ net29 net28 vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__a2111oi_2
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] _04086_ vssd1 vssd1 vccd1 vccd1
+ _04087_ sky130_fd_sc_hd__o21ai_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15075_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__or2_1
X_19952_ rbzero.pov.ready_buffer\[33\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-9\]
+ _03209_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__o221a_1
X_12287_ net38 _05043_ _05044_ net48 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a22o_1
XFILLER_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14026_ _05855_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__nand3_2
X_18903_ _02558_ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__nand2_1
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11238_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__buf_2
XFILLER_136_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19883_ rbzero.pov.ready_buffer\[73\] _03164_ _03155_ _03190_ vssd1 vssd1 vccd1 vccd1
+ _03191_ sky130_fd_sc_hd__o211a_1
XFILLER_171_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18834_ _02503_ _02505_ _02504_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__o21bai_1
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11169_ rbzero.othery\[3\] vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__inv_2
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18765_ _02450_ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__or2b_1
XFILLER_110_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15977_ _08601_ _08602_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__xnor2_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17716_ _10233_ _10280_ vssd1 vssd1 vccd1 vccd1 _10281_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14928_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.trackDistX\[1\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__mux2_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18696_ rbzero.wall_tracer.trackDistX\[11\] rbzero.wall_tracer.stepDistX\[11\] vssd1
+ vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__xor2_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17647_ _10209_ _10210_ vssd1 vssd1 vccd1 vccd1 _10212_ sky130_fd_sc_hd__and2_1
X_14859_ _07576_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17578_ _10127_ _10143_ vssd1 vssd1 vccd1 vccd1 _10144_ sky130_fd_sc_hd__nand2_1
XFILLER_51_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19317_ rbzero.spi_registers.new_vshift\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XFILLER_32_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16529_ _09171_ _09172_ vssd1 vssd1 vccd1 vccd1 _09173_ sky130_fd_sc_hd__xor2_1
XFILLER_176_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19248_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_sky\[2\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
XFILLER_192_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19179_ rbzero.floor_leak\[0\] _02732_ _02734_ _02722_ vssd1 vssd1 vccd1 vccd1 _00740_
+ sky130_fd_sc_hd__o211a_1
X_21210_ clknet_leaf_18_i_clk _00979_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21141_ clknet_leaf_60_i_clk _00910_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21072_ net162 _00841_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20023_ _04992_ _04037_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__nand2_1
XFILLER_150_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ clknet_leaf_13_i_clk _00694_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20856_ clknet_leaf_53_i_clk _00625_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20787_ clknet_leaf_16_i_clk _00556_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10540_ rbzero.tex_r0\[20\] rbzero.tex_r0\[19\] _03602_ vssd1 vssd1 vccd1 vccd1 _03607_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _03569_ vssd1 vssd1 vccd1 vccd1 _03571_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12210_ _04961_ _04960_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and2b_1
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21408_ net329 _01177_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13190_ _05814_ _05821_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _04909_ net62 _04911_ net12 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__o211a_1
XFILLER_194_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21339_ net260 _01108_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ _04840_ _04325_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nor2_1
XFILLER_81_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11023_ _03860_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__clkbuf_1
X_15900_ _08511_ _08543_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__nor2_1
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16880_ _08282_ _07994_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09521_ sky130_fd_sc_hd__or4_1
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _07995_ _07989_ _08475_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__or3_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _02144_ _02246_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__xnor2_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _08403_ _08404_ _08405_ vssd1 vssd1 vccd1 vccd1 _08407_ sky130_fd_sc_hd__nand3_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _05586_ _05587_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _10057_ _10066_ vssd1 vssd1 vccd1 vccd1 _10067_ sky130_fd_sc_hd__nand2_1
XFILLER_73_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14713_ _05779_ _07362_ _07372_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__o21ai_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _04263_ vssd1 vssd1 vccd1 vccd1 _04701_
+ sky130_fd_sc_hd__mux2_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _02176_ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__or2_1
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _07938_ _07939_ _08109_ vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__or3_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _08747_ _09699_ _08250_ vssd1 vssd1 vccd1 vccd1 _09999_ sky130_fd_sc_hd__o21ai_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _07350_ _07360_ _05793_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__mux2_1
X_11856_ rbzero.tex_g1\[9\] rbzero.tex_g1\[8\] _04350_ vssd1 vssd1 vccd1 vccd1 _04633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10807_ _03747_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14575_ _07305_ _07095_ _07096_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__and3_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17363_ _09368_ _09217_ vssd1 vssd1 vccd1 vccd1 _09930_ sky130_fd_sc_hd__nor2_1
X_11787_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _04262_ vssd1 vssd1 vccd1 vccd1 _04565_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19102_ _02684_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__clkbuf_1
X_16314_ _08290_ _08291_ _08958_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__a21bo_1
XFILLER_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13526_ _06256_ _06257_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10738_ rbzero.tex_g0\[54\] rbzero.tex_g0\[53\] _03706_ vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__mux2_1
X_17294_ _09854_ _09856_ _09855_ vssd1 vssd1 vccd1 vccd1 _09866_ sky130_fd_sc_hd__o21bai_1
XFILLER_186_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19033_ rbzero.pov.spi_buffer\[48\] rbzero.pov.ready_buffer\[48\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
X_13457_ _06152_ _06188_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or2b_1
X_16245_ _08881_ _08882_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__nor2_1
X_10669_ rbzero.tex_g1\[22\] rbzero.tex_g1\[23\] _03669_ vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__mux2_1
X_12408_ _05141_ _05172_ _05174_ net35 vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__o211a_1
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ _06046_ _06123_ _06122_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a21bo_1
X_16176_ _08674_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12339_ net27 net26 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__and2b_1
X_15127_ _07758_ _07769_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__nand2_1
XFILLER_173_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15058_ rbzero.debug_overlay.vplaneX\[-6\] _07708_ vssd1 vssd1 vccd1 vccd1 _07720_
+ sky130_fd_sc_hd__xor2_1
X_19935_ rbzero.debug_overlay.playerY\[3\] _03193_ _03229_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _01001_ sky130_fd_sc_hd__a211o_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _06240_ _06707_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__nor2_1
X_19866_ rbzero.debug_overlay.playerX\[1\] _03167_ rbzero.debug_overlay.playerX\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18817_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nand2_1
XFILLER_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19599__54 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
XFILLER_56_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19797_ _03127_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18748_ _02428_ _02430_ _02429_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a21boi_1
XFILLER_37_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03297_ clknet_0__03297_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03297_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18679_ _02364_ _02374_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20710_ clknet_leaf_16_i_clk _00001_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20641_ clknet_leaf_26_i_clk _00425_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20572_ _02721_ _03445_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__and3_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21124_ clknet_leaf_65_i_clk _00893_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21055_ clknet_leaf_57_i_clk _00824_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20006_ rbzero.pov.ready_buffer\[10\] _03239_ _03242_ _02906_ _02730_ vssd1 vssd1
+ vccd1 vccd1 _01047_ sky130_fd_sc_hd__o221a_1
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ gpout0.vpos\[4\] gpout0.vpos\[3\] _04488_ gpout0.vpos\[5\] vssd1 vssd1 vccd1
+ vccd1 _04489_ sky130_fd_sc_hd__or4b_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ clknet_leaf_64_i_clk _00677_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _05435_ _05436_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or3b_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _04004_ _04419_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__and3b_1
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20839_ clknet_leaf_26_i_clk _00608_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14360_ _06882_ _07034_ _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11572_ rbzero.tex_r1\[2\] _04350_ _04217_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a21o_1
XFILLER_156_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _06044_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__xor2_1
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10523_ rbzero.tex_r0\[28\] rbzero.tex_r0\[27\] _03591_ vssd1 vssd1 vccd1 vccd1 _03598_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 i_gpout2_sel[5] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_8
XFILLER_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14291_ _06798_ _06816_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__or2b_1
XFILLER_202_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13242_ _05856_ _05877_ _05888_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a21oi_1
X_16030_ _07980_ _08674_ _08020_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__or3_1
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10454_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _03558_ vssd1 vssd1 vccd1 vccd1 _03562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__inv_2
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10385_ _03523_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
X_12124_ net52 _04853_ _04857_ net50 _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a221o_1
XFILLER_112_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17981_ _01677_ _01683_ rbzero.wall_tracer.trackDistX\[4\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00593_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19720_ _03087_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
X_12055_ _04820_ _04823_ _04825_ _04827_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__o32a_1
X_16932_ _09425_ _09438_ _09572_ vssd1 vssd1 vccd1 vccd1 _09573_ sky130_fd_sc_hd__a21o_1
XFILLER_81_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03320_ _03320_ vssd1 vssd1 vccd1 vccd1 clknet_0__03320_ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11006_ _03851_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__clkbuf_1
X_19651_ _03051_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16863_ _09502_ _09503_ vssd1 vssd1 vccd1 vccd1 _09504_ sky130_fd_sc_hd__and2b_1
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18602_ _02293_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__xor2_1
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15814_ _08456_ _08457_ _08458_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__a21oi_1
X_19582_ clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__buf_1
XFILLER_65_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16794_ _09428_ _09435_ vssd1 vssd1 vccd1 vccd1 _09436_ sky130_fd_sc_hd__xnor2_2
XFILLER_46_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18533_ _02132_ _02134_ _02133_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__o21bai_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _08382_ _08388_ _08389_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__a21o_1
X_12957_ _05691_ _05673_ _05683_ _05693_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__or4_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20060__98 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__inv_2
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _04271_ vssd1 vssd1 vccd1 vccd1 _04684_
+ sky130_fd_sc_hd__mux2_1
X_18464_ _02033_ _02055_ _02031_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a21oi_1
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15676_ _08287_ _08285_ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__nand2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12888_ rbzero.wall_tracer.visualWallDist\[2\] _05571_ _04001_ vssd1 vssd1 vccd1
+ vccd1 _05625_ sky130_fd_sc_hd__a21oi_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _09686_ _09980_ _09981_ vssd1 vssd1 vccd1 vccd1 _09982_ sky130_fd_sc_hd__a21o_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _07309_ _07310_ _07312_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18395_ _01859_ _01863_ _01958_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11839_ rbzero.tex_g1\[47\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04616_
+ sky130_fd_sc_hd__a31o_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17346_ _09633_ _09636_ _09911_ vssd1 vssd1 vccd1 vccd1 _09913_ sky130_fd_sc_hd__and3_1
X_14558_ _07286_ _07292_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _05983_ _06245_ _06243_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _05531_ _09076_ vssd1 vssd1 vccd1 vccd1 _09851_ sky130_fd_sc_hd__nand2_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14489_ _07172_ _07221_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__a21oi_1
X_19016_ _02639_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__clkbuf_1
X_16228_ _08180_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16159_ _08766_ _08800_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19918_ rbzero.debug_overlay.playerY\[0\] _08030_ vssd1 vssd1 vccd1 vccd1 _03216_
+ sky130_fd_sc_hd__or2_1
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19849_ _03139_ _03162_ _03163_ _03157_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__o211a_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20125__157 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__inv_2
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20624_ clknet_leaf_52_i_clk _00408_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f3 sky130_fd_sc_hd__dfxtp_2
XFILLER_71_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20555_ rbzero.traced_texVinit\[0\] _09770_ _09771_ _09068_ vssd1 vssd1 vccd1 vccd1
+ _01408_ sky130_fd_sc_hd__a22o_1
XFILLER_138_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20486_ _03383_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__a21o_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21107_ net197 _00876_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21038_ clknet_leaf_2_i_clk _00807_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13860_ _06595_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__nand2_1
X_19578__35 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _05548_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__o21bai_1
X_13791_ _05824_ _06031_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nor2_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _05194_ _08172_ _08174_ _08002_ vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__a211o_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _05445_ _05489_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__xnor2_2
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15461_ _08086_ _08087_ _08105_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__and3_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _05419_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__and2b_1
XFILLER_203_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ rbzero.wall_tracer.mapX\[7\] _05525_ vssd1 vssd1 vccd1 vccd1 _09784_ sky130_fd_sc_hd__nor2_1
X_14412_ _06696_ _06698_ _07072_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__a21oi_1
X_11624_ rbzero.tex_r1\[35\] rbzero.tex_r1\[34\] _04350_ vssd1 vssd1 vccd1 vccd1 _04403_
+ sky130_fd_sc_hd__mux2_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18180_ _01879_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__xor2_1
X_15392_ _07502_ _08036_ _07933_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__mux2_2
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ _03477_ _04446_ vssd1 vssd1 vccd1 vccd1 _09761_ sky130_fd_sc_hd__nand2_1
X_11555_ rbzero.tex_r1\[9\] rbzero.tex_r1\[8\] _04291_ vssd1 vssd1 vccd1 vccd1 _04334_
+ sky130_fd_sc_hd__mux2_1
X_14343_ _07070_ _07079_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ rbzero.tex_r0\[36\] rbzero.tex_r0\[35\] _03580_ vssd1 vssd1 vccd1 vccd1 _03589_
+ sky130_fd_sc_hd__mux2_1
X_14274_ _07009_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__xnor2_1
X_17062_ _09694_ _09701_ vssd1 vssd1 vccd1 vccd1 _09702_ sky130_fd_sc_hd__xor2_2
X_11486_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__buf_6
XFILLER_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13225_ _05945_ _05949_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21oi_2
XFILLER_171_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16013_ _08656_ _08657_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__xor2_2
XFILLER_137_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10437_ rbzero.tex_r1\[2\] rbzero.tex_r1\[3\] _03549_ vssd1 vssd1 vccd1 vccd1 _03551_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13156_ _05801_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__clkbuf_4
X_10368_ _03514_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ net3 net4 net5 vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21oi_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__buf_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _01664_ _01666_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__or2_2
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10299_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__buf_2
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19703_ _03078_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12038_ _04809_ _04810_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__o21ba_1
X_16915_ _08873_ _09555_ _09421_ vssd1 vssd1 vccd1 vccd1 _09556_ sky130_fd_sc_hd__or3b_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17895_ _01596_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03303_ _03303_ vssd1 vssd1 vccd1 vccd1 clknet_0__03303_ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16846_ _09485_ _09486_ vssd1 vssd1 vccd1 vccd1 _09487_ sky130_fd_sc_hd__nand2_1
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19565_ rbzero.pov.spi_counter\[5\] _03031_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__and2_1
XFILLER_81_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ _08237_ _09279_ _08180_ vssd1 vssd1 vccd1 vccd1 _09419_ sky130_fd_sc_hd__a21o_1
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__inv_2
XFILLER_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18516_ _02109_ _02213_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__xor2_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _08306_ _08310_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19496_ _02973_ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nand2_1
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18447_ _01737_ _10238_ _09292_ _09991_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__or4_1
X_15659_ _08255_ _08303_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__nand2_1
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18378_ _01474_ _09215_ _01941_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__o31a_1
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ _09896_ vssd1 vssd1 vccd1 vccd1 _09897_ sky130_fd_sc_hd__inv_2
XFILLER_105_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20271_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__buf_1
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21656_ clknet_leaf_84_i_clk _01425_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20607_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__or2_1
XFILLER_165_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21587_ net508 _01356_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_75 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_75/HI o_rgb[3] sky130_fd_sc_hd__conb_1
XFILLER_71_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_86 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_86/HI o_rgb[18] sky130_fd_sc_hd__conb_1
XFILLER_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11340_ _04099_ _04069_ _04097_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__nor3_2
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20538_ rbzero.texV\[8\] _03327_ _03332_ _03429_ vssd1 vssd1 vccd1 vccd1 _01404_
+ sky130_fd_sc_hd__a22o_1
Xtop_ew_algofoogle_97 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_97/HI zeros[7] sky130_fd_sc_hd__conb_1
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ _04049_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nand2_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20469_ _03272_ _03370_ _03371_ _03250_ rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1
+ _01393_ sky130_fd_sc_hd__a32o_1
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _05690_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__inv_2
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14961_ _05201_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__buf_4
XFILLER_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16700_ _09324_ _09326_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__or2_2
XFILLER_102_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13912_ _06576_ _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nand2_1
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17680_ _10099_ _10244_ vssd1 vssd1 vccd1 vccd1 _10245_ sky130_fd_sc_hd__xnor2_1
X_14892_ _07602_ _04019_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__nand2_1
XFILLER_207_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16631_ _09269_ _09273_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__xnor2_1
X_13843_ _06259_ _06575_ _06578_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__or3_1
XFILLER_74_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19350_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__nor2_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20108__141 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__inv_2
X_16562_ _09059_ _08470_ _08546_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__or3_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13774_ _05944_ _06009_ _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__or3b_1
X_10986_ net48 rbzero.tex_b0\[63\] _03762_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__mux2_1
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18301_ _01966_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15513_ _05208_ _08157_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__or2_2
XFILLER_204_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12725_ _05424_ _05425_ _05427_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__o21a_1
X_19281_ _02795_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__clkbuf_1
X_16493_ _08981_ _07574_ _08234_ _09136_ _07970_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__a311o_1
XFILLER_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18232_ _01930_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__nand2_1
XFILLER_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15444_ _08030_ _08088_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__and2_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ _05388_ _05398_ _05399_ _05397_ rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1
+ vccd1 _05406_ sky130_fd_sc_hd__a32o_1
XFILLER_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _04384_ _04385_ _04226_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_1
X_18163_ _01739_ _01620_ _01862_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__o21ai_1
X_15375_ _05197_ rbzero.wall_tracer.stepDistX\[-7\] vssd1 vssd1 vccd1 vccd1 _08020_
+ sky130_fd_sc_hd__nor2_2
X_12587_ _05323_ _05288_ _05319_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__or3_1
XFILLER_184_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ _04821_ _09750_ _09751_ vssd1 vssd1 vccd1 vccd1 _09752_ sky130_fd_sc_hd__and3_1
XFILLER_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14326_ _06240_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__and3b_1
XFILLER_129_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _04317_ _04163_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__and2_1
X_18094_ _01793_ _01794_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17045_ _09141_ _09420_ _08194_ vssd1 vssd1 vccd1 vccd1 _09685_ sky130_fd_sc_hd__a21o_1
X_14257_ _06884_ _06915_ _06917_ _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__or4_2
X_11469_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _04213_ vssd1 vssd1 vccd1 vccd1 _04249_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13208_ _05856_ _05877_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a21o_2
XFILLER_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20154__183 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__inv_2
X_14188_ _06769_ _06671_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__nor2_1
XFILLER_140_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _05865_ _05870_ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__or3b_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ rbzero.pov.spi_buffer\[30\] rbzero.pov.ready_buffer\[30\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XFILLER_140_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _01647_ _01648_ _01649_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__and3_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17878_ _09661_ _09029_ _09165_ _01462_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__o22ai_1
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16829_ _09461_ _09465_ vssd1 vssd1 vccd1 vccd1 _09470_ sky130_fd_sc_hd__or2_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19548_ rbzero.pov.spi_counter\[0\] _03019_ _03021_ vssd1 vssd1 vccd1 vccd1 _00822_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_59_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ _02941_ _02944_ _02957_ _02959_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__o31a_1
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21510_ net431 _01279_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21441_ net362 _01210_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21372_ net293 _01141_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[15\] sky130_fd_sc_hd__dfxtp_1
X_20237__258 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__inv_2
XFILLER_190_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ rbzero.tex_g0\[6\] rbzero.tex_g0\[5\] _03762_ vssd1 vssd1 vccd1 vccd1 _03765_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ _03728_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12510_ rbzero.wall_tracer.trackDistY\[3\] _05264_ rbzero.wall_tracer.trackDistY\[-5\]
+ _05236_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
X_13490_ _06225_ _06226_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and2_1
XFILLER_198_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12441_ net71 rbzero.wall_tracer.state\[5\] _05190_ vssd1 vssd1 vccd1 vccd1 _05199_
+ sky130_fd_sc_hd__and3_1
XFILLER_139_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21639_ clknet_leaf_19_i_clk _01408_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12372_ net33 net32 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__nor2_2
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15160_ _07803_ _07808_ _07813_ _07676_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__o31ai_1
Xclkbuf_leaf_43_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14111_ _06843_ _06844_ _06846_ _06847_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__a22o_1
XFILLER_138_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11323_ rbzero.texV\[8\] _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__xor2_1
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15091_ _07736_ _07748_ _07749_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__or3_1
XFILLER_126_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ _06002_ _06758_ _06759_ _06770_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a31o_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11254_ _04031_ _04032_ _04002_ _04035_ _00000_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a41o_1
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18850_ _02517_ _02519_ _02518_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__o21bai_1
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11185_ rbzero.map_rom.f2 _03933_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__nand2_1
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17801_ _10244_ _01503_ _01504_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__a21o_1
XFILLER_122_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18781_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__and2_1
X_15993_ _08629_ _08637_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17732_ _10295_ _10296_ vssd1 vssd1 vccd1 vccd1 _10297_ sky130_fd_sc_hd__and2b_4
XFILLER_208_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14944_ rbzero.wall_tracer.visualWallDist\[6\] _07618_ vssd1 vssd1 vccd1 vccd1 _07639_
+ sky130_fd_sc_hd__or2_1
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17663_ _10225_ _10227_ vssd1 vssd1 vccd1 vccd1 _10228_ sky130_fd_sc_hd__nor2_1
X_14875_ _05737_ _05736_ _07588_ _07468_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__nor4_4
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19402_ _02886_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__and2_1
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16614_ _09009_ _09099_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__nand2_1
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13826_ _06335_ _06560_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a21oi_2
X_17594_ _10048_ _10159_ vssd1 vssd1 vccd1 vccd1 _10160_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19333_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__nor2_1
XFILLER_204_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16545_ _09055_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__inv_2
X_13757_ _06438_ _06455_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__xor2_1
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _03832_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19264_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_floor\[2\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
X_12708_ _05447_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__xor2_4
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16476_ _08283_ _08177_ _08264_ _08626_ vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__a2bb2o_1
X_13688_ _06376_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__or2b_1
X_18215_ _01897_ _01899_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__or2_1
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15427_ _07904_ _08071_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__nand2_1
X_19195_ _09753_ _02743_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__and2_1
X_12639_ _05388_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__nand2_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ _01840_ _01846_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__o21ai_1
XFILLER_106_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14309_ _06696_ _06667_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__nor2_1
X_18077_ _01611_ _01655_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15289_ _05349_ _05469_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17028_ _08570_ vssd1 vssd1 vccd1 vccd1 _09668_ sky130_fd_sc_hd__buf_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ rbzero.pov.spi_buffer\[22\] rbzero.pov.ready_buffer\[22\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20941_ clknet_leaf_67_i_clk _00710_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_96_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20872_ clknet_leaf_63_i_clk _00641_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21424_ net345 _01193_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21355_ net276 _01124_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21286_ clknet_leaf_31_i_clk _01055_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[4\] sky130_fd_sc_hd__dfxtp_4
XFILLER_150_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _05724_ _05683_ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__o21ba_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _04342_ vssd1 vssd1 vccd1 vccd1 _04717_
+ sky130_fd_sc_hd__mux2_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14660_ _07371_ _07396_ _05779_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__mux2_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11872_ rbzero.tex_g1\[21\] rbzero.tex_g1\[20\] _04336_ vssd1 vssd1 vccd1 vccd1 _04649_
+ sky130_fd_sc_hd__mux2_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _06304_ _06323_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__xnor2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10823_ rbzero.tex_g0\[14\] rbzero.tex_g0\[13\] _03751_ vssd1 vssd1 vccd1 vccd1 _03756_
+ sky130_fd_sc_hd__mux2_1
X_14591_ _07326_ _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__xnor2_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16330_ _08178_ _08194_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__nor2_1
X_13542_ _06150_ _06192_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__xnor2_2
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _03718_ vssd1 vssd1 vccd1 vccd1 _03720_
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16261_ _08902_ _08904_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__nand2_1
X_13473_ _06165_ _06158_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__or2b_1
X_10685_ _03683_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18000_ _09526_ _01576_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15212_ _07820_ rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1 vccd1 _07864_
+ sky130_fd_sc_hd__xnor2_1
X_12424_ _05188_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__buf_2
XFILLER_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16192_ _08828_ _08829_ _08831_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__or3b_1
XFILLER_126_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20372__379 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__inv_2
X_15143_ _07797_ _07798_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__xnor2_1
X_12355_ _05117_ _05119_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and3_1
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11306_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] rbzero.texV\[1\] rbzero.traced_texVinit\[1\]
+ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a221o_1
X_12286_ net23 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__inv_2
X_15074_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\]
+ rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__or4b_1
X_19951_ _03242_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__buf_2
XFILLER_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14025_ _06704_ _06760_ _06761_ _05825_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__o22ai_2
X_11237_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__buf_4
X_18902_ _02559_ rbzero.spi_registers.spi_counter\[0\] _02566_ _02568_ _02571_ vssd1
+ vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o2111a_1
XFILLER_171_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19882_ _03188_ _03185_ _02822_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a21o_1
XFILLER_136_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18833_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nand2_1
X_11168_ rbzero.otherx\[0\] _03919_ _03935_ rbzero.othery\[4\] _03956_ vssd1 vssd1
+ vccd1 vccd1 _03957_ sky130_fd_sc_hd__a221o_1
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18764_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nand2_1
XFILLER_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15976_ _08605_ _08606_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__xnor2_2
X_11099_ _03900_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20266__284 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__inv_2
X_17715_ _10277_ _10279_ vssd1 vssd1 vccd1 vccd1 _10280_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14927_ _07621_ _07626_ _07627_ _07620_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__o211a_1
XFILLER_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18695_ _02319_ _02320_ _02318_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__o21ai_1
XFILLER_64_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ _10209_ _10210_ vssd1 vssd1 vccd1 vccd1 _10211_ sky130_fd_sc_hd__nor2_1
X_14858_ rbzero.wall_tracer.stepDistY\[7\] _07575_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07576_ sky130_fd_sc_hd__mux2_1
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _06500_ _06493_ _06544_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__or4b_1
XFILLER_189_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17577_ _10140_ _10141_ _10137_ vssd1 vssd1 vccd1 vccd1 _10143_ sky130_fd_sc_hd__a21o_1
X_14789_ _05800_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__nand2_1
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19316_ _02814_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16528_ _08054_ _08425_ vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__nor2_1
XFILLER_32_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19247_ _02776_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__clkbuf_1
X_16459_ _08097_ vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__buf_4
XFILLER_118_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19178_ rbzero.spi_registers.new_leak\[0\] _02733_ vssd1 vssd1 vccd1 vccd1 _02734_
+ sky130_fd_sc_hd__or2_1
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18129_ _07974_ _09217_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__or2_1
XFILLER_191_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21140_ clknet_leaf_60_i_clk _00909_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21071_ net161 _00840_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20022_ _04021_ _04026_ _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__and3_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20924_ clknet_leaf_76_i_clk _00693_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ clknet_leaf_4_i_clk _00624_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20786_ clknet_leaf_21_i_clk _00555_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10470_ _03570_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21407_ net328 _01176_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _04910_ net61 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__or2_1
XFILLER_136_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21338_ net259 _01107_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ net6 _04841_ _04842_ net5 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a31o_1
X_21269_ clknet_leaf_65_i_clk _01038_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _03854_ vssd1 vssd1 vccd1 vccd1 _03860_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _07980_ _07929_ _07930_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__or3_1
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _08403_ _08404_ _08405_ vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__a21o_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ _05582_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__xor2_4
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17500_ _10064_ _10065_ vssd1 vssd1 vccd1 vccd1 _10066_ sky130_fd_sc_hd__and2_1
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _05963_ _07445_ _07446_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__o31a_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11924_ _04140_ _04683_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__or3_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _10094_ _09215_ _02072_ _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__o31a_1
XFILLER_206_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _08334_ _08336_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__xnor2_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _08377_ _08519_ _09699_ vssd1 vssd1 vccd1 vccd1 _09998_ sky130_fd_sc_hd__a21o_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _07378_ _07335_ _07336_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__or3b_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11855_ _04629_ _04630_ _04631_ _04379_ _04209_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__o221a_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10806_ rbzero.tex_g0\[22\] rbzero.tex_g0\[21\] _03740_ vssd1 vssd1 vccd1 vccd1 _03747_
+ sky130_fd_sc_hd__mux2_1
X_17362_ _09927_ _09928_ vssd1 vssd1 vccd1 vccd1 _09929_ sky130_fd_sc_hd__nand2_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14574_ _07309_ _07310_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nand2_1
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _04306_ _04559_ _04563_ _04371_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a211o_1
X_19101_ rbzero.spi_registers.spi_buffer\[6\] rbzero.spi_registers.spi_buffer\[5\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XFILLER_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16313_ _08292_ _07996_ _07959_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__or3_1
X_13525_ _06258_ _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17293_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09865_ sky130_fd_sc_hd__nand2_1
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10737_ _03710_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__clkbuf_1
X_19032_ _02647_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
X_16244_ _08827_ _08833_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__xnor2_1
X_13456_ _06150_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__and2b_1
X_10668_ _03674_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _05145_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or2_1
XFILLER_51_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ _08818_ _08819_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__or2_1
X_13387_ _06122_ _06046_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand3b_1
X_10599_ rbzero.tex_g1\[55\] rbzero.tex_g1\[56\] _03635_ vssd1 vssd1 vccd1 vccd1 _03638_
+ sky130_fd_sc_hd__mux2_1
XFILLER_115_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15126_ _07761_ _07771_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__nor2_1
X_12338_ net48 net39 net38 net40 _05082_ _05087_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__mux4_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15057_ _07719_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__clkbuf_1
X_19934_ rbzero.pov.ready_buffer\[56\] _03146_ _03227_ _03228_ _03197_ vssd1 vssd1
+ vccd1 vccd1 _03229_ sky130_fd_sc_hd__o221a_1
X_12269_ _04989_ _04990_ _05021_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_141_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14008_ _06245_ _06668_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__nor2_1
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19865_ rbzero.debug_overlay.playerX\[2\] rbzero.debug_overlay.playerX\[1\] _03167_
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or3_1
XFILLER_110_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18816_ _02496_ _01438_ rbzero.wall_tracer.trackDistY\[2\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00615_ sky130_fd_sc_hd__o2bb2a_1
X_19796_ rbzero.pov.spi_buffer\[71\] rbzero.pov.spi_buffer\[72\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15959_ _08601_ _08602_ _08603_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__a21oi_2
X_18747_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__and2_1
XFILLER_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03296_ clknet_0__03296_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03296_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18678_ _02367_ _02373_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17629_ _10192_ _10193_ vssd1 vssd1 vccd1 vccd1 _10194_ sky130_fd_sc_hd__nor2_1
XFILLER_211_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20640_ clknet_leaf_25_i_clk _00424_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20571_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__or2_1
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21123_ net213 _00892_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21054_ clknet_leaf_57_i_clk _00823_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20005_ rbzero.pov.ready_buffer\[9\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[0\]
+ _02730_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__o221a_1
XFILLER_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ clknet_leaf_64_i_clk _00676_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_203_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _04022_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__and2b_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ clknet_leaf_25_i_clk _00607_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20102__136 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__inv_2
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11571_ _04336_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__clkbuf_8
X_20769_ clknet_leaf_33_i_clk _00538_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _05995_ _05921_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o21ai_1
XFILLER_161_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10522_ _03597_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _07006_ _07026_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__xnor2_2
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10453_ _03561_ vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__clkbuf_1
X_13241_ _05939_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__buf_2
XFILLER_202_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10384_ rbzero.tex_r1\[27\] rbzero.tex_r1\[28\] _03516_ vssd1 vssd1 vccd1 vccd1 _03523_
+ sky130_fd_sc_hd__mux2_1
X_13172_ _05871_ _05905_ _05907_ _05908_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__o211a_2
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ net49 _04838_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__and2_1
XFILLER_123_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17980_ _01681_ _01682_ _09780_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12054_ _03473_ rbzero.row_render.wall\[0\] _04814_ vssd1 vssd1 vccd1 vccd1 _04828_
+ sky130_fd_sc_hd__and3b_1
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16931_ _09436_ _09437_ vssd1 vssd1 vccd1 vccd1 _09572_ sky130_fd_sc_hd__and2b_1
XFILLER_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11005_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _03843_ vssd1 vssd1 vccd1 vccd1 _03851_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19650_ rbzero.pov.spi_buffer\[1\] rbzero.pov.spi_buffer\[2\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
X_16862_ _09245_ _08075_ _08159_ _08150_ vssd1 vssd1 vccd1 vccd1 _09503_ sky130_fd_sc_hd__or4_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15813_ _08442_ _08455_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__nor2_1
X_18601_ _02296_ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nor2_1
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16793_ _08239_ _09434_ vssd1 vssd1 vccd1 vccd1 _09435_ sky130_fd_sc_hd__nor2_1
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18532_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__nand2_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _08375_ _08381_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__nor2_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ _05692_ _05636_ _05648_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__or3b_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11907_ _04232_ _04670_ _04674_ _04682_ _04244_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o311a_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _02141_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _08318_ _08309_ _08319_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__a21o_1
X_12887_ _05333_ _05334_ _04031_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__o21ai_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17414_ _08767_ _09552_ _09973_ _08283_ vssd1 vssd1 vccd1 vccd1 _09981_ sky130_fd_sc_hd__o22a_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14626_ _07095_ _07035_ _07099_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__a21oi_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _02084_ _02092_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__xnor2_1
X_11838_ rbzero.tex_g1\[46\] _04272_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__and2_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20378__385 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__inv_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _09633_ _09636_ _09911_ vssd1 vssd1 vccd1 vccd1 _09912_ sky130_fd_sc_hd__a21oi_2
X_14557_ _07285_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__xor2_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11769_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _04341_ vssd1 vssd1 vccd1 vccd1 _04547_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20077__113 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__inv_2
XFILLER_53_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13508_ _05940_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__clkbuf_4
XFILLER_140_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17276_ _09846_ _09847_ _09848_ vssd1 vssd1 vccd1 vccd1 _09850_ sky130_fd_sc_hd__a21oi_1
X_14488_ _07222_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__and2b_1
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19015_ rbzero.pov.spi_buffer\[39\] rbzero.pov.ready_buffer\[39\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16227_ _08170_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__clkbuf_4
X_13439_ _06080_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__clkinv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16158_ _08802_ _08579_ _08777_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__or3_1
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ rbzero.wall_tracer.rayAddendX\[1\] _07695_ _07767_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _07768_ sky130_fd_sc_hd__a22o_1
XFILLER_115_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16089_ _08726_ _08733_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__or2b_1
XFILLER_138_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19917_ rbzero.debug_overlay.playerY\[-1\] _03193_ _03215_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00997_ sky130_fd_sc_hd__a211o_1
XFILLER_64_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19848_ _08078_ _03143_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__nand2_1
XFILLER_110_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _03118_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20623_ clknet_leaf_52_i_clk _00407_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f4 sky130_fd_sc_hd__dfxtp_2
XFILLER_71_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20554_ _03441_ _03442_ rbzero.texV\[11\] net60 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_192_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20485_ _03379_ _03381_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__nand2_1
XFILLER_118_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21106_ net196 _00875_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21037_ clknet_leaf_77_i_clk _00806_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12810_ rbzero.wall_tracer.mapY\[8\] _05404_ _05547_ vssd1 vssd1 vccd1 vccd1 _05550_
+ sky130_fd_sc_hd__a21bo_1
X_13790_ _06382_ _06002_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nand2_1
XFILLER_62_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12741_ _05416_ _05442_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a31o_1
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ _08097_ _08104_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__nor2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12672_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nand2_1
XFILLER_169_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _07115_ _07119_ _07117_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__o21ba_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _04379_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__or2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15391_ _05355_ _05477_ _07893_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__mux2_1
XFILLER_129_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17130_ _03477_ _04446_ vssd1 vssd1 vccd1 vccd1 _09760_ sky130_fd_sc_hd__or2_1
X_14342_ _07077_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__xor2_1
X_11554_ _04326_ _04330_ _04331_ _04247_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__o221a_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10505_ _03588_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
X_17061_ _09696_ _09700_ vssd1 vssd1 vccd1 vccd1 _09701_ sky130_fd_sc_hd__xnor2_1
X_14273_ _06680_ _06708_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nor2_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _04126_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__buf_4
XFILLER_184_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16012_ _08578_ _08580_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_0__f__03299_ clknet_0__03299_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03299_
+ sky130_fd_sc_hd__clkbuf_16
X_13224_ _05800_ _05950_ _05955_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__o211a_2
X_10436_ _03550_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13155_ _05743_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__buf_2
XFILLER_100_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10367_ rbzero.tex_r1\[35\] rbzero.tex_r1\[36\] _03505_ vssd1 vssd1 vccd1 vccd1 _03514_
+ sky130_fd_sc_hd__mux2_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _04154_ _03477_ _04840_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__mux2_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13086_ _05800_ _05812_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__o21ai_4
X_10298_ gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__clkbuf_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ _01543_ _01545_ _01665_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__o21a_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19702_ rbzero.pov.spi_buffer\[26\] rbzero.pov.spi_buffer\[27\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
X_12037_ _04004_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__buf_2
X_16914_ _09554_ _09138_ _05198_ vssd1 vssd1 vccd1 vccd1 _09555_ sky130_fd_sc_hd__mux2_2
XFILLER_78_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17894_ _08275_ _08427_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__03302_ _03302_ vssd1 vssd1 vccd1 vccd1 clknet_0__03302_ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16845_ _08160_ _09352_ _09484_ vssd1 vssd1 vccd1 vccd1 _09486_ sky130_fd_sc_hd__or3_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19564_ _03033_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__clkbuf_1
X_16776_ _09117_ _09417_ vssd1 vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__nor2_1
XFILLER_111_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13988_ _06696_ _06677_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__nor2_1
XFILLER_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15727_ _08313_ _08324_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__xnor2_1
X_18515_ _02211_ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__nor2_1
XFILLER_74_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12939_ _05601_ _05604_ _05638_ _05649_ _05628_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__o41a_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19495_ _02904_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02974_
+ sky130_fd_sc_hd__or2_1
XFILLER_206_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18446_ _01971_ _02027_ _02036_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__o21ai_4
X_15658_ rbzero.wall_tracer.visualWallDist\[-11\] _08148_ _05198_ _08199_ vssd1 vssd1
+ vccd1 vccd1 _08303_ sky130_fd_sc_hd__and4_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ _07218_ _07323_ _07334_ _07332_ _07345_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__a311o_1
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18377_ _01939_ _01940_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__nand2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15589_ _08218_ _08232_ _08208_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__and3_1
XFILLER_147_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17328_ _04016_ _09739_ vssd1 vssd1 vccd1 vccd1 _09896_ sky130_fd_sc_hd__nand2_1
XFILLER_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17259_ _05531_ _09069_ vssd1 vssd1 vccd1 vccd1 _09835_ sky130_fd_sc_hd__nand2_1
XFILLER_88_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20131__162 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__inv_2
XFILLER_97_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21655_ clknet_leaf_87_i_clk _01424_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20606_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__nand2_1
XFILLER_166_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21586_ net507 _01355_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_76 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_76/HI o_rgb[4] sky130_fd_sc_hd__conb_1
XFILLER_181_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_87 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_87/HI o_rgb[19] sky130_fd_sc_hd__conb_1
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xtop_ew_algofoogle_98 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_98/HI zeros[8] sky130_fd_sc_hd__conb_1
X_20537_ _03426_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__xnor2_1
XFILLER_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20468_ _03367_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nand3_1
X_11270_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _04050_
+ sky130_fd_sc_hd__or2_1
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20214__237 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__inv_2
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14960_ rbzero.wall_tracer.visualWallDist\[11\] _07595_ _07649_ _07642_ vssd1 vssd1
+ vccd1 vccd1 _00466_ sky130_fd_sc_hd__o211a_1
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _06569_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14891_ _07601_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__clkinv_2
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16630_ _09271_ _09272_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__xnor2_1
X_13842_ _06259_ _06575_ _06578_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16561_ _09059_ _09193_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__and2b_1
X_13773_ _05823_ _06045_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__nor2_1
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ _03840_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18300_ _01998_ _01999_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__xor2_1
X_15512_ rbzero.wall_tracer.visualWallDist\[4\] _08148_ vssd1 vssd1 vccd1 vccd1 _08157_
+ sky130_fd_sc_hd__nand2_2
X_12724_ _05470_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__xnor2_4
X_19280_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_leak\[2\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16492_ _07566_ _07568_ _07571_ _08220_ _07575_ vssd1 vssd1 vccd1 vccd1 _09136_ sky130_fd_sc_hd__o41a_1
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20295__309 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__inv_2
XFILLER_188_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18231_ _01875_ _01857_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__or2b_1
X_15443_ rbzero.debug_overlay.playerY\[-2\] _08029_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ rbzero.wall_tracer.mapY\[5\] _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11606_ rbzero.tex_r1\[51\] rbzero.tex_r1\[50\] _04338_ vssd1 vssd1 vccd1 vccd1 _04385_
+ sky130_fd_sc_hd__mux2_1
X_18162_ _01739_ _01620_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__or3_1
XFILLER_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15374_ _04013_ _08017_ _08018_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__a21oi_4
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ _05338_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__and2_1
X_17113_ _04814_ _03474_ vssd1 vssd1 vccd1 vccd1 _09751_ sky130_fd_sc_hd__or2_1
X_14325_ _06245_ _06708_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__or2_1
XFILLER_157_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11537_ gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__buf_2
X_18093_ _01678_ _01680_ _01679_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__o21bai_1
XFILLER_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17044_ _08767_ _09417_ vssd1 vssd1 vccd1 vccd1 _09684_ sky130_fd_sc_hd__nor2_1
X_14256_ _06982_ _06989_ _06991_ _06992_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__a211oi_1
X_11468_ _04245_ _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux2_1
XFILLER_183_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13207_ _05700_ _05879_ _05881_ _05887_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a211o_2
X_10419_ _03541_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14187_ _06894_ _06896_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__xnor2_1
X_11399_ _04153_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__nor2_1
X_20189__214 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__inv_2
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13138_ _05703_ _05871_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__or3_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _02628_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__clkbuf_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _05777_ _05796_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__xnor2_1
X_17946_ _01523_ _01529_ _10271_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a21o_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17877_ _01578_ _01579_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16828_ rbzero.wall_tracer.texu\[3\] _09085_ _09468_ _09469_ _07642_ vssd1 vssd1
+ vccd1 vccd1 _00514_ sky130_fd_sc_hd__o221a_1
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19547_ rbzero.pov.spi_counter\[0\] _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 _03021_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16759_ _09252_ _09394_ _09399_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__and3_1
XFILLER_179_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19478_ _04034_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__nor2_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18429_ _01799_ _02024_ _02025_ _02023_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a221o_2
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21440_ net361 _01209_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21371_ net292 _01140_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19635__87 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__inv_2
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10770_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _03718_ vssd1 vssd1 vccd1 vccd1 _03728_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12440_ _05198_ _03914_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__nor2_1
XFILLER_185_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21638_ clknet_leaf_18_i_clk _01407_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12371_ net35 net36 net37 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__nor3_1
XFILLER_181_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21569_ net490 _01338_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ _06666_ _06678_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__nor2_1
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _04055_ _04054_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nand2_1
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15090_ _07748_ _07749_ _07736_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__o21ai_1
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14041_ _06012_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__and3_1
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11253_ _04034_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__buf_4
XFILLER_180_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ rbzero.map_rom.f2 rbzero.map_rom.f1 rbzero.map_rom.i_col\[4\] vssd1 vssd1
+ vccd1 vccd1 _03973_ sky130_fd_sc_hd__and3_1
XFILLER_122_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17800_ _09668_ _09552_ _09973_ _08802_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o22a_1
X_15992_ _08634_ _08636_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18780_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__nor2_1
XFILLER_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14943_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.trackDistX\[6\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__mux2_1
X_17731_ _10294_ _10184_ _10185_ vssd1 vssd1 vccd1 vccd1 _10296_ sky130_fd_sc_hd__or3_1
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14874_ _07452_ _07451_ _05892_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__mux2_1
X_17662_ _10070_ _10079_ _10226_ vssd1 vssd1 vccd1 vccd1 _10227_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ _02873_ _02884_ _02885_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__or3_1
X_13825_ _06561_ _06276_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__xor2_1
X_16613_ _09254_ _09255_ vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17593_ _10156_ _10158_ vssd1 vssd1 vccd1 vccd1 _10159_ sky130_fd_sc_hd__xor2_1
X_16544_ _09186_ _09187_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__xnor2_2
X_19332_ rbzero.pov.spi_done rbzero.pov.ready _02730_ _02823_ vssd1 vssd1 vccd1 vccd1
+ _00804_ sky130_fd_sc_hd__o211a_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13756_ _06491_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__nor2_1
X_10968_ rbzero.tex_b1\[8\] rbzero.tex_b1\[9\] _03828_ vssd1 vssd1 vccd1 vccd1 _03832_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12707_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] _05446_
+ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a21bo_1
XFILLER_204_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19263_ _02785_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16475_ _08284_ _08177_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__nor2_2
X_13687_ _06422_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__and2_1
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10899_ rbzero.tex_b1\[41\] rbzero.tex_b1\[42\] _03795_ vssd1 vssd1 vccd1 vccd1 _03796_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18214_ _01908_ _01914_ rbzero.wall_tracer.trackDistX\[6\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00595_ sky130_fd_sc_hd__o2bb2a_1
X_15426_ _08070_ rbzero.debug_overlay.playerY\[-3\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _08071_ sky130_fd_sc_hd__mux2_1
X_19194_ rbzero.spi_registers.new_sky\[1\] rbzero.color_sky\[1\] _02740_ vssd1 vssd1
+ vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
X_12638_ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__inv_2
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18145_ _01844_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__nand2_1
X_15357_ _07904_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__clkbuf_4
XFILLER_200_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12569_ _05321_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__and2_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14308_ _06134_ _06662_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__nor2_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18076_ _01653_ _01654_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__nor2_1
X_15288_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__buf_4
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17027_ _09665_ _09666_ vssd1 vssd1 vccd1 vccd1 _09667_ sky130_fd_sc_hd__nand2_1
X_14239_ _06970_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__xor2_1
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _02619_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17929_ _01613_ _01631_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__xor2_2
XFILLER_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20940_ clknet_leaf_67_i_clk _00709_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19640__90 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__inv_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20871_ clknet_leaf_63_i_clk _00640_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20243__263 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__inv_2
XFILLER_41_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21423_ net344 _01192_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21354_ net275 _01123_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20305_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__buf_1
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21285_ clknet_leaf_34_i_clk _01054_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20326__338 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__inv_2
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _04230_ _04711_ _04715_ _04242_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a211o_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ _04646_ _04647_ _04217_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__mux2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _06345_ _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nor2_1
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _03755_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _07203_ _07210_ _07154_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__a21oi_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13541_ _06193_ _06231_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__xor2_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _03719_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _08902_ _08904_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__nor2_1
X_13472_ _06168_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ rbzero.tex_g1\[15\] rbzero.tex_g1\[16\] _03680_ vssd1 vssd1 vccd1 vccd1 _03683_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _04034_ _07861_ _07862_ _07718_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__o31a_1
XFILLER_185_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__buf_2
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16191_ _08815_ _08835_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__xor2_1
XFILLER_166_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ _07786_ _07789_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__and2_1
X_12354_ _05101_ _05120_ _05121_ net31 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o211a_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20071__108 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__inv_2
X_11305_ rbzero.traced_texVinit\[1\] rbzero.texV\[1\] rbzero.texV\[0\] rbzero.traced_texVinit\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__o211a_1
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15073_ _07732_ _07733_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__xnor2_1
X_19950_ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__clkbuf_2
X_12285_ net46 _05046_ _05049_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a22o_1
XFILLER_142_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14024_ _05752_ _06658_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nand2_4
X_18901_ rbzero.spi_registers.spi_counter\[3\] _02564_ _02570_ vssd1 vssd1 vccd1 vccd1
+ _02571_ sky130_fd_sc_hd__o21a_1
XFILLER_84_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11236_ gpout0.hpos\[9\] _04009_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__and2_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19881_ _03188_ _03186_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__nor2_1
XFILLER_84_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18832_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__or2_1
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11167_ rbzero.otherx\[1\] rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__xor2_1
XFILLER_136_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18763_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__nor2_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19614__68 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
X_15975_ _08609_ _08611_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__xnor2_1
X_11098_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _03898_ vssd1 vssd1 vccd1 vccd1 _03900_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17714_ _10109_ _10151_ _10278_ vssd1 vssd1 vccd1 vccd1 _10279_ sky130_fd_sc_hd__a21bo_1
XFILLER_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14926_ rbzero.wall_tracer.visualWallDist\[0\] _07618_ vssd1 vssd1 vccd1 vccd1 _07627_
+ sky130_fd_sc_hd__or2_1
X_18694_ _09889_ _02388_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__or3b_1
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17645_ _09096_ _09359_ _10060_ _10059_ vssd1 vssd1 vccd1 vccd1 _10210_ sky130_fd_sc_hd__o31a_1
XFILLER_64_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14857_ _07468_ _07574_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__nand2b_4
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _06490_ _06493_ _06494_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__or3_1
XFILLER_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14788_ _05884_ _07477_ _07419_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__or3_1
X_17576_ _10137_ _10140_ _10141_ vssd1 vssd1 vccd1 vccd1 _10142_ sky130_fd_sc_hd__and3_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19315_ rbzero.spi_registers.new_vshift\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13739_ _06045_ _06009_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__nor2_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16527_ _09169_ _09170_ vssd1 vssd1 vccd1 vccd1 _09171_ sky130_fd_sc_hd__nand2_1
XFILLER_108_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19246_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_sky\[1\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ _09100_ _09101_ vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15409_ _08053_ vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__04835_ clknet_0__04835_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04835_
+ sky130_fd_sc_hd__clkbuf_16
X_19177_ rbzero.spi_registers.got_new_leak _02711_ vssd1 vssd1 vccd1 vccd1 _02733_
+ sky130_fd_sc_hd__nand2_1
X_16389_ _09032_ _09033_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__nand2_1
XFILLER_192_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18128_ _01827_ _01828_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20273__289 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__inv_2
X_18059_ _01757_ _01758_ _01759_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a21o_1
XFILLER_160_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21070_ net160 _00839_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20021_ _04990_ _04989_ _03258_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or4_1
XFILLER_141_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167__194 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__inv_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20923_ clknet_leaf_73_i_clk _00692_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20384__10 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20854_ clknet_leaf_1_i_clk _00623_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20785_ clknet_leaf_21_i_clk _00554_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_57_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21406_ net327 _01175_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21337_ net258 _01106_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ _04840_ _04666_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nand2_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21268_ clknet_leaf_62_i_clk _01037_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11021_ _03859_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21199_ clknet_leaf_48_i_clk _00968_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi sky130_fd_sc_hd__dfxtp_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _08337_ _08347_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__xnor2_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _05563_ _05566_ _05600_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__and3_1
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _07375_ _07447_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__or2_1
X_11923_ _04241_ _04690_ _04698_ _04207_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__o211a_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _08059_ _08335_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__nor2_1
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _07378_ _07349_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__nand2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17430_ _07601_ _09995_ _09996_ vssd1 vssd1 vccd1 vccd1 _09997_ sky130_fd_sc_hd__mux2_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11854_ rbzero.tex_g1\[13\] rbzero.tex_g1\[12\] _04337_ vssd1 vssd1 vccd1 vccd1 _04631_
+ sky130_fd_sc_hd__mux2_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _03746_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14573_ _07305_ _07093_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__xnor2_1
X_17361_ _09243_ _09029_ _09164_ _09096_ vssd1 vssd1 vccd1 vccd1 _09928_ sky130_fd_sc_hd__o22ai_1
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ _04560_ _04561_ _04562_ _04304_ _04253_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__o221a_1
XFILLER_41_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19100_ _02683_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__clkbuf_1
X_13524_ _06259_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nor2_1
X_16312_ _08550_ _08616_ _08673_ _08955_ _08956_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__o221ai_4
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17292_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09864_ sky130_fd_sc_hd__or2_1
X_10736_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _03706_ vssd1 vssd1 vccd1 vccd1 _03710_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19031_ rbzero.pov.spi_buffer\[47\] rbzero.pov.ready_buffer\[47\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
X_16243_ _08871_ _08887_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__nand2_1
X_13455_ _06189_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ rbzero.tex_g1\[23\] rbzero.tex_g1\[24\] _03669_ vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ _04883_ _04884_ _04886_ _04887_ _05143_ net34 vssd1 vssd1 vccd1 vccd1 _05173_
+ sky130_fd_sc_hd__mux4_1
X_16174_ _08816_ _08075_ _08817_ _08784_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__o22a_1
X_13386_ _06041_ _05991_ _05940_ _06078_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__o22ai_1
XFILLER_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10598_ _03637_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15125_ _07782_ vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__clkbuf_1
X_12337_ net46 _05103_ _05104_ _05099_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ rbzero.wall_tracer.rayAddendX\[-3\] _07717_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07719_ sky130_fd_sc_hd__mux2_1
X_19933_ rbzero.debug_overlay.playerY\[3\] _03223_ _02822_ vssd1 vssd1 vccd1 vccd1
+ _03228_ sky130_fd_sc_hd__a21o_1
X_12268_ _04886_ _04887_ _05021_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__mux2_1
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14007_ _06666_ _06708_ _06742_ _06743_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__o31ai_2
XFILLER_141_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__buf_2
X_19864_ rbzero.debug_overlay.playerX\[1\] _03143_ _03174_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00984_ sky130_fd_sc_hd__a211o_1
X_12199_ net17 net18 vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__nand2_1
XFILLER_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18815_ _05532_ _02494_ _02495_ _02399_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__o31a_1
XFILLER_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20309__322 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__inv_2
X_19795_ _03126_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18746_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__nor2_1
X_15958_ _08588_ _08600_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__03295_ clknet_0__03295_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03295_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14909_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.trackDistX\[-4\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__mux2_1
X_18677_ _02368_ _02372_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__xnor2_1
X_15889_ _08531_ _08532_ _08533_ vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17628_ _10085_ _10187_ _10191_ vssd1 vssd1 vccd1 vccd1 _10193_ sky130_fd_sc_hd__and3_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ _08747_ _09700_ vssd1 vssd1 vccd1 vccd1 _10125_ sky130_fd_sc_hd__nor2_1
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20570_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__nand2_1
XFILLER_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19229_ rbzero.spi_registers.new_vshift\[1\] _02763_ vssd1 vssd1 vccd1 vccd1 _02766_
+ sky130_fd_sc_hd__or2_1
XFILLER_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20355__364 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__inv_2
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21122_ net212 _00891_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21053_ clknet_leaf_57_i_clk _00822_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20004_ rbzero.pov.ready_buffer\[8\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[-1\]
+ _02730_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__o221a_1
XFILLER_101_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20906_ clknet_leaf_63_i_clk _00675_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20837_ clknet_leaf_24_i_clk _00606_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11570_ rbzero.tex_r1\[3\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and3_1
X_20768_ clknet_leaf_24_i_clk _00537_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_161_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10521_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _03591_ vssd1 vssd1 vccd1 vccd1 _03597_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20699_ clknet_leaf_5_i_clk _00483_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13240_ _05962_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__nand2_1
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10452_ rbzero.tex_r0\[62\] rbzero.tex_r0\[61\] _03558_ vssd1 vssd1 vccd1 vccd1 _03561_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13171_ _05884_ _05859_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__or2_1
X_10383_ _03522_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12122_ _04885_ _04888_ _04889_ _04893_ net4 net3 vssd1 vssd1 vccd1 vccd1 _04894_
+ sky130_fd_sc_hd__mux4_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12053_ rbzero.row_render.side _04821_ _04826_ _04814_ _04820_ vssd1 vssd1 vccd1
+ vccd1 _04827_ sky130_fd_sc_hd__o221ai_1
X_16930_ _09559_ _09570_ vssd1 vssd1 vccd1 vccd1 _09571_ sky130_fd_sc_hd__xnor2_2
XFILLER_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ _03850_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16861_ _09243_ _08159_ _08150_ _09245_ vssd1 vssd1 vccd1 vccd1 _09502_ sky130_fd_sc_hd__o22a_1
XFILLER_133_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18600_ _02179_ _02182_ _02295_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__and3_1
X_15812_ _08025_ _08013_ vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16792_ _09429_ _09433_ _05209_ vssd1 vssd1 vccd1 vccd1 _09434_ sky130_fd_sc_hd__a21o_2
XFILLER_93_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18531_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__or2_1
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12955_ _05642_ _05645_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__or2_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _08386_ _08387_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__xnor2_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11906_ _04332_ _04677_ _04681_ _04142_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a211o_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _02143_ _02159_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12886_ _05609_ _05619_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__or3_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _08263_ _08264_ _08307_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__and3_1
XFILLER_206_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17413_ _08284_ _09540_ vssd1 vssd1 vccd1 vccd1 _09980_ sky130_fd_sc_hd__nor2_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _07357_ _07361_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__or2_1
X_11837_ rbzero.tex_g1\[45\] rbzero.tex_g1\[44\] _04337_ vssd1 vssd1 vccd1 vccd1 _04614_
+ sky130_fd_sc_hd__mux2_1
X_18393_ _02086_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14556_ _07286_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__nor2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _08335_ _09359_ _09910_ _09624_ vssd1 vssd1 vccd1 vccd1 _09911_ sky130_fd_sc_hd__o31a_1
XFILLER_159_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11768_ _04542_ _04545_ _04208_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
XFILLER_201_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13507_ _05983_ _05940_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__or3_1
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10719_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _03624_ vssd1 vssd1 vccd1 vccd1 _03701_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14487_ _07177_ _07009_ _07223_ _07065_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a22o_1
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17275_ _09846_ _09847_ _09848_ vssd1 vssd1 vccd1 vccd1 _09849_ sky130_fd_sc_hd__and3_1
XFILLER_140_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11699_ rbzero.debug_overlay.vplaneY\[10\] _04453_ _04474_ _04477_ vssd1 vssd1 vccd1
+ vccd1 _04478_ sky130_fd_sc_hd__a211o_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19014_ _02594_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__buf_4
X_13438_ _05998_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__or2_1
X_16226_ _08870_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__inv_2
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16157_ _08111_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__buf_4
X_13369_ _06099_ _06102_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__nand3_1
XFILLER_155_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _07749_ _07766_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__xnor2_1
X_16088_ _08284_ _08128_ _08727_ _08732_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__o31ai_1
XFILLER_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15039_ _03913_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__clkbuf_4
X_19916_ _08089_ _03164_ _03193_ _03214_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a211oi_1
XFILLER_111_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19847_ rbzero.pov.ready_buffer\[66\] _08077_ _03146_ vssd1 vssd1 vccd1 vccd1 _03162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19778_ rbzero.pov.spi_buffer\[62\] rbzero.pov.spi_buffer\[63\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_209_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18729_ _02420_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20622_ clknet_leaf_73_i_clk _00406_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_189_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20279__295 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__inv_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20553_ _03436_ _03439_ _03440_ _09748_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a31o_1
XFILLER_165_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20484_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03384_
+ sky130_fd_sc_hd__nand2_1
XFILLER_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21105_ net195 _00874_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21036_ clknet_leaf_79_i_clk _00805_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _05486_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__xnor2_2
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__nor2_1
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ _07120_ _07126_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__or2_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ rbzero.tex_r1\[33\] rbzero.tex_r1\[32\] _04392_ vssd1 vssd1 vccd1 vccd1 _04401_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__buf_2
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14341_ _07017_ _07019_ _06774_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__o21ai_1
XFILLER_204_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _04208_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__buf_4
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10504_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _03580_ vssd1 vssd1 vccd1 vccd1 _03588_
+ sky130_fd_sc_hd__mux2_1
X_17060_ _08816_ _09699_ vssd1 vssd1 vccd1 vccd1 _09700_ sky130_fd_sc_hd__or2_1
X_14272_ _06675_ _06740_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__nor2_1
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11484_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _04263_ vssd1 vssd1 vccd1 vccd1 _04264_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16011_ _08634_ _08636_ _08655_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__a21bo_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13223_ _05901_ _05831_ _05956_ _05959_ _05871_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_1_0__f__03298_ clknet_0__03298_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03298_
+ sky130_fd_sc_hd__clkbuf_16
X_10435_ rbzero.tex_r1\[3\] rbzero.tex_r1\[4\] _03549_ vssd1 vssd1 vccd1 vccd1 _03550_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _05872_ _05890_ _05826_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__mux2_1
X_10366_ _03513_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12105_ net5 _04850_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__or2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _05814_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__or2_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _01546_ _01442_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__or2b_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19701_ _03077_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__clkbuf_1
X_12036_ _04317_ _04163_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nor2_1
X_16913_ rbzero.wall_tracer.stepDistX\[7\] vssd1 vssd1 vccd1 vccd1 _09554_ sky130_fd_sc_hd__clkinv_2
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17893_ _01594_ _01595_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__03301_ _03301_ vssd1 vssd1 vccd1 vccd1 clknet_0__03301_ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _08160_ _09480_ _09484_ _08162_ vssd1 vssd1 vccd1 vccd1 _09485_ sky130_fd_sc_hd__o22ai_1
XFILLER_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19563_ _03031_ _03020_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and3b_1
XFILLER_81_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16775_ _09416_ vssd1 vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__clkbuf_4
X_13987_ _06067_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18514_ _02205_ _02206_ _02210_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__and3_1
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15726_ _08327_ _08370_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__xnor2_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ _05659_ _05603_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__nand2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ _02904_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02973_
+ sky130_fd_sc_hd__nand2_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18445_ _02044_ _02052_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a21o_1
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _08300_ _08301_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__xnor2_2
X_12869_ _05603_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nand2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _07330_ _07342_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18376_ _02073_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__xor2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ _08218_ _08208_ _08232_ vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17327_ rbzero.wall_tracer.trackDistX\[-2\] _09817_ _09888_ _09895_ vssd1 vssd1 vccd1
+ vccd1 _00587_ sky130_fd_sc_hd__o22a_1
X_14539_ _07274_ _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__nor2_1
XFILLER_144_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17258_ _09830_ _09831_ _09832_ vssd1 vssd1 vccd1 vccd1 _09834_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16209_ _08519_ _08053_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__nor2_1
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17189_ rbzero.wall_tracer.mapX\[6\] _05512_ vssd1 vssd1 vccd1 vccd1 _09774_ sky130_fd_sc_hd__xor2_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21654_ clknet_3_7_0_i_clk _01423_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20605_ gpout3.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nor2_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21585_ net506 _01354_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_77 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_77/HI o_rgb[5] sky130_fd_sc_hd__conb_1
X_20536_ rbzero.traced_texa\[7\] rbzero.texV\[7\] _03427_ vssd1 vssd1 vccd1 vccd1
+ _03428_ sky130_fd_sc_hd__o21ai_1
XFILLER_166_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_88 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_88/HI o_rgb[20] sky130_fd_sc_hd__conb_1
XFILLER_165_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_99 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_99/HI zeros[9] sky130_fd_sc_hd__conb_1
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20467_ _03367_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__a21o_1
XFILLER_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13910_ _05752_ _05989_ _06053_ _06624_ _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__a41o_1
XFILLER_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21019_ clknet_leaf_67_i_clk _00788_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14890_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1 vccd1 vccd1 _07601_
+ sky130_fd_sc_hd__buf_4
XFILLER_130_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13841_ _06576_ _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__and2_1
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13772_ _06508_ _06481_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__xnor2_1
X_16560_ _05194_ _09202_ _09203_ _07642_ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__o211a_1
X_10984_ rbzero.tex_b1\[0\] rbzero.tex_b1\[1\] _03482_ vssd1 vssd1 vccd1 vccd1 _03840_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _08056_ _08063_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__and2_1
X_12723_ _05422_ _05429_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and2b_1
X_16491_ _09133_ _09134_ vssd1 vssd1 vccd1 vccd1 _09135_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18230_ _01874_ _01858_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or2b_1
XFILLER_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15442_ _08076_ _08085_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__nand2_1
X_12654_ _05397_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__clkbuf_4
XFILLER_130_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11605_ rbzero.tex_r1\[49\] rbzero.tex_r1\[48\] _04338_ vssd1 vssd1 vccd1 vccd1 _04384_
+ sky130_fd_sc_hd__mux2_1
X_18161_ _01859_ _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__nand2_1
XFILLER_180_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15373_ _07903_ rbzero.wall_tracer.stepDistY\[-7\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _08018_ sky130_fd_sc_hd__a21o_1
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ _05296_ _05297_ _05337_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__nand3b_1
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17112_ _09749_ vssd1 vssd1 vccd1 vccd1 _09750_ sky130_fd_sc_hd__clkbuf_4
X_14324_ _07060_ _06843_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nand2_1
X_11536_ gpout0.vpos\[5\] gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nand2_1
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18092_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__nand2_1
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14255_ _06962_ _06984_ _06988_ _06951_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__o22a_1
X_17043_ _09553_ _09557_ _09556_ vssd1 vssd1 vccd1 vccd1 _09683_ sky130_fd_sc_hd__a21bo_1
X_11467_ _04139_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__buf_4
XFILLER_143_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _05846_ _05940_ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__or3_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10418_ rbzero.tex_r1\[11\] rbzero.tex_r1\[12\] _03538_ vssd1 vssd1 vccd1 vccd1 _03541_
+ sky130_fd_sc_hd__mux2_1
X_14186_ _06921_ _06922_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11398_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] _04152_ vssd1 vssd1
+ vccd1 vccd1 _04178_ sky130_fd_sc_hd__nor3_1
XFILLER_124_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13137_ _05778_ _05872_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__o21a_1
XFILLER_139_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _03504_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18994_ rbzero.pov.spi_buffer\[29\] rbzero.pov.ready_buffer\[29\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13068_ _05721_ _05734_ _05796_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__mux2_1
X_17945_ _01643_ _01644_ _01646_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a21o_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12019_ _04379_ _04791_ _04792_ _04793_ _04209_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__o221a_1
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17876_ _09096_ _09703_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__nand2_1
XFILLER_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19615_ clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__buf_1
X_16827_ _09082_ _09467_ _05194_ vssd1 vssd1 vccd1 vccd1 _09469_ sky130_fd_sc_hd__a21o_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19546_ rbzero.pov.ss_buffer\[1\] _03555_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nor2_4
XFILLER_0_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16758_ _09252_ _09394_ _09399_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15709_ _08352_ _08353_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__nand2_1
X_19477_ _02941_ _02944_ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__o21a_1
XFILLER_179_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16689_ rbzero.debug_overlay.playerY\[-4\] vssd1 vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__clkinv_2
XFILLER_146_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18428_ _02125_ _02126_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__nand2_1
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18359_ _02056_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__nor2_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21370_ net291 _01139_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20183_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__buf_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20220__242 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__inv_2
XFILLER_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21637_ clknet_leaf_18_i_clk _01406_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12370_ _04738_ _05086_ _05098_ _05137_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__o2bb2a_2
XFILLER_166_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21568_ net489 _01337_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _04060_ _04063_ _04100_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__o21ba_1
XFILLER_126_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20519_ _03406_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__o21ai_1
XFILLER_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21499_ net420 _01268_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _06776_ _06658_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__nor2_1
XFILLER_180_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11252_ _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__buf_4
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ rbzero.map_rom.d6 _03942_ _03933_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_
+ sky130_fd_sc_hd__and4_1
XFILLER_161_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15991_ _08635_ _08561_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17730_ _10184_ _10185_ _10294_ vssd1 vssd1 vccd1 vccd1 _10295_ sky130_fd_sc_hd__o21a_1
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14942_ _07621_ _07636_ _07637_ _07620_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__o211a_1
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17661_ _10071_ _09961_ _10078_ vssd1 vssd1 vccd1 vccd1 _10226_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14873_ _07587_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19400_ _02884_ _02885_ _02873_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16612_ _07996_ _09103_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__or2_1
X_13824_ _06193_ _06231_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nand2_1
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17592_ _09955_ _10014_ _10157_ vssd1 vssd1 vccd1 vccd1 _10158_ sky130_fd_sc_hd__a21boi_1
XFILLER_211_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20303__317 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__inv_2
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19331_ _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16543_ _09046_ _09048_ _09045_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__a21boi_2
XFILLER_44_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13755_ _06467_ _06489_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__xor2_1
X_10967_ _03831_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19262_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_floor\[1\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
X_12706_ _05450_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__xnor2_2
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16474_ _08178_ _09117_ _08972_ _08973_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__o31ai_4
X_13686_ _06336_ _06375_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__xor2_1
X_10898_ _03646_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ _01912_ _01913_ _09780_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15425_ _08029_ _08069_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__and2_1
XFILLER_188_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19193_ rbzero.color_sky\[0\] _02740_ _02742_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__a21o_1
XFILLER_54_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12637_ rbzero.map_rom.a6 _05374_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__and2_1
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18144_ _10239_ _08423_ _01843_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__o21ai_1
XFILLER_129_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12568_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__nand2_1
X_15356_ _07999_ _08000_ _05496_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__mux2_1
XFILLER_200_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11519_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _04263_ vssd1 vssd1 vccd1 vccd1 _04299_
+ sky130_fd_sc_hd__mux2_1
X_14307_ _07005_ _06731_ _06700_ _07004_ _07003_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__o32ai_4
XFILLER_172_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18075_ _01775_ _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__or2_1
X_15287_ _07931_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12499_ rbzero.wall_tracer.trackDistY\[2\] vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__inv_2
X_17026_ _09661_ _08047_ _09662_ _09664_ vssd1 vssd1 vccd1 vccd1 _09666_ sky130_fd_sc_hd__a2bb2o_1
X_14238_ _06935_ _06963_ _06972_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__a31o_1
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ _06904_ _06903_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__and2b_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ rbzero.pov.spi_buffer\[21\] rbzero.pov.ready_buffer\[21\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XFILLER_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _01615_ _01630_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__xor2_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17859_ _01491_ _01455_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__or2b_1
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20870_ clknet_leaf_60_i_clk _00639_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19529_ _02994_ _02995_ _02998_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21422_ net343 _01191_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21353_ net274 _01122_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21284_ clknet_leaf_39_i_clk _01053_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11870_ rbzero.tex_g1\[17\] rbzero.tex_g1\[16\] _04211_ vssd1 vssd1 vccd1 vccd1 _04647_
+ sky130_fd_sc_hd__mux2_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _03751_ vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__mux2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ clknet_leaf_51_i_clk _00768_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13540_ _06193_ _06231_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__and3_1
XFILLER_198_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ rbzero.tex_g0\[48\] rbzero.tex_g0\[47\] _03718_ vssd1 vssd1 vccd1 vccd1 _03719_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _06199_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ _03682_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15210_ _07850_ _07854_ _07860_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__a21oi_1
X_12422_ net71 rbzero.wall_tracer.state\[9\] _03480_ vssd1 vssd1 vccd1 vccd1 _05187_
+ sky130_fd_sc_hd__and3_1
XFILLER_139_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16190_ _08827_ _08833_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12353_ net29 _05094_ net30 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__o21ai_1
X_15141_ _07785_ rbzero.wall_tracer.rayAddendX\[4\] vssd1 vssd1 vccd1 vccd1 _07797_
+ sky130_fd_sc_hd__xor2_1
XFILLER_126_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ rbzero.texV\[3\] _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__xor2_1
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15072_ _07721_ _07724_ _07722_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__a21bo_1
X_12284_ _04867_ _05034_ _05027_ net47 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a31o_1
XFILLER_181_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14023_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nand2_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18900_ rbzero.spi_registers.spi_counter\[1\] _02569_ vssd1 vssd1 vccd1 vccd1 _02570_
+ sky130_fd_sc_hd__xnor2_1
X_11235_ _04015_ _04019_ _03914_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a21oi_1
XFILLER_122_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19880_ rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__inv_2
XFILLER_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _02509_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
X_11166_ _03915_ _03918_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__o21a_1
XFILLER_132_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18762_ _02449_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15974_ _08584_ _08618_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__xnor2_4
X_11097_ _03899_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17713_ _10147_ _10150_ vssd1 vssd1 vccd1 vccd1 _10278_ sky130_fd_sc_hd__or2b_1
X_14925_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.trackDistX\[0\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__mux2_1
X_18693_ _02310_ _02313_ _02387_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__or3_1
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _10207_ _10208_ vssd1 vssd1 vccd1 vccd1 _10209_ sky130_fd_sc_hd__xnor2_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ _07433_ _07374_ _07573_ _07394_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__o211ai_4
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ _06505_ _06524_ _06525_ _06543_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__o211a_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _08872_ _10139_ _08266_ _09989_ vssd1 vssd1 vccd1 vccd1 _10141_ sky130_fd_sc_hd__a2bb2o_1
X_14787_ _05884_ _07516_ _07518_ _05800_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__a211o_1
XFILLER_95_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ _04772_ _04773_ _04225_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19314_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__buf_2
XFILLER_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16526_ _08112_ _08150_ _08331_ _08417_ vssd1 vssd1 vccd1 vccd1 _09170_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13738_ _05846_ _05823_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__nor2_1
XFILLER_182_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19245_ _02775_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__clkbuf_1
X_16457_ _07932_ _08097_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__or2_1
X_13669_ _05856_ _05877_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15408_ _07903_ _08048_ _08051_ _08052_ _05196_ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__o311a_2
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19176_ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__clkbuf_2
XFILLER_118_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16388_ _08053_ _08158_ _08418_ _08039_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_185_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18127_ _10094_ _09027_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nor2_1
X_15339_ rbzero.wall_tracer.visualWallDist\[-8\] _07983_ _07903_ vssd1 vssd1 vccd1
+ vccd1 _07984_ sky130_fd_sc_hd__mux2_1
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18058_ _01757_ _01758_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__nand3_1
XFILLER_126_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17009_ _09499_ _09506_ _09648_ vssd1 vssd1 vccd1 vccd1 _09649_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20020_ _04891_ _04887_ _04886_ _04890_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__or4b_1
XFILLER_154_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20922_ clknet_leaf_69_i_clk _00691_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ clknet_leaf_1_i_clk _00622_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20784_ clknet_leaf_21_i_clk _00553_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21405_ net326 _01174_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21336_ net257 _01105_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[43\] sky130_fd_sc_hd__dfxtp_1
X_20332__343 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__inv_2
XFILLER_191_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21267_ clknet_leaf_82_i_clk _01036_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11020_ rbzero.tex_b0\[48\] rbzero.tex_b0\[47\] _03854_ vssd1 vssd1 vccd1 vccd1 _03859_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21198_ clknet_leaf_48_i_clk _00967_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20149_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__buf_1
X_20057__95 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__inv_2
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _05591_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nand2_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _05741_ _07402_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__nand2_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _04692_ _04694_ _04697_ _04332_ _04371_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a221o_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _08054_ vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__clkbuf_4
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14641_ _05793_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__buf_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11853_ rbzero.tex_g1\[15\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04630_
+ sky130_fd_sc_hd__a31o_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _09243_ _08821_ _09028_ _09164_ vssd1 vssd1 vccd1 vccd1 _09927_ sky130_fd_sc_hd__or4_1
X_10804_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _03740_ vssd1 vssd1 vccd1 vccd1 _03746_
+ sky130_fd_sc_hd__mux2_1
X_14572_ _07095_ _07096_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__nand2_1
X_11784_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _04212_ vssd1 vssd1 vccd1 vccd1 _04562_
+ sky130_fd_sc_hd__mux2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16311_ _08617_ _08672_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__nand2_1
XFILLER_201_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13523_ _05991_ _06080_ _06134_ _05978_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__o22a_1
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ _03709_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__clkbuf_1
X_17291_ _04016_ vssd1 vssd1 vccd1 vccd1 _09863_ sky130_fd_sc_hd__clkbuf_4
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ _02646_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ _08885_ _08886_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__and2_1
X_13454_ _06069_ _06074_ _06089_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__a31oi_2
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10666_ _03673_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12405_ _04989_ gpout0.vpos\[5\] _04891_ _04890_ _05143_ net34 vssd1 vssd1 vccd1
+ vccd1 _05172_ sky130_fd_sc_hd__mux4_1
X_13385_ _06094_ _06096_ _06095_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__a21boi_1
XFILLER_154_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16173_ _08816_ _08075_ _08817_ _08784_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__nor4_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10597_ rbzero.tex_g1\[56\] rbzero.tex_g1\[57\] _03635_ vssd1 vssd1 vccd1 vccd1 _03637_
+ sky130_fd_sc_hd__mux2_1
XFILLER_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ rbzero.wall_tracer.rayAddendX\[2\] _07781_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07782_ sky130_fd_sc_hd__mux2_1
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12336_ _04867_ _05081_ net47 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ _04883_ _04884_ _05021_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15055_ _04029_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__buf_4
X_19932_ rbzero.debug_overlay.playerY\[3\] _03223_ vssd1 vssd1 vccd1 vccd1 _03227_
+ sky130_fd_sc_hd__nor2_1
X_14006_ _06659_ _06741_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__nand2_1
X_11218_ gpout0.hpos\[4\] gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__and2_1
X_19863_ _03911_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__buf_4
X_12198_ _04966_ net61 _04967_ net18 vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__o211a_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18814_ _02492_ _02493_ _02487_ _02489_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__o211a_1
X_11149_ rbzero.debug_overlay.playerY\[2\] _03934_ _03935_ rbzero.debug_overlay.playerY\[4\]
+ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a221o_1
XFILLER_96_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19794_ rbzero.pov.spi_buffer\[70\] rbzero.pov.spi_buffer\[71\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18745_ _02434_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15957_ _08562_ _08558_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__xnor2_2
XFILLER_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03294_ clknet_0__03294_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03294_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14908_ _07591_ _07612_ _07613_ _04039_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__o211a_1
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18676_ _02369_ _02371_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _08514_ _08530_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__nor2_1
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17627_ _10085_ _10187_ _10191_ vssd1 vssd1 vccd1 vccd1 _10192_ sky130_fd_sc_hd__a21oi_1
X_14839_ _07459_ _07444_ _07468_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__o21bai_4
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17558_ _09994_ _10002_ _10123_ vssd1 vssd1 vccd1 vccd1 _10124_ sky130_fd_sc_hd__a21bo_1
XFILLER_147_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _09113_ _09152_ vssd1 vssd1 vccd1 vccd1 _09153_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17489_ _10053_ _10054_ vssd1 vssd1 vccd1 vccd1 _10055_ sky130_fd_sc_hd__nand2_1
XFILLER_177_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19228_ rbzero.spi_registers.vshift\[0\] _02762_ _02764_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00758_ sky130_fd_sc_hd__o211a_1
XFILLER_192_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19159_ rbzero.spi_registers.new_other\[1\] _02712_ vssd1 vssd1 vccd1 vccd1 _02720_
+ sky130_fd_sc_hd__or2_1
XFILLER_121_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21121_ net211 _00890_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21052_ clknet_leaf_3_i_clk _00821_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20003_ rbzero.pov.ready_buffer\[7\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-2\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__a221o_1
XFILLER_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ clknet_leaf_62_i_clk _00674_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ clknet_leaf_28_i_clk _00605_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20767_ clknet_leaf_32_i_clk _00536_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ _03596_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20698_ clknet_leaf_5_i_clk _00482_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _03560_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _05800_ _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__or2_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10382_ rbzero.tex_r1\[28\] rbzero.tex_r1\[29\] _03516_ vssd1 vssd1 vccd1 vccd1 _03522_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12121_ _04890_ _04891_ _04892_ gpout0.vpos\[0\] _04852_ _04846_ vssd1 vssd1 vccd1
+ vccd1 _04893_ sky130_fd_sc_hd__mux4_1
XFILLER_191_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21319_ net240 _01088_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ rbzero.row_render.texu\[5\] rbzero.row_render.texu\[4\] _03473_ vssd1 vssd1
+ vccd1 vccd1 _04826_ sky130_fd_sc_hd__mux2_1
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11003_ rbzero.tex_b0\[56\] rbzero.tex_b0\[55\] _03843_ vssd1 vssd1 vccd1 vccd1 _03850_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16860_ _09096_ _08427_ vssd1 vssd1 vccd1 vccd1 _09501_ sky130_fd_sc_hd__nor2_1
XFILLER_120_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15811_ _08442_ _08455_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__xor2_1
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16791_ _09085_ _09431_ _09432_ _08235_ vssd1 vssd1 vccd1 vccd1 _09433_ sky130_fd_sc_hd__o31ai_4
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18530_ _02226_ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__or2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _07996_ _08194_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__nor2_1
X_12954_ _05690_ _05634_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__or2_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11905_ _04678_ _04679_ _04680_ _04345_ _04253_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__o221a_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _02144_ _02158_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _08263_ _08264_ _08307_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__a21o_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _04001_ _05490_ _05620_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__o2bb2a_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17412_ _09694_ _09701_ _09978_ vssd1 vssd1 vccd1 vccd1 _09979_ sky130_fd_sc_hd__a21bo_1
XFILLER_61_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _05893_ _07360_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__and2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _02089_ _02090_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__xor2_1
XFILLER_92_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _04611_ _04612_ _04304_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__mux2_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _08331_ _09621_ vssd1 vssd1 vccd1 vccd1 _09910_ sky130_fd_sc_hd__nand2_1
XFILLER_198_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14555_ _07287_ _07288_ _07291_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__o21a_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _04543_ _04544_ _04138_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_1
XFILLER_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20339__349 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__inv_2
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _06241_ _06242_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__nand2_1
X_17274_ _09838_ _09840_ _09839_ vssd1 vssd1 vccd1 vccd1 _09848_ sky130_fd_sc_hd__o21bai_1
X_10718_ _03700_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14486_ _06689_ _06708_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__nor2_1
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11698_ rbzero.debug_overlay.vplaneY\[-6\] _04475_ _04454_ rbzero.debug_overlay.vplaneY\[-5\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a221o_1
X_19013_ _02637_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16225_ _08868_ _08869_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__or2_1
X_13437_ _05943_ _06000_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__and2b_1
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10649_ _03664_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16156_ _08766_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__or2_1
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _06103_ _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_41_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15107_ _07764_ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__or2_1
X_12319_ _05083_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16087_ _08728_ _08731_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__or2b_1
XFILLER_114_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13299_ _06032_ _06033_ _06034_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__nand3_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15038_ _07700_ _07701_ _03914_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__a21oi_1
X_19915_ rbzero.pov.ready_buffer\[52\] _03164_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__nor2_1
XFILLER_190_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_i_clk clknet_opt_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19846_ _03139_ _03160_ _03161_ _03157_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__o211a_1
XFILLER_111_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16989_ _08075_ _08821_ _09028_ _08425_ vssd1 vssd1 vccd1 vccd1 _09629_ sky130_fd_sc_hd__or4_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19777_ _03117_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__clkbuf_1
X_20084__119 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__inv_2
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18728_ rbzero.wall_tracer.trackDistY\[-9\] _02419_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02420_ sky130_fd_sc_hd__mux2_1
XFILLER_209_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18659_ _01860_ _09027_ _09350_ _01498_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__o22ai_1
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20621_ clknet_leaf_74_i_clk _00405_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_row\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20552_ _03436_ _03439_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20483_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03383_
+ sky130_fd_sc_hd__or2_1
XFILLER_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_156_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21104_ net194 _00873_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21035_ clknet_leaf_64_i_clk _00804_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready sky130_fd_sc_hd__dfxtp_1
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nand2_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11621_ _04230_ _04395_ _04399_ _04371_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a211o_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20819_ clknet_leaf_6_i_clk _00588_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14340_ _07075_ _07076_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__and2_1
X_11552_ rbzero.tex_r1\[13\] rbzero.tex_r1\[12\] _04291_ vssd1 vssd1 vccd1 vccd1 _04331_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10503_ _03587_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14271_ _06245_ _06663_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__nor2_1
X_11483_ _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__clkbuf_8
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16010_ _08637_ _08629_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__or2b_1
Xclkbuf_1_0__f__03297_ clknet_0__03297_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03297_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10434_ _03482_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__buf_4
X_13222_ _05931_ _05911_ _05958_ _05928_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__o211a_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10365_ rbzero.tex_r1\[36\] rbzero.tex_r1\[37\] _03505_ vssd1 vssd1 vccd1 vccd1 _03513_
+ sky130_fd_sc_hd__mux2_1
X_13153_ _05773_ _05733_ _05792_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12104_ net4 _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__or2_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13084_ _05815_ _05819_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__mux2_1
XFILLER_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17961_ _01560_ _01663_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__xor2_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12035_ gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__clkbuf_4
XFILLER_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19700_ rbzero.pov.spi_buffer\[25\] rbzero.pov.spi_buffer\[26\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03077_ sky130_fd_sc_hd__mux2_1
X_16912_ _09117_ _09552_ vssd1 vssd1 vccd1 vccd1 _09553_ sky130_fd_sc_hd__nor2_2
X_17892_ _08202_ _01475_ _01476_ _08259_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__o22ai_1
XFILLER_104_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03300_ _03300_ vssd1 vssd1 vccd1 vccd1 clknet_0__03300_ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16843_ _09483_ vssd1 vssd1 vccd1 vccd1 _09484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19562_ rbzero.pov.spi_counter\[3\] rbzero.pov.spi_counter\[2\] _03022_ rbzero.pov.spi_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a31o_1
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16774_ _08242_ _09129_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__and2_1
XFILLER_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ _06720_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__or2b_1
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18513_ _02205_ _02206_ _02210_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a21oi_1
X_15725_ _08349_ _08369_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__xnor2_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _05667_ _05650_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__xor2_1
X_19493_ _02972_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18444_ _02049_ _02051_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__nor2_1
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15656_ _07601_ _08148_ _05198_ _08199_ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__and4_1
X_12868_ _05563_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__nand2_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _07218_ _07323_ _07216_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__a21oi_1
X_18375_ _10094_ _09215_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__nor2_1
X_11819_ rbzero.tex_g1\[51\] rbzero.tex_g1\[50\] _04212_ vssd1 vssd1 vccd1 vccd1 _04596_
+ sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15587_ _07568_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__inv_2
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ rbzero.wall_tracer.mapY\[7\] _05397_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_
+ sky130_fd_sc_hd__o21a_1
X_17326_ _09889_ _09893_ _09894_ _09780_ vssd1 vssd1 vccd1 vccd1 _09895_ sky130_fd_sc_hd__a31o_1
X_14538_ _07233_ _07249_ _07247_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__a21oi_1
XFILLER_202_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17257_ _09830_ _09831_ _09832_ vssd1 vssd1 vccd1 vccd1 _09833_ sky130_fd_sc_hd__and3_1
X_14469_ _07131_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__nor2_1
XFILLER_146_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16208_ _08847_ _08852_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__nand2_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17188_ _09773_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16139_ _08519_ _08674_ _08112_ _08377_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__o22a_1
XFILLER_170_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19829_ _03139_ _03147_ _03149_ _02765_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__o211a_1
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21653_ clknet_leaf_46_i_clk _01422_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20604_ _03466_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21584_ net505 _01353_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20535_ rbzero.traced_texa\[7\] rbzero.texV\[7\] _03422_ vssd1 vssd1 vccd1 vccd1
+ _03427_ sky130_fd_sc_hd__a21o_1
XFILLER_166_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_78 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_78/HI o_rgb[8] sky130_fd_sc_hd__conb_1
XFILLER_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_89 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_89/HI o_rgb[21] sky130_fd_sc_hd__conb_1
XFILLER_119_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20466_ _03362_ _03364_ _03363_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__o21bai_1
XFILLER_174_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21018_ clknet_leaf_69_i_clk _00787_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13840_ _05752_ _05921_ _06053_ _05974_ _05989_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a32o_1
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__nand2_1
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ _03839_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15510_ _08043_ _08055_ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__and2b_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12722_ _05423_ _05428_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__or2_2
X_16490_ _07598_ _08230_ _08147_ _08984_ vssd1 vssd1 vccd1 vccd1 _09134_ sky130_fd_sc_hd__or4_1
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _08076_ _08085_ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__or2_1
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _05403_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _04210_ _04377_ _04382_ _04232_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a211o_1
XFILLER_129_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18160_ _01860_ _10238_ _09973_ _01737_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o22ai_1
XFILLER_157_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ _07933_ _07524_ _08016_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__o21ai_1
X_12584_ _05297_ _05337_ _05296_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _03555_ _04037_ vssd1 vssd1 vccd1 vccd1 _09749_ sky130_fd_sc_hd__nor2_1
X_14323_ _05982_ _06658_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__nor2_1
X_11535_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or2b_4
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18091_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__or2_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ _09409_ _09543_ _09681_ vssd1 vssd1 vccd1 vccd1 _09682_ sky130_fd_sc_hd__a21bo_1
X_14254_ _06951_ _06988_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__a21o_1
X_11466_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _04213_ vssd1 vssd1 vccd1 vccd1 _04246_
+ sky130_fd_sc_hd__mux2_1
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13205_ _05941_ _05910_ _05923_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__o21ai_1
X_10417_ _03540_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
X_14185_ _06666_ _06690_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__nor2_1
X_11397_ gpout0.hpos\[9\] _04158_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__o21a_1
XFILLER_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20115__148 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__inv_2
X_13136_ _05791_ _05795_ _05591_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__or3b_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10348_ rbzero.tex_r1\[44\] rbzero.tex_r1\[45\] _03494_ vssd1 vssd1 vccd1 vccd1 _03504_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _02594_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__clkbuf_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13067_ _05591_ _05803_ _05791_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__mux2_1
X_17944_ _01643_ _01644_ _01646_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__nand3_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12018_ rbzero.tex_b1\[47\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04793_
+ sky130_fd_sc_hd__a31o_1
X_17875_ _09249_ _01576_ _01577_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__o21ba_1
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _09082_ _09467_ vssd1 vssd1 vccd1 vccd1 _09468_ sky130_fd_sc_hd__nor2_1
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16757_ _09397_ _09398_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__xnor2_1
X_19545_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] vssd1 vssd1 vccd1
+ vccd1 _03019_ sky130_fd_sc_hd__nor2b_4
XFILLER_111_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13969_ _06613_ _06563_ _06600_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__or3_1
XFILLER_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15708_ _08022_ _08035_ _08046_ _08112_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_1_1__f__03045_ clknet_0__03045_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03045_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_94_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16688_ _09207_ _09330_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__xnor2_4
X_19476_ _02938_ _02956_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__xor2_1
XFILLER_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _07924_ vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__buf_4
X_18427_ _02122_ _02124_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__nand2_1
XFILLER_62_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ _01977_ _01997_ _01975_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17309_ _09879_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18289_ _08802_ _10139_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__nor2_1
XFILLER_147_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21636_ clknet_leaf_37_i_clk _01405_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21567_ net488 _01336_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11320_ _04069_ _04097_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__o21a_1
X_20518_ _03411_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__nand2_1
XFILLER_193_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21498_ net419 _01267_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11251_ rbzero.vga_sync.vsync _03555_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nor2_8
X_20449_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] _03354_ vssd1 vssd1 vccd1 vccd1
+ _03355_ sky130_fd_sc_hd__o21ai_1
XFILLER_118_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11182_ rbzero.map_rom.f3 rbzero.map_rom.f2 rbzero.map_rom.a6 rbzero.map_rom.i_row\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a22o_1
XFILLER_180_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15990_ _07958_ _08041_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__or2_1
XFILLER_125_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14941_ rbzero.wall_tracer.visualWallDist\[5\] _07618_ vssd1 vssd1 vccd1 vccd1 _07637_
+ sky130_fd_sc_hd__or2_1
XFILLER_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17660_ _10215_ _10224_ vssd1 vssd1 vccd1 vccd1 _10225_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14872_ rbzero.wall_tracer.stepDistY\[10\] _07586_ _05188_ vssd1 vssd1 vccd1 vccd1
+ _07587_ sky130_fd_sc_hd__mux2_1
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16611_ _09252_ _09253_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__nand2_1
X_13823_ _06378_ _06558_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__a21o_1
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17591_ _10011_ _10013_ vssd1 vssd1 vccd1 vccd1 _10157_ sky130_fd_sc_hd__or2b_1
XFILLER_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ _09183_ _09185_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__xnor2_2
XFILLER_62_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19330_ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__clkbuf_4
X_13754_ _06483_ _06485_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__nand2_1
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10966_ rbzero.tex_b1\[9\] rbzero.tex_b1\[10\] _03828_ vssd1 vssd1 vccd1 vccd1 _03831_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19261_ _02784_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _05451_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nand2_1
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16473_ _08194_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__buf_4
XFILLER_204_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13685_ _06379_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__nor2_1
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10897_ _03794_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18212_ _01909_ _01910_ _01911_ _05204_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__o31a_1
X_15424_ rbzero.debug_overlay.playerY\[-3\] _07952_ vssd1 vssd1 vccd1 vccd1 _08069_
+ sky130_fd_sc_hd__nand2_1
X_19192_ rbzero.spi_registers.new_sky\[0\] rbzero.spi_registers.got_new_sky _02711_
+ _02741_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a31o_1
X_12636_ rbzero.map_rom.a6 _05374_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__or2_1
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18143_ _10239_ _08423_ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__or3_1
X_15355_ rbzero.debug_overlay.playerX\[-7\] vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__inv_2
XFILLER_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12567_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__or2_1
XFILLER_157_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14306_ _07042_ _06995_ _07039_ _07038_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a31o_1
XFILLER_102_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11518_ _04294_ _04297_ _04210_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__mux2_1
X_18074_ _01773_ _01774_ _01733_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a21oi_1
XFILLER_184_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15286_ _07929_ _07930_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__or2_2
XFILLER_116_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12498_ _05251_ rbzero.wall_tracer.trackDistX\[-2\] _05252_ rbzero.wall_tracer.trackDistX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__o22a_1
XFILLER_176_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17025_ _09661_ _08047_ _09662_ _09664_ vssd1 vssd1 vccd1 vccd1 _09665_ sky130_fd_sc_hd__or4bb_2
X_14237_ _06844_ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__and2_1
X_11449_ _04123_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__buf_4
XFILLER_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14168_ _06903_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__and2b_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _05852_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a21o_1
XFILLER_124_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14099_ _06823_ _06834_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__or2b_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _02618_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17927_ _01622_ _01629_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__xnor2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17858_ _01457_ _01490_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16809_ _09347_ _09450_ vssd1 vssd1 vccd1 vccd1 _09451_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17789_ _10247_ _10250_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__nor2_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19528_ _03003_ _03004_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__nor2_1
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19459_ _02927_ _02938_ _02939_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__nor3_1
XFILLER_210_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21421_ net342 _01190_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21352_ net273 _01121_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21283_ clknet_leaf_42_i_clk _01052_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20250__269 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__inv_2
XFILLER_143_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _03754_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20144__174 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__inv_2
X_20998_ clknet_leaf_52_i_clk _00767_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10751_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__clkbuf_4
XFILLER_198_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ _06200_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ rbzero.tex_g1\[16\] rbzero.tex_g1\[17\] _03680_ vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12421_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__inv_4
X_21619_ clknet_leaf_32_i_clk _01388_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15140_ _07756_ _07789_ _07790_ _07796_ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a31o_1
X_12352_ _04154_ _03477_ _05087_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__mux2_1
XFILLER_194_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11303_ _04079_ _04078_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__nand2_1
X_15071_ _07729_ _07731_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__nand2_1
X_12283_ _04867_ _05027_ _05042_ _05049_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__and4_1
XFILLER_181_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14022_ _06641_ _06642_ _06615_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__a21o_2
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11234_ _04018_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18830_ rbzero.wall_tracer.trackDistY\[4\] _02508_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02509_ sky130_fd_sc_hd__mux2_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _03939_ _03952_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o21a_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15973_ _08615_ _08614_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__and2b_1
X_11096_ rbzero.tex_b0\[12\] rbzero.tex_b0\[11\] _03898_ vssd1 vssd1 vccd1 vccd1 _03899_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18761_ rbzero.wall_tracer.trackDistY\[-5\] _02448_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02449_ sky130_fd_sc_hd__mux2_1
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17712_ _10254_ _10276_ vssd1 vssd1 vccd1 vccd1 _10277_ sky130_fd_sc_hd__xnor2_1
X_14924_ _07621_ _07624_ _07625_ _07620_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__o211a_1
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18692_ _02310_ _02313_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__o21a_1
XFILLER_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ _07433_ _07421_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nand2_1
XFILLER_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17643_ _09249_ _09359_ vssd1 vssd1 vccd1 vccd1 _10208_ sky130_fd_sc_hd__nor2_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ _06522_ _06524_ _06526_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or4_1
X_17574_ _08872_ _08873_ _09991_ _10139_ vssd1 vssd1 vccd1 vccd1 _10140_ sky130_fd_sc_hd__or4_1
X_14786_ _05884_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__nor2_1
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _04250_ vssd1 vssd1 vccd1 vccd1 _04773_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19313_ rbzero.spi_registers.spi_done _03480_ _02563_ vssd1 vssd1 vccd1 vccd1 _02812_
+ sky130_fd_sc_hd__and3_1
X_16525_ _08112_ _08329_ _08419_ vssd1 vssd1 vccd1 vccd1 _09169_ sky130_fd_sc_hd__or3_1
X_13737_ _06473_ _06445_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10949_ rbzero.tex_b1\[17\] rbzero.tex_b1\[18\] _03817_ vssd1 vssd1 vccd1 vccd1 _03822_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ _09009_ _09099_ vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__xnor2_1
X_19244_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_sky\[0\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
X_13668_ _06400_ _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _07903_ rbzero.wall_tracer.stepDistY\[-10\] vssd1 vssd1 vccd1 vccd1 _08052_
+ sky130_fd_sc_hd__nand2_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19175_ rbzero.spi_registers.got_new_leak _02708_ vssd1 vssd1 vccd1 vccd1 _02731_
+ sky130_fd_sc_hd__and2_1
X_12619_ _05331_ _05335_ _05340_ _05370_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__o41ai_4
X_16387_ _08331_ _08420_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__nand2_1
X_13599_ _06302_ _06329_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18126_ _08275_ _09165_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__nor2_1
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ _07982_ rbzero.debug_overlay.playerY\[-8\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _07983_ sky130_fd_sc_hd__mux2_1
X_18057_ _10110_ _09991_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__nor2_1
X_15269_ rbzero.debug_overlay.playerX\[-5\] _07898_ vssd1 vssd1 vccd1 vccd1 _07914_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ _09387_ _09390_ _09505_ vssd1 vssd1 vccd1 vccd1 _09648_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18959_ _02609_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19605__59 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20921_ clknet_leaf_69_i_clk _00690_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20852_ clknet_leaf_92_i_clk _00621_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20783_ clknet_leaf_21_i_clk _00552_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21404_ net325 _01173_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21335_ net256 _01104_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21266_ clknet_leaf_62_i_clk _01035_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21197_ clknet_leaf_64_i_clk _00966_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12970_ _05593_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11921_ _04695_ _04696_ _04139_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__mux2_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _07106_ _07107_ _07041_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__and3_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ rbzero.tex_g1\[14\] _04272_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__and2_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _03745_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14571_ _07306_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__nand2_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ rbzero.tex_g0\[56\] _04350_ _04224_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a21o_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16310_ _08951_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__a21oi_4
X_13522_ _06080_ _06134_ _05921_ _05989_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__and4bb_1
XFILLER_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17290_ _09862_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__clkbuf_1
X_10734_ rbzero.tex_g0\[56\] rbzero.tex_g0\[55\] _03706_ vssd1 vssd1 vccd1 vccd1 _03709_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _08884_ _08865_ _08876_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__nand3_1
X_13453_ _06077_ _06088_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__and2b_1
XFILLER_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ rbzero.tex_g1\[24\] rbzero.tex_g1\[25\] _03669_ vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12404_ _05141_ _05166_ _05168_ _05170_ _05153_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__o221a_1
XFILLER_139_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16172_ _08674_ _08112_ _08747_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__nor3_1
X_13384_ _06112_ _06118_ _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a21bo_1
XFILLER_182_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10596_ _03636_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15123_ _07772_ _07773_ _07780_ _07676_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__a2bb2o_1
X_12335_ _05083_ _05082_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__and2b_1
XFILLER_115_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15054_ _07676_ _07708_ _07709_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__a31o_1
X_19931_ rbzero.debug_overlay.playerY\[2\] _03198_ _03226_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _01000_ sky130_fd_sc_hd__o211a_1
X_12266_ _05032_ _05033_ _05034_ _05024_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__o31a_1
XFILLER_99_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ _06659_ _06741_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__xnor2_1
X_11217_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__buf_2
X_19862_ _03141_ _03171_ _03172_ _03173_ _03155_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__o311a_1
Xoutput70 net122 vssd1 vssd1 vccd1 vccd1 o_tex_sclk sky130_fd_sc_hd__clkbuf_1
X_12197_ _04966_ _04666_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__nand2_1
XFILLER_123_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_150_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18813_ _02487_ _02489_ _02492_ _02493_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a211oi_1
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11148_ rbzero.debug_overlay.playerY\[2\] _03934_ _03936_ rbzero.debug_overlay.playerX\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__a2bb2o_1
X_19793_ _03125_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18744_ rbzero.wall_tracer.trackDistY\[-7\] _02433_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02434_ sky130_fd_sc_hd__mux2_1
X_15956_ _08588_ _08600_ vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__xor2_2
X_11079_ rbzero.tex_b0\[20\] rbzero.tex_b0\[19\] _03887_ vssd1 vssd1 vccd1 vccd1 _03890_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03293_ clknet_0__03293_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03293_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14907_ rbzero.wall_tracer.visualWallDist\[-5\] _07595_ vssd1 vssd1 vccd1 vccd1 _07613_
+ sky130_fd_sc_hd__or2_1
X_15887_ _08484_ _08479_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18675_ _02259_ _02267_ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a21oi_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17626_ _10189_ _10190_ vssd1 vssd1 vccd1 vccd1 _10191_ sky130_fd_sc_hd__nand2_1
X_14838_ _07561_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14769_ rbzero.wall_tracer.stepDistY\[-9\] _07502_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07503_ sky130_fd_sc_hd__mux2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17557_ _10001_ _10000_ vssd1 vssd1 vccd1 vccd1 _10123_ sky130_fd_sc_hd__or2b_1
XFILLER_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16508_ _09149_ _09151_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__xnor2_1
X_17488_ _09368_ _09483_ _09910_ vssd1 vssd1 vccd1 vccd1 _10054_ sky130_fd_sc_hd__or3_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19227_ _02721_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__clkbuf_4
X_16439_ _09080_ _09082_ _05194_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__a21o_1
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19158_ rbzero.othery\[0\] _02710_ _02719_ _02714_ vssd1 vssd1 vccd1 vccd1 _00734_
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18109_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
X_19089_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.mosi _02677_ vssd1
+ vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
X_21120_ net210 _00889_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21051_ clknet_leaf_3_i_clk _00820_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20002_ rbzero.pov.ready_buffer\[6\] _03239_ _03242_ _04471_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01043_ sky130_fd_sc_hd__o221a_1
XFILLER_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ clknet_leaf_80_i_clk _00673_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ clknet_leaf_28_i_clk _00604_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20766_ clknet_leaf_33_i_clk _00535_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20697_ clknet_leaf_5_i_clk _00481_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10450_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _03558_ vssd1 vssd1 vccd1 vccd1 _03560_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20256__275 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__inv_2
XFILLER_109_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10381_ _03521_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
X_12120_ gpout0.vpos\[1\] vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21318_ net239 _01087_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12051_ _04814_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__nor2_1
X_21249_ clknet_leaf_80_i_clk _01018_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_77_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _03849_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15810_ _08451_ _08453_ _08454_ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__a21oi_2
X_16790_ _07575_ _07579_ _08983_ _07582_ vssd1 vssd1 vccd1 vccd1 _09432_ sky130_fd_sc_hd__o31a_1
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15741_ _08384_ _08385_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__nand2_1
X_12953_ _05632_ _05637_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__or2b_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11904_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _04290_ vssd1 vssd1 vccd1 vccd1 _04680_
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15672_ _08314_ _08315_ _08316_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__a21bo_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _02149_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__xnor2_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12884_ rbzero.wall_tracer.visualWallDist\[1\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05621_ sky130_fd_sc_hd__a21o_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _07358_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__xnor2_2
X_17411_ _08872_ _09977_ _09700_ vssd1 vssd1 vccd1 vccd1 _09978_ sky130_fd_sc_hd__or3_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _08257_ _08423_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__nor2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ rbzero.tex_g1\[41\] rbzero.tex_g1\[40\] _04350_ vssd1 vssd1 vccd1 vccd1 _04612_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _09656_ _09617_ vssd1 vssd1 vccd1 vccd1 _09909_ sky130_fd_sc_hd__or2b_1
XFILLER_187_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14554_ _07289_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__nand2_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _04129_ vssd1 vssd1 vccd1 vccd1 _04544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ _05974_ _06240_ _06161_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__or3_1
X_17273_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09847_ sky130_fd_sc_hd__nand2_1
X_10717_ net47 rbzero.tex_g0\[63\] _03624_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__mux2_1
X_14485_ _07172_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11697_ rbzero.debug_overlay.vplaneY\[-8\] _04466_ _04458_ rbzero.debug_overlay.vplaneY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a22o_1
X_19012_ rbzero.pov.spi_buffer\[38\] rbzero.pov.ready_buffer\[38\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
X_16224_ _08170_ _08572_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__or2_1
X_13436_ _06082_ _06087_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nand2_1
X_10648_ rbzero.tex_g1\[32\] rbzero.tex_g1\[33\] _03658_ vssd1 vssd1 vccd1 vccd1 _03664_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16155_ _08778_ _08798_ _08799_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__a21oi_1
X_13367_ _06100_ _06101_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__xor2_1
XFILLER_177_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10579_ _03627_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15106_ _07751_ _07754_ _07763_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__and3_1
X_12318_ _05081_ _05084_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__and3_1
XFILLER_114_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16086_ _08729_ _08730_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__xnor2_1
X_13298_ _06032_ _06033_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__a21o_1
XFILLER_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15037_ _07697_ _07698_ _07699_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__o21ai_1
X_19914_ rbzero.debug_overlay.playerY\[-2\] _03198_ _03213_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00996_ sky130_fd_sc_hd__o211a_1
X_12249_ net18 net19 _05002_ _05009_ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__o311a_2
XFILLER_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19845_ _08067_ _03143_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nand2_1
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19776_ rbzero.pov.spi_buffer\[61\] rbzero.pov.spi_buffer\[62\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03117_ sky130_fd_sc_hd__mux2_1
X_16988_ _08821_ _09028_ _08425_ _09243_ vssd1 vssd1 vccd1 vccd1 _09628_ sky130_fd_sc_hd__o22a_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18727_ _09863_ _02417_ _02418_ _09835_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__o31ai_1
X_15939_ _08566_ _08583_ _08492_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__a21oi_4
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19595__50 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
X_18658_ _02263_ _02264_ _02261_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a21boi_1
XFILLER_58_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17609_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _10175_ sky130_fd_sc_hd__nand2_1
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18589_ _02254_ _02285_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__xor2_1
XFILLER_149_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20620_ clknet_leaf_71_i_clk _00404_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.a6 sky130_fd_sc_hd__dfxtp_2
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20551_ rbzero.traced_texa\[11\] rbzero.texV\[11\] vssd1 vssd1 vccd1 vccd1 _03440_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_165_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20482_ _03272_ _03381_ _03382_ _03250_ rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1
+ _01395_ sky130_fd_sc_hd__a32o_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21103_ net193 _00872_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21034_ clknet_leaf_51_i_clk _00803_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vshift
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11620_ _04379_ _04396_ _04397_ _04398_ _04209_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__o221a_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20818_ clknet_leaf_7_i_clk _00587_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ rbzero.tex_r1\[15\] _04327_ _04328_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_
+ sky130_fd_sc_hd__a31o_1
XFILLER_196_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20749_ clknet_leaf_35_i_clk _00518_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10502_ rbzero.tex_r0\[38\] rbzero.tex_r0\[37\] _03580_ vssd1 vssd1 vccd1 vccd1 _03587_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14270_ _06762_ _06765_ _06764_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a21bo_1
XFILLER_109_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11482_ _04211_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__buf_6
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03296_ clknet_0__03296_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03296_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ _05688_ _05792_ _05957_ _05778_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a211o_1
X_10433_ _03548_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13152_ _05856_ _05877_ _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a21o_2
XFILLER_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10364_ _03512_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12103_ _04813_ _04811_ _04006_ _03475_ net2 net3 vssd1 vssd1 vccd1 vccd1 _04875_
+ sky130_fd_sc_hd__mux4_1
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13083_ _05797_ _05809_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__nand2_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17960_ _01660_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12034_ _04808_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_4
X_16911_ _09551_ vssd1 vssd1 vccd1 vccd1 _09552_ sky130_fd_sc_hd__buf_2
X_17891_ _08259_ _08202_ _08157_ _08149_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__or4_1
XFILLER_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16842_ _09482_ vssd1 vssd1 vccd1 vccd1 _09483_ sky130_fd_sc_hd__buf_2
XFILLER_66_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19561_ rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\] _03028_ vssd1 vssd1
+ vccd1 vccd1 _03031_ sky130_fd_sc_hd__and3_1
X_13985_ _06719_ _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__and2_1
XFILLER_168_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16773_ _09407_ _09414_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__xor2_2
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18512_ _02208_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__nand2_1
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15724_ _08367_ _08368_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__nand2_1
X_12936_ _05657_ _05658_ _05663_ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or4_2
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ rbzero.wall_tracer.rayAddendY\[6\] _02971_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _02972_ sky130_fd_sc_hd__mux2_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _02139_ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__nor2b_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12867_ rbzero.wall_tracer.visualWallDist\[4\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05604_ sky130_fd_sc_hd__a21o_1
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ rbzero.wall_tracer.visualWallDist\[-11\] _08148_ _05198_ _08254_ vssd1 vssd1
+ vccd1 vccd1 _08300_ sky130_fd_sc_hd__and4_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _07329_ _07330_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__nand3b_2
X_11818_ rbzero.tex_g1\[49\] rbzero.tex_g1\[48\] _04212_ vssd1 vssd1 vccd1 vccd1 _04595_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18374_ _01939_ _02071_ _02072_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a21o_1
X_15586_ _08230_ rbzero.wall_tracer.stepDistY\[5\] vssd1 vssd1 vccd1 vccd1 _08231_
+ sky130_fd_sc_hd__nand2_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ rbzero.wall_tracer.mapY\[6\] _05397_ _05538_ vssd1 vssd1 vccd1 vccd1 _05540_
+ sky130_fd_sc_hd__a21bo_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _07197_ _07195_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__xor2_1
X_17325_ _09890_ _09891_ _09892_ vssd1 vssd1 vccd1 vccd1 _09894_ sky130_fd_sc_hd__o21ai_1
X_11749_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _04271_ vssd1 vssd1 vccd1 vccd1 _04527_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14468_ _06724_ _06760_ _07117_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__or3_1
X_17256_ _09823_ _09821_ _09822_ vssd1 vssd1 vccd1 vccd1 _09832_ sky130_fd_sc_hd__a21bo_1
XFILLER_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13419_ _06154_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__or2_1
XFILLER_190_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16207_ _08840_ _08846_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__or2_1
XFILLER_162_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17187_ rbzero.wall_tracer.wall\[1\] rbzero.row_render.wall\[1\] _07830_ vssd1 vssd1
+ vccd1 vccd1 _09773_ sky130_fd_sc_hd__mux2_1
XFILLER_190_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ _06698_ _06740_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__nor2_1
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16138_ _08748_ _08745_ _08746_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16069_ _08697_ _08712_ _08713_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19828_ _03148_ _03143_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__nand2_1
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19759_ rbzero.pov.spi_buffer\[53\] rbzero.pov.spi_buffer\[54\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21652_ clknet_leaf_43_i_clk _01421_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20603_ _02721_ _03464_ _03465_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__and3_1
X_21583_ net504 _01352_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20534_ _03424_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and2b_1
XFILLER_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_79 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_79/HI o_rgb[9] sky130_fd_sc_hd__conb_1
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20465_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03368_
+ sky130_fd_sc_hd__nand2_1
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20368__376 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__inv_2
X_21017_ clknet_leaf_69_i_clk _00786_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20067__104 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__inv_2
XFILLER_134_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13770_ _06488_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__and2_1
X_10982_ rbzero.tex_b1\[1\] rbzero.tex_b1\[2\] _03482_ vssd1 vssd1 vccd1 vccd1 _03839_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12721_ _05430_ _05433_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__xor2_4
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19574__31 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15440_ _08084_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__or3_1
Xclkbuf_2_0_0_i_clk clknet_1_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ _05402_ rbzero.map_rom.i_row\[4\] _05283_ vssd1 vssd1 vccd1 vccd1 _05403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _04378_ _04380_ _04381_ _04219_ _04230_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__o221a_1
XFILLER_141_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15371_ _07933_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__nand2_1
XFILLER_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _05301_ _05336_ _05305_ _05309_ _05299_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o311ai_4
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_55_i_clk clknet_opt_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14322_ _07058_ _07001_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__xnor2_1
X_17110_ _03474_ _09748_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__nor2_1
X_11534_ _04047_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__inv_2
X_18090_ _09807_ _01790_ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__or3_1
XFILLER_156_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ _09114_ _09126_ _09544_ vssd1 vssd1 vccd1 vccd1 _09681_ sky130_fd_sc_hd__or3_1
X_14253_ _06986_ _06987_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__and2b_1
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _04213_ vssd1 vssd1 vccd1 vccd1 _04245_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _05889_ _05900_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nand2_1
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ rbzero.tex_r1\[12\] rbzero.tex_r1\[13\] _03538_ vssd1 vssd1 vccd1 vccd1 _03540_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14184_ _06919_ _06920_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__nand2_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11396_ rbzero.row_render.size\[9\] _04155_ rbzero.row_render.size\[10\] vssd1 vssd1
+ vccd1 vccd1 _04176_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13135_ _05705_ _05707_ _05791_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10347_ _03503_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _02626_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _05593_ _05706_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__xor2_2
X_17943_ _10271_ _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12017_ rbzero.tex_b1\[46\] _04272_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__and2_1
XFILLER_94_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17874_ _09391_ _09480_ _09484_ _09249_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__o22a_1
XFILLER_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16825_ _09465_ _09466_ vssd1 vssd1 vccd1 vccd1 _09467_ sky130_fd_sc_hd__nor2_1
XFILLER_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19544_ _03914_ _03018_ _03009_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16756_ _08282_ _09103_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__or2_1
XFILLER_98_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _06704_ _06658_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03044_ clknet_0__03044_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03044_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15707_ _08022_ _08034_ _08045_ _08112_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__or4_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _05650_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nor2_1
X_19475_ _02904_ _04471_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__xor2_1
X_13899_ _06248_ _06581_ _06583_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a21o_1
X_16687_ _09328_ _09329_ vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__and2_2
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18426_ _02122_ _02124_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__or2_2
X_15638_ _07913_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__buf_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18357_ _02033_ _02055_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _08002_ _08207_ _08210_ _08213_ _07945_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__a221o_1
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17308_ rbzero.wall_tracer.trackDistX\[-4\] _09878_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09879_ sky130_fd_sc_hd__mux2_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18288_ _09668_ _09991_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__nor2_1
XFILLER_175_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17239_ _05413_ vssd1 vssd1 vccd1 vccd1 _09817_ sky130_fd_sc_hd__clkbuf_4
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21635_ clknet_leaf_37_i_clk _01404_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21566_ net487 _01335_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20517_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__nand2_1
XFILLER_197_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21497_ net418 _01266_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11250_ rbzero.wall_tracer.state\[0\] vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__inv_2
XFILLER_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20448_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] _03349_ vssd1 vssd1 vccd1 vccd1
+ _03354_ sky130_fd_sc_hd__a21o_1
XFILLER_134_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11181_ rbzero.wall_tracer.state\[1\] _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__nand2_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14940_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.trackDistX\[5\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__mux2_1
XFILLER_75_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14871_ _07468_ _07585_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__or2b_2
XFILLER_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16610_ _08383_ _08111_ _08570_ _08282_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__o22ai_1
X_13822_ _06278_ _06334_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17590_ _10088_ _10155_ vssd1 vssd1 vccd1 vccd1 _10156_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13753_ _06467_ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__and2b_1
X_16541_ _09025_ _09049_ _09184_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__a21oi_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10965_ _03830_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__nand2_1
X_19260_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_floor\[0\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ _06391_ _06419_ _06420_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a21oi_2
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16472_ _08962_ _08963_ _09115_ vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__a21bo_1
X_10896_ rbzero.tex_b1\[42\] rbzero.tex_b1\[43\] _03784_ vssd1 vssd1 vccd1 vccd1 _03794_
+ sky130_fd_sc_hd__mux2_1
XFILLER_176_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18211_ _01909_ _01910_ _01911_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12635_ _05387_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__clkbuf_1
X_15423_ _08066_ _08067_ _05495_ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__mux2_1
X_19191_ _03555_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__buf_4
X_20121__153 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__inv_2
XFILLER_169_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18142_ _01841_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__xnor2_1
X_15354_ _07897_ _07998_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__nand2_1
XFILLER_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12566_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__xor2_1
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11517_ _04295_ _04296_ _04247_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
X_14305_ _06882_ _07034_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__nand2_1
XFILLER_157_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15285_ _05197_ rbzero.wall_tracer.stepDistX\[-4\] vssd1 vssd1 vccd1 vccd1 _07930_
+ sky130_fd_sc_hd__nor2_1
X_18073_ _01733_ _01773_ _01774_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__and3_1
X_12497_ rbzero.wall_tracer.trackDistY\[-3\] vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__inv_2
XFILLER_141_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14236_ _06964_ _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17024_ _08383_ _09103_ _09663_ vssd1 vssd1 vccd1 vccd1 _09664_ sky130_fd_sc_hd__or3_1
X_11448_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _04214_ vssd1 vssd1 vccd1 vccd1 _04228_
+ sky130_fd_sc_hd__mux2_1
XFILLER_172_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14167_ _06741_ _06888_ _06889_ _06891_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a22o_1
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] vssd1 vssd1 vccd1
+ vccd1 _04159_ sky130_fd_sc_hd__xnor2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13118_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__buf_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _06823_ _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__xnor2_1
X_18975_ rbzero.pov.spi_buffer\[20\] rbzero.pov.ready_buffer\[20\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _05725_ _05657_ _05658_ _05663_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__or4_1
XFILLER_117_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17926_ _01626_ _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__xor2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17857_ _10189_ _01452_ _01451_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__o21bai_1
XFILLER_67_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20396__21 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16808_ _09448_ _09449_ vssd1 vssd1 vccd1 vccd1 _09450_ sky130_fd_sc_hd__xor2_1
X_17788_ _01455_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19527_ _03002_ _03000_ _03001_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__and3_1
X_16739_ _09379_ _09380_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__nand2_1
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20204__228 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__inv_2
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19458_ _02938_ _02939_ _02927_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o21a_1
XFILLER_90_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18409_ _01936_ _01937_ _01935_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__o21a_1
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19389_ _02865_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__xnor2_1
XFILLER_194_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21420_ net341 _01189_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20096__130 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__inv_2
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21351_ net272 _01120_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21282_ clknet_leaf_42_i_clk _01051_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20997_ clknet_leaf_52_i_clk _00766_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _03556_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__buf_4
XFILLER_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20179__205 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__inv_2
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10681_ _03681_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12420_ _05138_ _05140_ _05178_ _05186_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__o2bb2a_2
X_21618_ clknet_leaf_32_i_clk _01387_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12351_ net28 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__or2_1
XFILLER_51_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21549_ net470 _01318_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11302_ _04077_ _04080_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15070_ _07730_ rbzero.wall_tracer.rayAddendX\[-1\] vssd1 vssd1 vccd1 vccd1 _07731_
+ sky130_fd_sc_hd__nand2_1
X_12282_ _05042_ _05045_ _05048_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a211o_1
XFILLER_119_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ _06615_ _06641_ _06642_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__nand3_4
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ _03969_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__or2_1
XFILLER_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ rbzero.wall_tracer.visualWallDist\[11\] vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__inv_2
XFILLER_150_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18760_ _09863_ _02446_ _02447_ _09869_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o31ai_1
X_15972_ _08550_ _08616_ vssd1 vssd1 vccd1 vccd1 _08617_ sky130_fd_sc_hd__xor2_2
X_11095_ _03556_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17711_ _10273_ _10275_ vssd1 vssd1 vccd1 vccd1 _10276_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14923_ rbzero.wall_tracer.visualWallDist\[-1\] _07618_ vssd1 vssd1 vccd1 vccd1 _07625_
+ sky130_fd_sc_hd__or2_1
X_18691_ _02382_ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__xor2_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17642_ _09391_ _10205_ _10206_ vssd1 vssd1 vccd1 vccd1 _10207_ sky130_fd_sc_hd__o21ba_1
XFILLER_91_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14854_ _07572_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__clkbuf_1
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13805_ _05825_ _06031_ _06527_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__o31a_1
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17573_ _10138_ _09565_ _05198_ vssd1 vssd1 vccd1 vccd1 _10139_ sky130_fd_sc_hd__mux2_4
X_14785_ _07490_ _07493_ _05952_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__mux2_1
X_11997_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _04250_ vssd1 vssd1 vccd1 vccd1 _04772_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19312_ rbzero.spi_registers.got_new_other _02730_ _02728_ _02801_ vssd1 vssd1 vccd1
+ vccd1 _00796_ sky130_fd_sc_hd__a31o_1
XFILLER_205_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16524_ _09003_ _09006_ vssd1 vssd1 vccd1 vccd1 _09168_ sky130_fd_sc_hd__nand2_1
XFILLER_204_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13736_ _06045_ _06016_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nor2_1
X_10948_ _03821_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19243_ _02773_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16455_ _07977_ _08109_ vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__nor2_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13667_ _06356_ _06401_ _06402_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__o22a_1
XFILLER_143_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10879_ _03785_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ rbzero.wall_tracer.side _08049_ _08050_ rbzero.wall_tracer.state\[3\] vssd1
+ vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__o211a_1
X_12618_ _05327_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nand2_2
X_19174_ rbzero.spi_registers.new_vinf _02726_ _02728_ _02729_ _02730_ vssd1 vssd1
+ vccd1 vccd1 _00739_ sky130_fd_sc_hd__o311a_1
X_13598_ _06278_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__nand2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _08416_ _08420_ _08426_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__a21bo_1
XFILLER_129_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18125_ _01824_ _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__xnor2_1
X_12549_ _05301_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__nor2_1
X_15337_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__xor2_1
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18056_ _08895_ _08767_ _01524_ _10139_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__or4_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _03953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__buf_2
XFILLER_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17007_ _09639_ _09646_ vssd1 vssd1 vccd1 vccd1 _09647_ sky130_fd_sc_hd__xnor2_1
X_14219_ _06924_ _06930_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__or2b_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15199_ _07835_ _07838_ _07836_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__a21boi_1
XFILLER_141_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18958_ rbzero.pov.spi_buffer\[12\] rbzero.pov.ready_buffer\[12\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17909_ _01507_ _01509_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__nor2_1
X_18889_ rbzero.spi_registers.spi_counter\[3\] vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__inv_2
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20920_ clknet_leaf_70_i_clk _00689_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20128__159 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__inv_2
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20851_ clknet_leaf_93_i_clk _00620_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20782_ clknet_leaf_22_i_clk _00551_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21403_ net324 _01172_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21334_ net255 _01103_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21265_ clknet_leaf_82_i_clk _01034_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20216_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__buf_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21196_ clknet_leaf_64_i_clk _00965_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _04271_ vssd1 vssd1 vccd1 vccd1 _04696_
+ sky130_fd_sc_hd__mux2_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _04610_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__nor2_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ rbzero.tex_g0\[24\] rbzero.tex_g0\[23\] _03740_ vssd1 vssd1 vccd1 vccd1 _03745_
+ sky130_fd_sc_hd__mux2_1
X_14570_ _07295_ _07300_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__xor2_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11782_ rbzero.tex_g0\[57\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__and3_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13521_ _05990_ _06067_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__or2_1
X_20390__16 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
XFILLER_159_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _03708_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13452_ _06152_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16240_ _08865_ _08876_ _08884_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__a21o_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10664_ _03672_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ _05149_ _05169_ _05145_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a21o_1
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13383_ _06045_ _06114_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__or3_1
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16171_ _08594_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__clkbuf_4
XFILLER_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ rbzero.tex_g1\[57\] rbzero.tex_g1\[58\] _03635_ vssd1 vssd1 vccd1 vccd1 _03636_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ net31 _05099_ _05101_ _04867_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__or4b_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15122_ _07778_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__xor2_1
XFILLER_181_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15053_ _07676_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__nor2_1
X_19930_ rbzero.pov.ready_buffer\[55\] _03141_ _03192_ _03225_ vssd1 vssd1 vccd1 vccd1
+ _03226_ sky130_fd_sc_hd__a211o_1
X_12265_ net24 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__inv_2
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20233__254 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__inv_2
XFILLER_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _06704_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__nor2_1
X_11216_ _04001_ _04002_ _04003_ _03914_ rbzero.wall_tracer.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _00011_ sky130_fd_sc_hd__a311o_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19861_ rbzero.pov.ready_buffer\[69\] _03145_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__or2_1
X_12196_ _04961_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__clkbuf_4
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 o_reset sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 o_vsync sky130_fd_sc_hd__buf_2
X_18812_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__nor2_1
XFILLER_110_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11147_ rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__clkinv_2
XFILLER_150_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19792_ rbzero.pov.spi_buffer\[69\] rbzero.pov.spi_buffer\[70\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XFILLER_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ _02431_ _02432_ _09851_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _03889_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__clkbuf_1
X_15955_ _08589_ _08598_ _08599_ vssd1 vssd1 vccd1 vccd1 _08600_ sky130_fd_sc_hd__a21oi_2
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03292_ clknet_0__03292_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03292_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14906_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.trackDistX\[-5\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__mux2_1
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18674_ _02265_ _02266_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__and2b_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _08514_ _08530_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__xor2_2
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _10064_ _10067_ _10188_ vssd1 vssd1 vccd1 vccd1 _10190_ sky130_fd_sc_hd__nand3_1
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14837_ rbzero.wall_tracer.stepDistY\[1\] _07560_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07561_ sky130_fd_sc_hd__mux2_1
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17556_ _10112_ _10121_ vssd1 vssd1 vccd1 vccd1 _10122_ sky130_fd_sc_hd__xnor2_2
X_14768_ _07487_ _07455_ _07488_ _07501_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a211o_1
XFILLER_211_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16507_ _08970_ _08994_ _09150_ vssd1 vssd1 vccd1 vccd1 _09151_ sky130_fd_sc_hd__a21bo_1
X_13719_ _06454_ _06439_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__or2b_1
XFILLER_177_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17487_ _09368_ _09480_ _09483_ _08329_ vssd1 vssd1 vccd1 vccd1 _10053_ sky130_fd_sc_hd__o22ai_1
XFILLER_189_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14699_ _05892_ _07395_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__nand2_1
XFILLER_147_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19226_ rbzero.spi_registers.new_vshift\[0\] _02763_ vssd1 vssd1 vccd1 vccd1 _02764_
+ sky130_fd_sc_hd__or2_1
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16438_ _09080_ _09082_ vssd1 vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__nor2_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19157_ rbzero.spi_registers.new_other\[0\] _02712_ vssd1 vssd1 vccd1 vccd1 _02719_
+ sky130_fd_sc_hd__or2_1
X_16369_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__nand2_1
XFILLER_30_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18108_ _01808_ _01704_ _01702_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19088_ _02676_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__clkbuf_4
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ _01738_ _01740_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nand2_1
XFILLER_172_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21050_ clknet_leaf_2_i_clk _00819_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20001_ rbzero.pov.ready_buffer\[5\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-4\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__a221o_1
XFILLER_119_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ clknet_leaf_81_i_clk _00672_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20834_ clknet_leaf_27_i_clk _00603_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20765_ clknet_leaf_32_i_clk _00534_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20696_ clknet_leaf_6_i_clk _00480_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ rbzero.tex_r1\[29\] rbzero.tex_r1\[30\] _03516_ vssd1 vssd1 vccd1 vccd1 _03521_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21317_ net238 _01086_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ rbzero.row_render.texu\[1\] rbzero.row_render.texu\[0\] _03473_ vssd1 vssd1
+ vccd1 vccd1 _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_137_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21248_ clknet_leaf_80_i_clk _01017_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11001_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _03843_ vssd1 vssd1 vccd1 vccd1 _03849_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21179_ clknet_leaf_74_i_clk _00948_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04835_ clknet_0__04835_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04835_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _07977_ _08276_ _07981_ _07989_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__or4_1
X_12952_ _05638_ _05649_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__or3_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ rbzero.tex_b0\[2\] _04262_ _04126_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a21o_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _07913_ _07924_ _07995_ _07932_ vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__or4_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _04030_ _05332_ _05341_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__and3_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _09976_ vssd1 vssd1 vccd1 vccd1 _09977_ sky130_fd_sc_hd__clkbuf_4
X_14622_ _07304_ _07308_ _07315_ _07302_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__a31o_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _02087_ _02088_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nand2_1
XFILLER_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ rbzero.tex_g1\[43\] rbzero.tex_g1\[42\] _04350_ vssd1 vssd1 vccd1 vccd1 _04611_
+ sky130_fd_sc_hd__mux2_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _09609_ _09612_ _09907_ vssd1 vssd1 vccd1 vccd1 _09908_ sky130_fd_sc_hd__a21o_2
XFILLER_92_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14553_ _07287_ _07288_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__xor2_1
X_11765_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _04129_ vssd1 vssd1 vccd1 vccd1 _04543_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _06239_ _06240_ _06202_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__o21bai_1
XFILLER_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ _03699_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__clkbuf_1
X_17272_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09846_ sky130_fd_sc_hd__or2_1
XFILLER_105_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14484_ _07176_ _07178_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__xor2_1
X_11696_ _04420_ _04447_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__and2_2
XFILLER_186_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19011_ _02636_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16223_ _08180_ _08491_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__or2_1
X_13435_ _06170_ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__xor2_1
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _03663_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13366_ _05939_ _06016_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nor2_1
XFILLER_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16154_ _08779_ _08797_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__nor2_1
X_10578_ rbzero.tex_r0\[2\] rbzero.tex_r0\[1\] _03624_ vssd1 vssd1 vccd1 vccd1 _03627_
+ sky130_fd_sc_hd__mux2_1
X_15105_ _07751_ _07754_ _07763_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__a21oi_1
X_12317_ net29 net28 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nor2_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13297_ _05988_ _05980_ _05991_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a21oi_1
XFILLER_182_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16085_ _08124_ _08490_ _07924_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12248_ _04972_ _05011_ _05017_ net18 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a211o_1
X_15036_ _07697_ _07698_ _07699_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__or3_1
X_19913_ _08080_ _02823_ _03197_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__o211ai_1
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19844_ rbzero.pov.ready_buffer\[65\] _08066_ _03146_ vssd1 vssd1 vccd1 vccd1 _03160_
+ sky130_fd_sc_hd__mux2_1
X_12179_ gpout0.vpos\[4\] gpout0.vpos\[5\] _04891_ gpout0.vpos\[9\] net8 net10 vssd1
+ vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__mux4_1
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19775_ _03116_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16987_ _08823_ _09164_ vssd1 vssd1 vccd1 vccd1 _09627_ sky130_fd_sc_hd__nor2_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18726_ _02414_ _02415_ _02416_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a21oi_1
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15938_ _08568_ _08582_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__or2b_1
XFILLER_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18657_ _02144_ _02246_ _02352_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15869_ _08451_ _08453_ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__xnor2_2
XFILLER_37_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17608_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _10174_ sky130_fd_sc_hd__or2_1
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18588_ _02268_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__xor2_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _08178_ _09674_ _09965_ _10104_ vssd1 vssd1 vccd1 vccd1 _10105_ sky130_fd_sc_hd__o31a_1
XFILLER_178_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20550_ _09750_ _03438_ _03439_ _03250_ rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1
+ _01406_ sky130_fd_sc_hd__a32o_1
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19209_ _09753_ _02752_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__and2_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20481_ _03378_ _03379_ _03373_ _03377_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a211o_1
XFILLER_146_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21102_ net192 _00871_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21033_ clknet_leaf_51_i_clk _00802_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20262__280 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__inv_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20817_ clknet_leaf_7_i_clk _00586_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11550_ _04126_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__buf_4
X_20748_ clknet_leaf_39_i_clk _00517_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10501_ _03586_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _04213_ vssd1 vssd1 vccd1 vccd1 _04261_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20679_ clknet_leaf_2_i_clk _00463_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[8\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _05640_ _05792_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__03295_ clknet_0__03295_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03295_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10432_ rbzero.tex_r1\[4\] rbzero.tex_r1\[5\] _03538_ vssd1 vssd1 vccd1 vccd1 _03548_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13151_ _05700_ _05879_ _05881_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a211oi_4
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ rbzero.tex_r1\[37\] rbzero.tex_r1\[38\] _03505_ vssd1 vssd1 vccd1 vccd1 _03512_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ net5 net4 _04873_ net6 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a31o_1
XFILLER_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _05816_ _05818_ _05806_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__mux2_1
XFILLER_152_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _04314_ _04807_ _04521_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__o21a_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16910_ _08237_ _09279_ vssd1 vssd1 vccd1 vccd1 _09551_ sky130_fd_sc_hd__and2_1
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17890_ _01499_ _01501_ _01497_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a21bo_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16841_ _05211_ _09481_ vssd1 vssd1 vccd1 vccd1 _09482_ sky130_fd_sc_hd__or2_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19560_ rbzero.pov.spi_counter\[3\] _03028_ _03030_ _03026_ vssd1 vssd1 vccd1 vccd1
+ _00825_ sky130_fd_sc_hd__o211a_1
XFILLER_93_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20345__355 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__inv_2
X_16772_ _09408_ _09413_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__xnor2_1
X_13984_ _06710_ _06713_ _06718_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__nand3_1
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18511_ _02078_ _02081_ _02207_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__nand3_1
X_15723_ _08350_ _08351_ _08366_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__nand3_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _05665_ _05666_ _05670_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a22o_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19491_ _02967_ _02970_ _04033_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _10271_ _02028_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__nand2_1
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _08256_ _08258_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _04031_ _05372_ _05602_ _04001_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a211o_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _07340_ _07341_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__and2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _04594_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_6
X_18373_ _01498_ _09027_ _09162_ _10239_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__o22a_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _08002_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__clkbuf_4
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ rbzero.wall_tracer.mapY\[7\] _05397_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__and2_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _09890_ _09891_ _09892_ vssd1 vssd1 vccd1 vccd1 _09893_ sky130_fd_sc_hd__or3_1
X_14536_ _07250_ _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__or2_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11748_ _04523_ _04524_ _04525_ _04139_ _04208_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__o221a_1
XFILLER_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09831_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14467_ _06689_ _06761_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__or2_1
XFILLER_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11679_ _04434_ _04447_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__and2_2
X_16206_ _08850_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__inv_2
X_13418_ _06015_ _06031_ _05982_ _05974_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__o22a_1
XFILLER_139_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17186_ _09772_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__clkbuf_1
X_14398_ _07114_ _07127_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or2_1
X_16137_ _08748_ _08745_ _08746_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__and3_1
X_13349_ _06081_ _06085_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20090__125 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__inv_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16068_ _08698_ _08711_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__and2b_1
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__nor2_1
XFILLER_97_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19827_ rbzero.debug_overlay.playerX\[-8\] vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__inv_2
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19758_ _03107_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18709_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _02401_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__and4_1
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19689_ _03071_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03289_ _03289_ vssd1 vssd1 vccd1 vccd1 clknet_0__03289_ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21651_ clknet_leaf_43_i_clk _01420_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20602_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__or2_1
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21582_ net503 _01351_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20533_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03425_
+ sky130_fd_sc_hd__nand2_1
XFILLER_123_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20464_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03367_
+ sky130_fd_sc_hd__or2_1
XFILLER_192_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21016_ clknet_leaf_68_i_clk _00785_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_leak
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10981_ _03838_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ _05421_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__xnor2_2
XFILLER_128_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ rbzero.debug_overlay.playerY\[4\] _05401_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05402_ sky130_fd_sc_hd__mux2_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11602_ rbzero.tex_r1\[59\] rbzero.tex_r1\[58\] _04338_ vssd1 vssd1 vccd1 vccd1 _04381_
+ sky130_fd_sc_hd__mux2_1
X_12582_ _05289_ _05295_ _05303_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__and3_1
X_15370_ _05351_ _05475_ _07893_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__mux2_1
XFILLER_196_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ _07055_ _07057_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11533_ _04206_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nand2_1
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17040_ _09659_ _09679_ vssd1 vssd1 vccd1 vccd1 _09680_ sky130_fd_sc_hd__xnor2_2
X_14252_ _06951_ _06962_ _06984_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__or4_1
XFILLER_144_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11464_ _04121_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__buf_4
XFILLER_137_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13203_ _05923_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__xnor2_4
X_10415_ _03539_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
X_14183_ _06709_ _06918_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__or2_1
X_11395_ _04154_ _04157_ _04158_ gpout0.hpos\[9\] _04174_ vssd1 vssd1 vccd1 vccd1
+ _04175_ sky130_fd_sc_hd__a221o_1
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ rbzero.tex_r1\[45\] rbzero.tex_r1\[46\] _03494_ vssd1 vssd1 vccd1 vccd1 _03503_
+ sky130_fd_sc_hd__mux2_1
X_13134_ _05700_ _05703_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nor2_2
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18991_ rbzero.pov.spi_buffer\[28\] rbzero.pov.ready_buffer\[28\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_152_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _05710_ _05715_ _05718_ _05713_ _05777_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_
+ sky130_fd_sc_hd__mux4_1
X_17942_ _10133_ _10135_ _10126_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a21boi_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12016_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _04392_ vssd1 vssd1 vccd1 vccd1 _04791_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17873_ _09391_ _09351_ _09483_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__or3_1
X_16824_ _09463_ _09464_ vssd1 vssd1 vccd1 vccd1 _09466_ sky130_fd_sc_hd__and2_1
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19543_ rbzero.wall_tracer.rayAddendY\[11\] _03017_ vssd1 vssd1 vccd1 vccd1 _03018_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16755_ _09395_ _09396_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__xnor2_1
X_13967_ _06031_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _08323_ _08317_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__or2b_1
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03043_ clknet_0__03043_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03043_
+ sky130_fd_sc_hd__clkbuf_16
X_12918_ _05652_ _05654_ _05567_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21oi_1
X_19474_ _07678_ _02953_ _02954_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and3_1
XFILLER_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20404__5 clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
X_16686_ _09208_ _09327_ vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__or2_1
XFILLER_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ _06586_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18425_ _02006_ _02008_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__o21a_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ _07977_ vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__clkbuf_4
X_12849_ _05570_ _05360_ _05585_ _05561_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__o211a_1
XFILLER_62_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18356_ _02035_ _02054_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__xnor2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _08002_ _08212_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__nor2_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17307_ _09812_ _09876_ _09877_ vssd1 vssd1 vccd1 vccd1 _09878_ sky130_fd_sc_hd__o21ai_1
X_14519_ _07231_ _07255_ _05752_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__o21a_1
XFILLER_175_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18287_ _01985_ _01986_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__and2_1
XFILLER_148_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15499_ _08138_ _08142_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__nor2_1
XFILLER_175_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17238_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09813_ _09814_ vssd1 vssd1 vccd1 vccd1 _09816_ sky130_fd_sc_hd__a22oi_1
XFILLER_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17169_ rbzero.traced_texa\[-2\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a22o_1
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21634_ clknet_leaf_37_i_clk _01403_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21565_ net486 _01334_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20374__381 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__inv_2
X_20516_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03411_
+ sky130_fd_sc_hd__or2_1
XFILLER_154_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21496_ net417 _01265_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20447_ _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__and2b_1
XFILLER_181_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11180_ _03955_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__and2_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14870_ _05737_ _05736_ _07584_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__or3_2
XFILLER_208_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13821_ _06425_ _06555_ _06557_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a21bo_1
XFILLER_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16540_ _09022_ _09024_ vssd1 vssd1 vccd1 vccd1 _09184_ sky130_fd_sc_hd__nor2_1
X_13752_ _06468_ _06482_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a21bo_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ rbzero.tex_b1\[10\] rbzero.tex_b1\[11\] _03828_ vssd1 vssd1 vccd1 vccd1 _03830_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12703_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__or2_1
X_16471_ _08282_ _09114_ _08964_ vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__or3_1
X_13683_ _06418_ _06393_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__and2b_1
XFILLER_189_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10895_ _03793_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18210_ _01793_ _01795_ _01794_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a21boi_1
XFILLER_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15422_ rbzero.debug_overlay.playerX\[-3\] vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__inv_2
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19190_ rbzero.spi_registers.got_new_sky _02707_ vssd1 vssd1 vccd1 vccd1 _02740_
+ sky130_fd_sc_hd__nand2_2
X_12634_ _05386_ _03933_ _05284_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__mux2_1
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ _08257_ _01476_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__nor2_1
X_15353_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] rbzero.debug_overlay.playerX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _05308_ _05312_ _05314_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__o211a_1
XFILLER_184_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14304_ _06995_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__xor2_4
XFILLER_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11516_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _04291_ vssd1 vssd1 vccd1 vccd1 _04296_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18072_ _01770_ _01771_ _01772_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a21o_1
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15284_ _07925_ _07927_ _07928_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__a21oi_2
XFILLER_89_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12496_ rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__inv_2
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ _08202_ _08203_ _08129_ vssd1 vssd1 vccd1 vccd1 _09663_ sky130_fd_sc_hd__a21o_1
X_14235_ _06938_ _06971_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__and2_1
X_11447_ rbzero.tex_r0\[56\] _04214_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__a21o_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14166_ _06853_ _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__or2_1
X_11378_ rbzero.row_render.size\[9\] _04155_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nor2_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10329_ _03482_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__clkbuf_4
X_13117_ _05812_ _05821_ _05799_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__mux2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _06825_ _06832_ _06833_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__a21o_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _02617_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _05701_ _05682_ _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__or3_1
X_17925_ _09674_ _09417_ _01504_ _01627_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__o31a_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17856_ _01553_ _01559_ rbzero.wall_tracer.trackDistX\[3\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00592_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16807_ _09239_ _09317_ _09315_ vssd1 vssd1 vccd1 vccd1 _09449_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17787_ _01457_ _01490_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14999_ rbzero.wall_tracer.stepDistX\[6\] _07571_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07670_ sky130_fd_sc_hd__mux2_1
XFILLER_81_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19526_ _03000_ _03001_ _03002_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a21oi_1
X_16738_ _09263_ _09349_ _09378_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__nand3_1
X_19457_ rbzero.debug_overlay.vplaneY\[0\] rbzero.debug_overlay.vplaneY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__and2_1
XFILLER_62_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16669_ _09309_ _09310_ _09266_ vssd1 vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__a21o_1
X_18408_ _01965_ _01929_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__or2b_1
XFILLER_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19388_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nand2_1
XFILLER_194_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18339_ _02036_ _02037_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__nand2_1
XFILLER_72_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21350_ net271 _01119_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21281_ clknet_leaf_34_i_clk _01050_ vssd1 vssd1 vccd1 vccd1 rbzero.hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20094_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__buf_1
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19631__83 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__inv_2
XFILLER_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20996_ clknet_leaf_52_i_clk _00765_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_69_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_198_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ rbzero.tex_g1\[17\] rbzero.tex_g1\[18\] _03680_ vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21617_ clknet_leaf_33_i_clk _01386_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12350_ _04813_ _04811_ _04006_ _03475_ _05083_ _05082_ vssd1 vssd1 vccd1 vccd1 _05118_
+ sky130_fd_sc_hd__mux4_1
X_21548_ net469 _01317_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11301_ _04077_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nor2_1
X_12281_ _04021_ _05047_ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and3_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21479_ net400 _01248_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14020_ _06755_ _06756_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__nor2_1
XFILLER_84_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _04016_ _03997_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__or2_2
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11163_ _03946_ _03949_ _03950_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__or4_1
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15971_ _08584_ _08614_ _08615_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__a21oi_2
X_11094_ _03897_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17710_ _10122_ _10146_ _10274_ vssd1 vssd1 vccd1 vccd1 _10275_ sky130_fd_sc_hd__a21o_1
X_14922_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.trackDistX\[-1\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__mux2_1
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18690_ _02383_ _02385_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__xnor2_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _09526_ _09029_ _09165_ _09245_ vssd1 vssd1 vccd1 vccd1 _10206_ sky130_fd_sc_hd__o22a_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14853_ rbzero.wall_tracer.stepDistY\[6\] _07571_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07572_ sky130_fd_sc_hd__mux2_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _06534_ _06538_ _06539_ _06540_ _06518_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__a311o_1
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17572_ rbzero.wall_tracer.stepDistX\[10\] vssd1 vssd1 vccd1 vccd1 _10138_ sky130_fd_sc_hd__inv_2
X_14784_ _07498_ _07489_ _05952_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__mux2_1
XFILLER_205_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11996_ _04232_ _04758_ _04762_ _04770_ _04244_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__o311a_1
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19311_ _02811_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16523_ _09033_ _09035_ _09032_ vssd1 vssd1 vccd1 vccd1 _09167_ sky130_fd_sc_hd__a21bo_1
X_13735_ _06382_ _06153_ _06469_ _06470_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__a22o_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10947_ rbzero.tex_b1\[18\] rbzero.tex_b1\[19\] _03817_ vssd1 vssd1 vccd1 vccd1 _03821_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19242_ _02561_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__or2_1
X_16454_ _09095_ _09097_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__and2_1
X_13666_ _06356_ _06401_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ rbzero.tex_b1\[51\] rbzero.tex_b1\[52\] _03784_ vssd1 vssd1 vccd1 vccd1 _03785_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15405_ rbzero.wall_tracer.side rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1
+ vccd1 _08050_ sky130_fd_sc_hd__nand2_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _05324_ _05325_ _05326_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a21bo_1
X_19173_ _05190_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__buf_4
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _09029_ _08162_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__nor2_2
X_13597_ _06279_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__and2_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18124_ _09391_ _09703_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__and2_1
X_15336_ _07980_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__clkbuf_4
X_12548_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__nor2_1
XFILLER_157_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18055_ _08895_ _01524_ _10266_ _08767_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__o22ai_1
X_15267_ _05206_ _07902_ _07910_ _07911_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__a22o_2
XANTENNA_2 _04021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _05233_ _05216_ _05213_ _05230_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or4_1
XFILLER_172_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _09640_ _09645_ vssd1 vssd1 vccd1 vccd1 _09646_ sky130_fd_sc_hd__xnor2_1
X_14218_ _06892_ _06954_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15198_ _07849_ _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__nand2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14149_ _06860_ _06874_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20210__233 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__inv_2
XFILLER_140_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957_ _02608_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17908_ _01609_ _01610_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__and2_1
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18888_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__nor2b_2
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17839_ _01454_ _01542_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20850_ clknet_leaf_93_i_clk _00619_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19509_ _03913_ _02986_ _02987_ _07855_ rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__a32o_1
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20781_ clknet_leaf_21_i_clk _00550_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21402_ net323 _01171_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21333_ net254 _01102_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21264_ clknet_leaf_62_i_clk _01033_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21195_ clknet_leaf_64_i_clk _00964_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20185__210 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__inv_2
XFILLER_170_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11850_ _04244_ _04618_ _04626_ _04116_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a31o_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _03744_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11781_ _04557_ _04558_ _04218_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20979_ clknet_leaf_52_i_clk _00748_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ _06214_ _06217_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__and2b_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10732_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _03706_ vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ _06172_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ rbzero.tex_g1\[25\] rbzero.tex_g1\[26\] _03669_ vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12402_ _04813_ _04811_ _05143_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__mux2_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16170_ _08813_ _08814_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__or2_1
X_13382_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__nand2_1
XFILLER_166_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10594_ _03482_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15121_ _07754_ _07763_ _07764_ _07749_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__o2bb2ai_1
X_12333_ _05100_ net28 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__nand2_1
XFILLER_166_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15052_ _07712_ _07714_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__xnor2_1
X_12264_ net22 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__inv_2
XFILLER_181_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__clkbuf_4
X_11215_ rbzero.wall_tracer.state\[11\] vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__inv_2
X_12195_ _04962_ _04963_ _04964_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__and3_1
X_19860_ rbzero.debug_overlay.playerX\[1\] _03167_ vssd1 vssd1 vccd1 vccd1 _03172_
+ sky130_fd_sc_hd__and2_1
XFILLER_134_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 o_rgb[14] sky130_fd_sc_hd__buf_2
XFILLER_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18811_ _05254_ _08186_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__nor2_1
X_11146_ rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__inv_2
X_19791_ _03124_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11077_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _03887_ vssd1 vssd1 vccd1 vccd1 _03889_
+ sky130_fd_sc_hd__mux2_1
X_15954_ _08590_ _08597_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__nor2_1
X_18742_ _02428_ _02429_ _02430_ _05531_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a31o_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03291_ clknet_0__03291_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03291_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14905_ _07591_ _07610_ _07611_ _04039_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__o211a_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18673_ _01737_ _01524_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__or2_1
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _08526_ _08528_ _08529_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__a21oi_2
XFILLER_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17624_ _10064_ _10067_ _10188_ vssd1 vssd1 vccd1 vccd1 _10189_ sky130_fd_sc_hd__a21o_1
XFILLER_97_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19610__64 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _10119_ _10120_ vssd1 vssd1 vccd1 vccd1 _10121_ sky130_fd_sc_hd__or2b_1
XFILLER_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _05814_ _07496_ _07500_ _07486_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a211oi_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11979_ _04242_ _04745_ _04753_ _04207_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__o211a_1
XFILLER_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _08991_ _08993_ vssd1 vssd1 vccd1 vccd1 _09150_ sky130_fd_sc_hd__or2b_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13718_ _06439_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__xor2_1
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17486_ _09971_ _09957_ vssd1 vssd1 vccd1 vccd1 _10052_ sky130_fd_sc_hd__or2b_1
XFILLER_189_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14698_ _07106_ _07419_ _07420_ _07423_ _05892_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__a311o_1
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19225_ rbzero.spi_registers.got_new_vshift _02711_ vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__nand2_1
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16437_ _09081_ vssd1 vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__clkbuf_4
X_13649_ _06339_ _06383_ _06384_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19156_ rbzero.otherx\[4\] _02710_ _02718_ _02714_ vssd1 vssd1 vccd1 vccd1 _00733_
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16368_ _09011_ _09012_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18107_ _01701_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__inv_2
XFILLER_121_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _04013_ _07962_ _07963_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__a21oi_4
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19087_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ _02567_ _02558_ _02557_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__o311a_1
X_16299_ _08764_ _08807_ _08811_ _08940_ _08943_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__a32oi_4
X_18038_ _01739_ _10238_ _09552_ _01737_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__o22ai_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20000_ rbzero.pov.ready_buffer\[4\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-5\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__a221o_1
XFILLER_87_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19989_ rbzero.pov.ready_buffer\[15\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-5\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__a221o_1
XFILLER_80_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20902_ clknet_leaf_81_i_clk _00671_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ clknet_leaf_27_i_clk _00602_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20764_ clknet_leaf_32_i_clk _00533_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20695_ clknet_leaf_6_i_clk _00479_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20217__239 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__inv_2
XFILLER_191_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21316_ net237 _01085_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21247_ clknet_leaf_80_i_clk _01016_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_172_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11000_ _03848_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21178_ clknet_leaf_74_i_clk _00947_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__inv_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ rbzero.tex_b0\[3\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and3_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15670_ _07959_ _07941_ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__nor2_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _05610_ _05612_ _05615_ _05601_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a2111o_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _07316_ _07317_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__xnor2_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _04242_ _04601_ _04609_ _04207_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__o211a_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _09486_ _09495_ vssd1 vssd1 vccd1 vccd1 _09907_ sky130_fd_sc_hd__and2b_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _07058_ _06999_ _07000_ _07057_ _07055_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__o32ai_2
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _04540_ _04541_ _04126_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _06159_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__clkbuf_4
XFILLER_144_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17271_ _09845_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ rbzero.tex_g1\[0\] rbzero.tex_g1\[1\] _03691_ vssd1 vssd1 vccd1 vccd1 _03699_
+ sky130_fd_sc_hd__mux2_1
X_14483_ _07168_ _07219_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__nand2_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ rbzero.debug_overlay.vplaneY\[-7\] _04455_ _04465_ rbzero.debug_overlay.vplaneY\[-1\]
+ _04040_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a221o_1
XFILLER_186_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19010_ net511 rbzero.pov.ready_buffer\[37\] _02627_ vssd1 vssd1 vccd1 vccd1 _02636_
+ sky130_fd_sc_hd__mux2_1
X_16222_ _08865_ _08866_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__and2_1
X_13434_ _06004_ _06005_ _06019_ _06020_ _06001_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a32o_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10646_ rbzero.tex_g1\[33\] rbzero.tex_g1\[34\] _03658_ vssd1 vssd1 vccd1 vccd1 _03663_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16153_ _08779_ _08797_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__nand2_1
X_13365_ _06100_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or2_1
X_10577_ _03626_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _04462_ rbzero.debug_overlay.vplaneX\[-7\] vssd1 vssd1 vccd1 vccd1 _07763_
+ sky130_fd_sc_hd__xnor2_1
X_20157__186 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__inv_2
X_12316_ _05082_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__nor2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16084_ _07912_ _08125_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__or2_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13296_ _05939_ _05975_ _05962_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__or3b_1
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15035_ _07680_ _07693_ _07681_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__o21ai_1
X_19912_ rbzero.pov.ready_buffer\[51\] _02823_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__nand2_1
X_12247_ _04996_ _05013_ _05016_ net16 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o22a_1
XFILLER_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19843_ _03139_ _03158_ _03159_ _03157_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__o211a_1
X_12178_ _04883_ _04884_ gpout0.vpos\[6\] _04887_ _04910_ net10 vssd1 vssd1 vccd1
+ vccd1 _04949_ sky130_fd_sc_hd__mux4_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11129_ rbzero.wall_tracer.visualWallDist\[10\] rbzero.wall_tracer.visualWallDist\[9\]
+ _03916_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or4_1
X_19774_ rbzero.pov.spi_buffer\[60\] rbzero.pov.spi_buffer\[61\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_1
X_16986_ _09624_ _09625_ vssd1 vssd1 vccd1 vccd1 _09626_ sky130_fd_sc_hd__and2_1
XFILLER_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18725_ _02414_ _02415_ _02416_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__and3_1
XFILLER_77_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _08578_ _08580_ _08581_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__o21ai_2
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15868_ _08456_ _08457_ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__xnor2_1
X_18656_ _02247_ _02236_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__and2b_1
XFILLER_37_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20322__334 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__inv_2
XFILLER_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17607_ _10172_ vssd1 vssd1 vccd1 vccd1 _10173_ sky130_fd_sc_hd__inv_2
XFILLER_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14819_ rbzero.wall_tracer.stepDistY\[-3\] _07545_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07547_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18587_ _02282_ _02283_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__nor2_1
X_15799_ _08379_ _08443_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__xor2_4
XFILLER_184_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17538_ _09670_ _09964_ vssd1 vssd1 vccd1 vccd1 _10104_ sky130_fd_sc_hd__nand2_1
XFILLER_177_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17469_ _09817_ vssd1 vssd1 vccd1 vccd1 _10036_ sky130_fd_sc_hd__buf_2
XFILLER_177_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19208_ rbzero.spi_registers.new_floor\[0\] rbzero.color_floor\[0\] _02751_ vssd1
+ vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20480_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__inv_2
XFILLER_158_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19139_ _04037_ _02705_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21101_ net191 _00870_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21032_ clknet_leaf_51_i_clk _00801_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20297__311 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__inv_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ clknet_leaf_8_i_clk _00585_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20747_ clknet_leaf_36_i_clk _00516_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _03580_ vssd1 vssd1 vccd1 vccd1 _03586_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ _04219_ _04259_ _04254_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o21a_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20678_ clknet_leaf_3_i_clk _00462_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[7\]
+ sky130_fd_sc_hd__dfxtp_4
Xclkbuf_1_0__f__03294_ clknet_0__03294_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03294_
+ sky130_fd_sc_hd__clkbuf_16
X_10431_ _03547_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ _05883_ _05886_ _05798_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__o21a_1
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10362_ _03511_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12101_ _04317_ _04853_ _04838_ _03473_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _05690_ _05796_ _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__o21a_1
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _04805_ _04806_ _04206_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__mux2_1
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16840_ rbzero.wall_tracer.visualWallDist\[10\] _04015_ vssd1 vssd1 vccd1 vccd1 _09481_
+ sky130_fd_sc_hd__nand2_1
XFILLER_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16771_ _09411_ _09412_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__xor2_1
X_13983_ _06674_ _06679_ _06673_ _06683_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a22oi_2
XFILLER_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15722_ _08350_ _08351_ _08366_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__a21o_1
X_18510_ _02078_ _02081_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a21o_1
X_12934_ _05563_ _05653_ _05669_ _05650_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a211o_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _02968_ _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__xor2_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _02028_ _01645_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__and2b_1
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15653_ _08262_ _08278_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__xnor2_2
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ rbzero.wall_tracer.visualWallDist\[5\] _04031_ vssd1 vssd1 vccd1 vccd1 _05602_
+ sky130_fd_sc_hd__nor2_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _07206_ _07339_ _07338_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__or3_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20163__190 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__inv_2
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11816_ _04591_ _04593_ _04324_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21ba_1
X_18372_ _01498_ _09162_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nor2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _08216_ _08228_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__xnor2_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _05533_ _05537_ _05538_ _05284_ rbzero.wall_tracer.mapY\[6\] vssd1 vssd1
+ vccd1 vccd1 _00413_ sky130_fd_sc_hd__a32o_1
XFILLER_199_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _09880_ _09882_ _09881_ vssd1 vssd1 vccd1 vccd1 _09892_ sky130_fd_sc_hd__a21boi_1
XFILLER_183_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14535_ _07252_ _07267_ _07271_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__o21a_1
XFILLER_159_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11747_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _04271_ vssd1 vssd1 vccd1 vccd1 _04525_
+ sky130_fd_sc_hd__mux2_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17254_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09830_ sky130_fd_sc_hd__or2_1
XFILLER_202_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ _07132_ _07201_ _07202_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__o21ai_1
XFILLER_159_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ rbzero.debug_overlay.vplaneX\[-5\] _04454_ _04455_ rbzero.debug_overlay.vplaneX\[-7\]
+ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__a221o_1
XFILLER_186_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _08845_ _08847_ _08849_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__a21o_1
X_13417_ _05752_ _06153_ _05976_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__and3_1
X_10629_ rbzero.tex_g1\[41\] rbzero.tex_g1\[42\] _03647_ vssd1 vssd1 vccd1 vccd1 _03654_
+ sky130_fd_sc_hd__mux2_1
X_17185_ rbzero.wall_tracer.wall\[0\] rbzero.row_render.wall\[0\] _07830_ vssd1 vssd1
+ vccd1 vccd1 _09772_ sky130_fd_sc_hd__mux2_1
X_14397_ _07114_ _07127_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__nand2_1
XFILLER_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16136_ _08743_ _08750_ vssd1 vssd1 vccd1 vccd1 _08781_ sky130_fd_sc_hd__or2_1
X_13348_ _06041_ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__nor2_1
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16067_ _08698_ _08711_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__xnor2_1
X_13279_ _06011_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15018_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__or2_1
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19826_ rbzero.pov.ready_buffer\[60\] _07985_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19757_ rbzero.pov.spi_buffer\[52\] rbzero.pov.spi_buffer\[53\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_49_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16969_ _09485_ _09486_ _09497_ _09608_ vssd1 vssd1 vccd1 vccd1 _09609_ sky130_fd_sc_hd__a31o_1
XFILLER_204_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18708_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__nand2_1
X_19688_ rbzero.pov.spi_buffer\[19\] rbzero.pov.spi_buffer\[20\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _02333_ _02334_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21650_ clknet_leaf_18_i_clk _01419_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20601_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__nand2_1
XFILLER_71_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21581_ net502 _01350_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20532_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03424_
+ sky130_fd_sc_hd__nor2_1
XFILLER_119_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20463_ _03272_ _03365_ _03366_ _03327_ rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1
+ _01392_ sky130_fd_sc_hd__a32o_1
XFILLER_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21015_ clknet_leaf_67_i_clk _00784_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10980_ rbzero.tex_b1\[2\] rbzero.tex_b1\[3\] _03828_ vssd1 vssd1 vccd1 vccd1 _03838_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12650_ _05398_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ rbzero.tex_r1\[56\] _04273_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a21o_1
XFILLER_208_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12581_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or2_1
XFILLER_157_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14320_ _07013_ _07014_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__o21a_1
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ rbzero.color_sky\[0\] rbzero.color_floor\[0\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04312_ sky130_fd_sc_hd__mux2_1
XFILLER_184_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _06986_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11463_ _04230_ _04236_ _04240_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__a211o_1
XFILLER_172_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__buf_4
X_10414_ rbzero.tex_r1\[13\] rbzero.tex_r1\[14\] _03538_ vssd1 vssd1 vccd1 vccd1 _03539_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14182_ _06709_ _06918_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__nand2_1
XFILLER_183_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ gpout0.hpos\[7\] _04159_ _04157_ gpout0.hpos\[8\] _04173_ vssd1 vssd1 vccd1
+ vccd1 _04174_ sky130_fd_sc_hd__o221a_1
XFILLER_174_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20351__360 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__inv_2
XFILLER_178_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _05820_ _05866_ _05869_ _05813_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__o211a_1
XFILLER_125_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10345_ _03502_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
X_18990_ _02625_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13064_ _05796_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__clkbuf_4
X_17941_ _01641_ _01642_ _01634_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a21o_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12015_ _04788_ _04789_ _04304_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__mux2_1
XFILLER_39_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17872_ _01494_ _01512_ _01574_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20269__287 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__inv_2
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16823_ _09463_ _09464_ vssd1 vssd1 vccd1 vccd1 _09465_ sky130_fd_sc_hd__nor2_1
XFILLER_207_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19542_ _07677_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__nor2_1
X_13966_ _06685_ _06695_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__a21oi_2
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16754_ _08111_ _08264_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__and2b_1
XFILLER_207_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03042_ clknet_0__03042_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03042_
+ sky130_fd_sc_hd__clkbuf_16
X_15705_ _08320_ _08322_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__nand2_1
X_12917_ _05563_ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__nand2_1
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16685_ _09208_ _09327_ vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__nand2_1
X_19473_ _02951_ _02952_ _02950_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a21o_1
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13897_ _06632_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__and2_1
XFILLER_206_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18424_ _02009_ _01917_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or2b_1
X_15636_ _08249_ _08280_ vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__xor2_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ rbzero.wall_tracer.visualWallDist\[-6\] rbzero.wall_tracer.rcp_sel\[2\] vssd1
+ vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or2_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18355_ _02038_ _02053_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__xnor2_1
X_15567_ _07894_ _05331_ _08211_ _07970_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__o211a_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ rbzero.map_rom.i_col\[4\] _05523_ _05414_ vssd1 vssd1 vccd1 vccd1 _05524_
+ sky130_fd_sc_hd__mux2_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _07230_ _07229_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__and2b_1
X_17306_ _09807_ _09331_ vssd1 vssd1 vccd1 vccd1 _09877_ sky130_fd_sc_hd__or2_1
X_15498_ _08138_ _08142_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__xor2_1
X_18286_ _01860_ _01620_ _01984_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__o21ai_1
XFILLER_175_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ _07114_ _07185_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__nor2_1
XFILLER_147_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17237_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09813_ _09814_ vssd1 vssd1 vccd1 vccd1 _09815_ sky130_fd_sc_hd__and4_1
XFILLER_175_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17168_ _07679_ vssd1 vssd1 vccd1 vccd1 _09769_ sky130_fd_sc_hd__buf_2
XFILLER_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16119_ _08719_ _08763_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__xor2_2
XFILLER_66_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17099_ _09737_ _09738_ vssd1 vssd1 vccd1 vccd1 _09739_ sky130_fd_sc_hd__xnor2_4
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19809_ _03133_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03309_ clknet_0__03309_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03309_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21633_ clknet_leaf_37_i_clk _01402_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21564_ net485 _01333_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20515_ rbzero.texV\[4\] _03327_ _03332_ _03410_ vssd1 vssd1 vccd1 vccd1 _01400_
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21495_ net416 _01264_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20446_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _03352_
+ sky130_fd_sc_hd__nand2_1
XFILLER_107_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _06279_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__xnor2_2
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _06486_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__nand2_1
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10963_ _03829_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12702_ _05446_ _05447_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__o21a_1
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16470_ _07959_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__clkbuf_4
X_13682_ _06393_ _06418_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__xnor2_1
X_10894_ rbzero.tex_b1\[43\] rbzero.tex_b1\[44\] _03784_ vssd1 vssd1 vccd1 vccd1 _03793_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ _08027_ _08065_ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__nand2_1
X_12633_ rbzero.debug_overlay.playerY\[2\] _05385_ _05204_ vssd1 vssd1 vccd1 vccd1
+ _05386_ sky130_fd_sc_hd__mux2_1
XFILLER_197_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ _07977_ _07981_ _07989_ _07996_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__o22ai_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18140_ _01498_ _01475_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__nor2_1
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__inv_2
X_14303_ _07035_ _07038_ _07039_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__nor3b_2
X_11515_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _04291_ vssd1 vssd1 vccd1 vccd1 _04295_
+ sky130_fd_sc_hd__mux2_1
X_18071_ _01770_ _01771_ _01772_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nand3_1
XFILLER_129_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15283_ _07904_ rbzero.wall_tracer.stepDistY\[-4\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _07928_ sky130_fd_sc_hd__a21o_1
X_12495_ rbzero.wall_tracer.trackDistY\[-5\] _05236_ rbzero.wall_tracer.trackDistY\[-6\]
+ _05237_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__o221a_1
XFILLER_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17022_ _08204_ _09103_ _08493_ _08383_ vssd1 vssd1 vccd1 vccd1 _09662_ sky130_fd_sc_hd__o22ai_1
X_14234_ _06805_ _06678_ _06937_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__o21bai_1
X_20275__291 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__inv_2
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__buf_4
XFILLER_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14165_ _06680_ _06690_ _06672_ _06675_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__o22a_1
X_11377_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__and2_1
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ _05794_ _05828_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__or2_2
X_10328_ _03493_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14096_ _06826_ _06831_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__nor2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ rbzero.pov.spi_buffer\[19\] rbzero.pov.ready_buffer\[19\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XFILLER_124_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _05719_ _05721_ _05705_ _05783_ _05710_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o32a_1
XFILLER_117_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17924_ _10244_ _01503_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _09889_ _01558_ _09781_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _09382_ _09447_ vssd1 vssd1 vccd1 vccd1 _09448_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17786_ _01471_ _01489_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__xor2_1
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14998_ _07669_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19525_ _02906_ rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 _03002_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16737_ _09263_ _09349_ _09378_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__a21o_1
X_13949_ _06665_ _06670_ _06684_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__nand3_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19456_ rbzero.debug_overlay.vplaneY\[0\] rbzero.debug_overlay.vplaneY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__nor2_1
X_16668_ _09266_ _09309_ _09310_ vssd1 vssd1 vccd1 vccd1 _09311_ sky130_fd_sc_hd__nand3_1
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18407_ _01964_ _01932_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__or2b_1
X_15619_ _08199_ _08201_ _08203_ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__a21bo_2
X_19387_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__nand2_1
XFILLER_188_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16599_ _09124_ _09116_ vssd1 vssd1 vccd1 vccd1 _09242_ sky130_fd_sc_hd__or2b_1
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18338_ _01971_ _01968_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__or2b_1
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18269_ _10110_ _01524_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__nor2_1
XFILLER_129_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21280_ clknet_leaf_31_i_clk _01049_ vssd1 vssd1 vccd1 vccd1 rbzero.vga_sync.vsync
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20995_ clknet_leaf_58_i_clk _00764_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21616_ clknet_3_5_0_i_clk _01385_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21547_ net468 _01316_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ rbzero.texV\[3\] _04078_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a21boi_1
XFILLER_181_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12280_ net21 net20 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and2_2
XFILLER_166_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21478_ net399 _01247_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11231_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__clkinv_4
XFILLER_181_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20429_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03338_
+ sky130_fd_sc_hd__or2_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03045_ clknet_0__03045_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03045_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11162_ rbzero.wall_tracer.mapX\[11\] rbzero.wall_tracer.mapX\[10\] rbzero.wall_tracer.mapY\[7\]
+ rbzero.wall_tracer.mapY\[6\] vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or4_1
XFILLER_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15970_ _08585_ _08613_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__nor2_1
X_11093_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _03887_ vssd1 vssd1 vccd1 vccd1 _03897_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14921_ _07621_ _07622_ _07623_ _07620_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__o211a_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _08705_ _09029_ _09165_ vssd1 vssd1 vccd1 vccd1 _10205_ sky130_fd_sc_hd__or3_1
XFILLER_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14852_ _07394_ _07433_ _07418_ _07468_ _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__a311o_4
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _06503_ _06516_ _06517_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__a21oi_1
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14783_ _00004_ _07514_ _07515_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17571_ _09117_ _09977_ vssd1 vssd1 vccd1 vccd1 _10137_ sky130_fd_sc_hd__nor2_1
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11995_ _04306_ _04765_ _04769_ _04241_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a211o_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ rbzero.spi_registers.new_other\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _02800_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__mux2_1
XFILLER_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13734_ _06382_ _06153_ _06469_ _06470_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__nand4_1
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16522_ _09029_ _08160_ _09165_ _08162_ vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__o22a_1
XFILLER_95_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10946_ _03820_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19241_ rbzero.spi_registers.spi_done _03480_ _02560_ vssd1 vssd1 vccd1 vccd1 _02772_
+ sky130_fd_sc_hd__nand3_1
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _06041_ _06016_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__or2_1
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16453_ _09096_ _08356_ _09094_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__o21ai_1
XFILLER_189_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10877_ _03646_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _05342_ _05345_ _05365_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4b_1
X_15404_ rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__inv_2
XFILLER_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16384_ _09028_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__buf_2
X_19172_ rbzero.spi_registers.got_new_vinf _02711_ rbzero.row_render.vinf vssd1 vssd1
+ vccd1 vccd1 _02729_ sky130_fd_sc_hd__a21o_1
X_13596_ _06331_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__and2b_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18123_ _01822_ _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__or2_1
X_15335_ rbzero.debug_overlay.playerX\[-9\] _05206_ _07979_ vssd1 vssd1 vccd1 vccd1
+ _07980_ sky130_fd_sc_hd__a21oi_4
X_12547_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__and2_1
XFILLER_185_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _10131_ _10132_ _01525_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a21o_4
X_15266_ rbzero.wall_tracer.visualWallDist\[-6\] _04013_ _05195_ vssd1 vssd1 vccd1
+ vccd1 _07911_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12478_ _05219_ _05221_ _05223_ _05225_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__or4_1
XANTENNA_3 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14217_ _06900_ _06899_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__and2b_1
XFILLER_126_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17005_ _09641_ _09644_ vssd1 vssd1 vccd1 vccd1 _09645_ sky130_fd_sc_hd__xnor2_1
X_11429_ _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__buf_4
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ _07730_ _07833_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__nand2_1
XFILLER_67_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _06858_ _06876_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14079_ _06799_ _06814_ _06815_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__a21bo_1
X_18956_ rbzero.pov.spi_buffer\[11\] rbzero.pov.ready_buffer\[11\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
X_17907_ _01573_ _01608_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__or2_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18887_ net70 _03555_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__nor2_4
XFILLER_187_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17838_ _01539_ _01541_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__xor2_1
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17769_ _10240_ _10242_ _10237_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a21bo_1
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19508_ _02984_ _02985_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__or2_1
XFILLER_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20780_ clknet_leaf_22_i_clk _00549_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19439_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[2\] _02896_
+ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__o21bai_1
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03039_ _03039_ vssd1 vssd1 vccd1 vccd1 clknet_0__03039_ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20291__306 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__inv_2
X_21401_ net322 _01170_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21332_ net253 _01101_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21263_ clknet_leaf_61_i_clk _01032_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21194_ clknet_leaf_64_i_clk _00963_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _03740_ vssd1 vssd1 vccd1 vccd1 _03744_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11780_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _04262_ vssd1 vssd1 vccd1 vccd1 _04558_
+ sky130_fd_sc_hd__mux2_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20978_ clknet_leaf_49_i_clk _00747_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ _03707_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13450_ _06173_ _06186_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__xor2_1
XFILLER_139_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10662_ _03671_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ net34 _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and2_1
X_13381_ _06114_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__xnor2_2
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10593_ _03634_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ _07776_ _07777_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__or2_1
XFILLER_194_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12332_ net29 vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__inv_2
XFILLER_127_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _07713_ _07699_ _07698_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__a21oi_1
X_12263_ net21 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__inv_2
XFILLER_182_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ _06615_ _06738_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__or2_1
XFILLER_141_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11214_ rbzero.wall_tracer.state\[8\] vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__inv_2
XFILLER_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12194_ net18 net19 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__nor2_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18810_ _02491_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__clkbuf_1
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 o_rgb[15] sky130_fd_sc_hd__buf_2
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11145_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__inv_2
X_19790_ rbzero.pov.spi_buffer\[68\] rbzero.pov.spi_buffer\[69\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XFILLER_123_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18741_ _02428_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1__f__03290_ clknet_0__03290_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03290_
+ sky130_fd_sc_hd__clkbuf_16
X_11076_ _03888_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__clkbuf_1
X_15953_ _08590_ _08597_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__xor2_1
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14904_ rbzero.wall_tracer.visualWallDist\[-6\] _07595_ vssd1 vssd1 vccd1 vccd1 _07611_
+ sky130_fd_sc_hd__or2_1
X_18672_ _08047_ _09565_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__nor2_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _08517_ _08525_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__nor2_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17623_ _10053_ _10056_ _10054_ vssd1 vssd1 vccd1 vccd1 _10188_ sky130_fd_sc_hd__a21boi_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _07468_ _07557_ _07558_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__or3b_1
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _10118_ _10114_ vssd1 vssd1 vccd1 vccd1 _10120_ sky130_fd_sc_hd__or2b_1
XFILLER_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ _07473_ _07499_ _05814_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__a21oi_1
X_11978_ _04254_ _04748_ _04752_ _04371_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a211o_1
XFILLER_205_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16505_ _09125_ _09148_ vssd1 vssd1 vccd1 vccd1 _09149_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13717_ _06440_ _06452_ _06453_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21oi_1
X_10929_ _03811_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__clkbuf_1
X_14697_ _07394_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nand2_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17485_ _09958_ _09970_ vssd1 vssd1 vccd1 vccd1 _10051_ sky130_fd_sc_hd__nand2_1
XFILLER_205_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19224_ _02761_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__clkbuf_2
X_16436_ _05397_ _05503_ _07971_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__mux2_1
X_13648_ _06339_ _06383_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ rbzero.spi_registers.new_other\[10\] _02712_ vssd1 vssd1 vccd1 vccd1 _02718_
+ sky130_fd_sc_hd__or2_1
X_13579_ _06309_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__nand2_1
X_16367_ _07941_ _08097_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__or2_1
XFILLER_118_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18106_ _01705_ _01714_ _01712_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a21o_1
XFILLER_185_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15318_ _07903_ rbzero.wall_tracer.stepDistY\[-6\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _07963_ sky130_fd_sc_hd__a21o_1
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16298_ _08811_ _08942_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__xnor2_2
XFILLER_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19086_ _02675_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18037_ _08242_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__buf_2
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__buf_4
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_68_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20134__165 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__inv_2
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19988_ rbzero.pov.ready_buffer\[14\] _03252_ _03253_ rbzero.debug_overlay.vplaneX\[-6\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__o221a_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18939_ rbzero.pov.spi_buffer\[3\] rbzero.pov.ready_buffer\[3\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20901_ clknet_leaf_83_i_clk _00670_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ clknet_leaf_26_i_clk _00601_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20763_ clknet_leaf_32_i_clk _00532_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20694_ clknet_leaf_8_i_clk _00478_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21315_ net236 _01084_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21246_ clknet_leaf_80_i_clk _01015_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21177_ clknet_leaf_74_i_clk _00946_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12950_ _05685_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__xnor2_4
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11901_ _04675_ _04676_ _04139_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__mux2_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _05561_ _05461_ _05616_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o22a_2
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _05793_ _07356_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__and2_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11832_ _04306_ _04604_ _04608_ _04371_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a211o_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14551_ _07080_ _07082_ _07084_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__o21a_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _04129_ vssd1 vssd1 vccd1 vccd1 _04541_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _06015_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__clkbuf_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _03698_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__clkbuf_1
X_14482_ _07164_ _07167_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__nand2_1
X_17270_ rbzero.wall_tracer.trackDistX\[-8\] _09844_ _05414_ vssd1 vssd1 vccd1 vccd1
+ _09845_ sky130_fd_sc_hd__mux2_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _04471_ _04463_ _04459_ rbzero.debug_overlay.vplaneY\[0\] _04472_ vssd1 vssd1
+ vccd1 vccd1 _04473_ sky130_fd_sc_hd__a221o_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13433_ _06168_ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__or2_1
X_16221_ _08860_ _08864_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__nand2_1
X_10645_ _03662_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16152_ _08780_ _08781_ _08792_ _08794_ _08796_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__a32oi_2
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ _05946_ _05961_ _06007_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or3_1
XFILLER_194_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10576_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _03624_ vssd1 vssd1 vccd1 vccd1 _03626_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ net26 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15103_ _07758_ _07759_ _07760_ _07757_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__a22o_1
X_16083_ _07958_ _08572_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__or2_1
X_13295_ _05978_ _06031_ _05962_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__o21bai_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__and2_1
X_19911_ rbzero.debug_overlay.playerY\[-3\] _03198_ _03211_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00995_ sky130_fd_sc_hd__o211a_1
X_12246_ _04977_ _05014_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__o21ai_1
XFILLER_170_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19842_ _07949_ _03143_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__nand2_1
XFILLER_111_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ _04908_ _04943_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ rbzero.wall_tracer.visualWallDist\[4\] rbzero.wall_tracer.visualWallDist\[3\]
+ rbzero.wall_tracer.visualWallDist\[2\] rbzero.wall_tracer.visualWallDist\[1\] vssd1
+ vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or4_1
XFILLER_122_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19773_ _03115_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
X_16985_ _09620_ _09623_ vssd1 vssd1 vccd1 vccd1 _09625_ sky130_fd_sc_hd__or2_1
X_18724_ _02407_ _02408_ _02409_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__o21bai_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _03879_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__clkbuf_1
X_15936_ _08569_ _08577_ vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__or2_1
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18655_ _02139_ _02248_ _02140_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21a_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _08460_ _08461_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__xnor2_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ _05203_ _10171_ vssd1 vssd1 vccd1 vccd1 _10172_ sky130_fd_sc_hd__or2_1
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14818_ _05188_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__buf_4
X_18586_ _02269_ _02270_ _02281_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__and3_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _08259_ _08238_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__nor2_2
XFILLER_45_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17537_ _10101_ _10102_ vssd1 vssd1 vccd1 vccd1 _10103_ sky130_fd_sc_hd__xor2_1
X_14749_ _07468_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__or2_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17468_ _05532_ _10033_ _10034_ _09817_ vssd1 vssd1 vccd1 vccd1 _10035_ sky130_fd_sc_hd__o31a_1
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19207_ rbzero.spi_registers.got_new_floor _02707_ vssd1 vssd1 vccd1 vccd1 _02751_
+ sky130_fd_sc_hd__nand2_2
X_16419_ _09061_ _09062_ _09063_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__and3_1
XFILLER_121_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17399_ _08178_ _09103_ vssd1 vssd1 vccd1 vccd1 _09966_ sky130_fd_sc_hd__or2_1
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19138_ gpout0.vpos\[3\] _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__and2_1
XFILLER_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19069_ rbzero.pov.spi_buffer\[65\] rbzero.pov.ready_buffer\[65\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21100_ net190 _00869_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21031_ clknet_leaf_51_i_clk _00800_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19586__42 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_103_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20815_ clknet_leaf_25_i_clk _00584_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20746_ clknet_leaf_37_i_clk _00515_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20677_ clknet_leaf_3_i_clk _00461_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_104_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03293_ clknet_0__03293_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03293_
+ sky130_fd_sc_hd__clkbuf_16
X_10430_ rbzero.tex_r1\[5\] rbzero.tex_r1\[6\] _03538_ vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10361_ rbzero.tex_r1\[38\] rbzero.tex_r1\[39\] _03505_ vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ gpout0.hpos\[3\] _04855_ _04857_ _04163_ vssd1 vssd1 vccd1 vccd1 _04872_
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ _05634_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__or4_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ rbzero.color_sky\[5\] rbzero.color_floor\[5\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04806_ sky130_fd_sc_hd__mux2_1
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21229_ clknet_leaf_74_i_clk _00998_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_137_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16770_ _09114_ _08178_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__or2_1
X_13982_ _06710_ _06713_ _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a21o_1
XFILLER_74_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20306__319 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__inv_2
X_15721_ _08358_ _08365_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__xnor2_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12933_ _05650_ _05669_ _05654_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o21bai_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__or2_1
X_15652_ _08281_ _08296_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__xnor2_2
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _05577_ _05579_ _05582_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a211o_2
XFILLER_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _07206_ _07338_ _07339_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__o21ai_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _04206_ _04592_ _04314_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a21o_1
X_18371_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__xnor2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _05534_ _05536_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__nand2_1
X_15583_ _08217_ _08225_ _08227_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__o21a_1
XFILLER_42_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09891_ sky130_fd_sc_hd__and2_1
X_14534_ _07268_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__or2b_1
XFILLER_144_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11746_ rbzero.tex_g0\[15\] _04135_ _04136_ _04126_ vssd1 vssd1 vccd1 vccd1 _04524_
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17253_ _09829_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__clkbuf_1
X_14465_ _07147_ _07152_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__or2b_1
X_11677_ rbzero.debug_overlay.vplaneX\[-6\] _04420_ _04447_ vssd1 vssd1 vccd1 vccd1
+ _04456_ sky130_fd_sc_hd__and3_1
XFILLER_70_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16204_ _08778_ _08848_ vssd1 vssd1 vccd1 vccd1 _08849_ sky130_fd_sc_hd__xnor2_1
X_13416_ _05988_ _05980_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__nand2_4
XFILLER_31_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ _03653_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14396_ _07129_ _07132_ _06239_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a21oi_1
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17184_ rbzero.traced_texa\[11\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__a22o_1
XFILLER_155_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13347_ _06059_ _06060_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__and2_1
XFILLER_127_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16135_ _08743_ _08750_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__nand2_1
X_10559_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _03613_ vssd1 vssd1 vccd1 vccd1 _03617_
+ sky130_fd_sc_hd__mux2_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13278_ _05750_ _05684_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__nor2_2
XFILLER_143_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16066_ _08700_ _08709_ _08710_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__a21o_1
XFILLER_170_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12229_ net44 _04963_ _04978_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__and3_1
XFILLER_130_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15017_ _07680_ _07681_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__and2b_1
XFILLER_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19825_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__buf_4
XFILLER_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19756_ _03106_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__clkbuf_1
X_16968_ _09486_ _09495_ vssd1 vssd1 vccd1 vccd1 _09608_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18707_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__or2_1
XFILLER_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15919_ _08492_ _08494_ vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__nand2_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19687_ _03047_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20246__266 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__inv_2
X_16899_ _08985_ _09420_ vssd1 vssd1 vccd1 vccd1 _09540_ sky130_fd_sc_hd__and2_1
X_18638_ _09141_ _08423_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__nor2_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18569_ _02071_ _02172_ _02174_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a21bo_1
X_20600_ gpout2.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21580_ net501 _01349_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20531_ rbzero.texV\[7\] _03327_ _03332_ _03423_ vssd1 vssd1 vccd1 vccd1 _01403_
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20462_ _03362_ _03363_ _03364_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_4_0_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_4_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20393_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__buf_1
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21014_ clknet_leaf_68_i_clk _00783_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ _04224_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__buf_4
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _05322_ _05332_ _05320_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a21oi_1
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11531_ _04206_ _04270_ _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand3b_2
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20729_ clknet_leaf_85_i_clk _00498_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _06953_ _06959_ _06958_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__a21o_1
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11462_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__buf_4
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13201_ _05925_ _05927_ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__a21bo_1
XFILLER_99_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10413_ _03482_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__clkbuf_4
X_14181_ _06704_ _06672_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nor2_1
XFILLER_171_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11393_ gpout0.hpos\[7\] _04159_ _04171_ _04172_ vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13132_ _05820_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__nand2_1
X_10344_ rbzero.tex_r1\[46\] rbzero.tex_r1\[47\] _03494_ vssd1 vssd1 vccd1 vccd1 _03502_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13063_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__clkbuf_4
X_17940_ _01634_ _01641_ _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nand3_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ rbzero.tex_b1\[41\] rbzero.tex_b1\[40\] _04392_ vssd1 vssd1 vccd1 vccd1 _04789_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17871_ _01496_ _01511_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__nor2_1
XFILLER_61_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16822_ _09335_ _09337_ _09334_ vssd1 vssd1 vccd1 vccd1 _09464_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19541_ _02906_ _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16753_ _08383_ _08570_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__nor2_1
X_13965_ _06700_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__nand2_1
XFILLER_185_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03041_ clknet_0__03041_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03041_
+ sky130_fd_sc_hd__clkbuf_16
X_15704_ _08337_ _08347_ _08348_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__a21o_1
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12916_ rbzero.wall_tracer.visualWallDist\[7\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05653_ sky130_fd_sc_hd__a21o_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19472_ _02950_ _02951_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__nand3_1
XFILLER_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16684_ _09324_ _09326_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__xor2_1
XFILLER_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13896_ _06620_ _06631_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__nand2_1
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18423_ _02120_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__nand2_1
XFILLER_73_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ _08262_ _08278_ _08279_ vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__a21oi_2
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _05475_ _05583_ _05561_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__mux2_2
XFILLER_185_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _02044_ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__xor2_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _07894_ _05454_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__nand2_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ rbzero.debug_overlay.playerX\[4\] _05522_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_148_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19580__37 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _09874_ _09875_ vssd1 vssd1 vccd1 vccd1 _09876_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _07060_ _06843_ _07066_ _07253_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__a31o_1
X_18285_ _01860_ _01620_ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__or3_1
X_11729_ rbzero.debug_overlay.playerY\[-6\] _04475_ _04498_ _04507_ vssd1 vssd1 vccd1
+ vccd1 _04508_ sky130_fd_sc_hd__a211o_1
XFILLER_202_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15497_ _08113_ _08139_ _08140_ _08141_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__o22a_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17236_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _09814_ sky130_fd_sc_hd__nand2_1
X_14448_ _07112_ _07113_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__and2_1
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ rbzero.traced_texa\[-3\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__a22o_1
X_14379_ _06698_ _07072_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nor2_1
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _08737_ _08761_ _08762_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__a21oi_2
XFILLER_192_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _09594_ _09596_ _09592_ vssd1 vssd1 vccd1 vccd1 _09738_ sky130_fd_sc_hd__a21oi_2
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16049_ _08682_ _08689_ _08691_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__and3_1
XFILLER_130_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19808_ net52 rbzero.pov.sclk_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1 _03133_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03308_ clknet_0__03308_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03308_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19739_ _03097_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21632_ clknet_leaf_37_i_clk _01401_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21563_ net484 _01332_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20514_ _03406_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21494_ net415 _01263_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20445_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _03351_
+ sky130_fd_sc_hd__nor2_1
XFILLER_107_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20229__250 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__inv_2
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13750_ _06468_ _06482_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__xor2_1
X_10962_ rbzero.tex_b1\[11\] rbzero.tex_b1\[12\] _03828_ vssd1 vssd1 vccd1 vccd1 _03829_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ rbzero.debug_overlay.facingX\[10\] _05448_ vssd1 vssd1 vccd1 vccd1 _05449_
+ sky130_fd_sc_hd__nand2_1
X_13681_ _06394_ _06416_ _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__o21a_1
X_10893_ _03792_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15420_ rbzero.debug_overlay.playerX\[-3\] _07946_ vssd1 vssd1 vccd1 vccd1 _08065_
+ sky130_fd_sc_hd__nand2_1
X_12632_ _05383_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15351_ _07995_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__clkbuf_4
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _05315_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__or2_1
XFILLER_129_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11514_ _04292_ _04293_ _04266_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_1
X_14302_ _07036_ _07037_ _06882_ _07034_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__a211o_1
XFILLER_156_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18070_ _01632_ _01651_ _01650_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a21o_1
XFILLER_54_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12494_ rbzero.wall_tracer.trackDistY\[-6\] _05237_ rbzero.wall_tracer.trackDistY\[-7\]
+ _05238_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a221o_1
X_15282_ _07541_ _07926_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07927_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17021_ _07976_ vssd1 vssd1 vccd1 vccd1 _09661_ sky130_fd_sc_hd__clkbuf_4
X_14233_ _06944_ _06969_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__nand2_1
XFILLER_172_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11445_ _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__buf_6
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14164_ _06892_ _06899_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11376_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] rbzero.row_render.size\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__nand3_1
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13115_ _05847_ _05848_ _05851_ _05700_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a211o_2
X_10327_ rbzero.tex_r1\[54\] rbzero.tex_r1\[55\] _03483_ vssd1 vssd1 vccd1 vccd1 _03493_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14095_ _06826_ _06831_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__xor2_1
X_18972_ _02594_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13046_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__xnor2_2
XFILLER_117_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17923_ _01624_ _01625_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__xnor2_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17854_ _01556_ _01557_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16805_ _09445_ _09446_ vssd1 vssd1 vccd1 vccd1 _09447_ sky130_fd_sc_hd__xor2_1
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17785_ _01487_ _01488_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__nor2_1
X_14997_ rbzero.wall_tracer.stepDistX\[5\] _07568_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07669_ sky130_fd_sc_hd__mux2_1
XFILLER_19_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19524_ rbzero.wall_tracer.rayAddendY\[8\] rbzero.wall_tracer.rayAddendY\[7\] _02906_
+ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__o21ai_1
X_16736_ _09362_ _09377_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__xnor2_1
X_13948_ _06665_ _06670_ _06684_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__a21o_1
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19455_ _02923_ _02925_ _02935_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16667_ _09305_ _09306_ _09308_ vssd1 vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__a21o_1
X_13879_ _06273_ _06593_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__nand2_1
XFILLER_179_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18406_ _02102_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__xor2_1
X_15618_ rbzero.debug_overlay.playerX\[-9\] _08147_ _07979_ vssd1 vssd1 vccd1 vccd1
+ _08263_ sky130_fd_sc_hd__a21o_2
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19386_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__or2_1
X_16598_ _09118_ _09123_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__nand2_1
XFILLER_203_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18337_ _01756_ _01970_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__nand2_1
X_20358__367 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__inv_2
X_15549_ _08008_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_148_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18268_ _01879_ _01880_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a21bo_1
XFILLER_135_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _09779_ _09798_ _09799_ _09781_ rbzero.wall_tracer.mapX\[10\] vssd1 vssd1
+ vccd1 vccd1 _00575_ sky130_fd_sc_hd__a32o_1
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18199_ _01897_ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20161_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__buf_1
XFILLER_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20387__13 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XFILLER_66_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ clknet_leaf_51_i_clk _00763_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21615_ clknet_leaf_22_i_clk _01384_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21546_ net467 _01315_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21477_ net398 _01246_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[56\] sky130_fd_sc_hd__dfxtp_1
X_11230_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__buf_6
X_20428_ rbzero.texV\[-10\] _03175_ _03332_ _03337_ vssd1 vssd1 vccd1 vccd1 _01386_
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03044_ clknet_0__03044_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03044_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11161_ rbzero.wall_tracer.mapY\[9\] rbzero.wall_tracer.mapY\[8\] rbzero.wall_tracer.mapY\[11\]
+ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or4_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11092_ _03896_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14920_ rbzero.wall_tracer.visualWallDist\[-2\] _07618_ vssd1 vssd1 vccd1 vccd1 _07623_
+ sky130_fd_sc_hd__or2_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _05742_ _07383_ _07390_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__a2111oi_2
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13802_ _06406_ _06531_ _06530_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__nand3b_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _10133_ _10135_ vssd1 vssd1 vccd1 vccd1 _10136_ sky130_fd_sc_hd__and2_1
XFILLER_75_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ rbzero.wall_tracer.stepDistY\[-8\] _00004_ vssd1 vssd1 vccd1 vccd1 _07515_
+ sky130_fd_sc_hd__nor2_1
X_11994_ _04766_ _04767_ _04768_ _04225_ _04229_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__o221a_1
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16521_ _09164_ vssd1 vssd1 vccd1 vccd1 _09165_ sky130_fd_sc_hd__clkbuf_4
XFILLER_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13733_ _06057_ _06031_ _05945_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__o21ai_1
X_10945_ rbzero.tex_b1\[19\] rbzero.tex_b1\[20\] _03817_ vssd1 vssd1 vccd1 vccd1 _03820_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19240_ _02771_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16452_ _08821_ vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__clkbuf_4
X_13664_ _05990_ _06009_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or2_1
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10876_ _03783_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ _07486_ _07455_ _07483_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _08048_ sky130_fd_sc_hd__a211oi_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__buf_4
X_12615_ _05367_ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nand2_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _08147_ _09027_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__or2_2
X_13595_ _06148_ _06147_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__xnor2_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18122_ _01462_ _09526_ _09621_ rbzero.wall_tracer.visualWallDist\[10\] vssd1 vssd1
+ vccd1 vccd1 _01823_ sky130_fd_sc_hd__and4bb_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ rbzero.debug_overlay.playerY\[-9\] _04013_ _05196_ _07978_ vssd1 vssd1 vccd1
+ vccd1 _07979_ sky130_fd_sc_hd__o211a_2
XFILLER_40_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12546_ _05296_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__and2_1
XFILLER_200_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18053_ _01636_ _01639_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15265_ _07904_ _07909_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__nand2_1
XFILLER_184_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ _05216_ _05229_ _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o21a_1
XANTENNA_4 _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17004_ _09642_ _09643_ vssd1 vssd1 vccd1 vccd1 _09644_ sky130_fd_sc_hd__and2b_1
X_14216_ _06951_ _06952_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__nor2_1
XFILLER_125_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11428_ _04141_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__buf_4
X_15196_ _07847_ _07848_ _07833_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__o21bai_1
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14147_ _06856_ _06879_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11359_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__clkbuf_8
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14078_ _06813_ _06800_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or2b_1
X_18955_ _02607_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13029_ _05765_ _05576_ _05657_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__o21ba_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _01573_ _01608_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__nand2_1
XFILLER_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18886_ _02556_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17837_ _10233_ _10280_ _01540_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__a21boi_1
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17768_ _10074_ _10217_ _10219_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19507_ _02984_ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__nand2_1
X_16719_ _09358_ _09360_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__xor2_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17699_ _10257_ _10263_ vssd1 vssd1 vccd1 vccd1 _10264_ sky130_fd_sc_hd__xor2_2
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19438_ rbzero.wall_tracer.rayAddendY\[2\] rbzero.wall_tracer.rayAddendY\[1\] rbzero.debug_overlay.vplaneY\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03038_ _03038_ vssd1 vssd1 vccd1 vccd1 clknet_0__03038_ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19369_ _07676_ _02849_ _02850_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a31o_1
X_21400_ net321 _01169_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21331_ net252 _01100_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21262_ clknet_leaf_60_i_clk _01031_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21193_ clknet_leaf_79_i_clk _00962_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20111__144 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__inv_2
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ clknet_leaf_51_i_clk _00746_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ rbzero.tex_g0\[58\] rbzero.tex_g0\[57\] _03706_ vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ rbzero.tex_g1\[26\] rbzero.tex_g1\[27\] _03669_ vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12400_ _04154_ _03477_ _05143_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__mux2_1
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13380_ _06115_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__and3_1
XFILLER_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10592_ rbzero.tex_g1\[58\] rbzero.tex_g1\[59\] _03549_ vssd1 vssd1 vccd1 vccd1 _03634_
+ sky130_fd_sc_hd__mux2_1
XFILLER_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12331_ _05082_ _05087_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nand2_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21529_ net450 _01298_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12262_ net23 _05023_ _05026_ _05030_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__o211a_1
X_15050_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__or2_1
XFILLER_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ _06614_ _06598_ _06599_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__and3_1
X_11213_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__clkbuf_4
X_12193_ net17 net16 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__nor2_1
XFILLER_150_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11144_ rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__clkbuf_4
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 o_rgb[22] sky130_fd_sc_hd__buf_2
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18740_ _02421_ _02423_ _02422_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__o21bai_1
X_11075_ rbzero.tex_b0\[22\] rbzero.tex_b0\[21\] _03887_ vssd1 vssd1 vccd1 vccd1 _03888_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15952_ _08593_ _08595_ _08596_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__o21a_1
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20086__121 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__inv_2
X_14903_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.trackDistX\[-6\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__mux2_1
X_18671_ _02144_ _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _08527_ _08474_ vssd1 vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__xnor2_2
XFILLER_114_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17622_ _10087_ _10050_ vssd1 vssd1 vccd1 vccd1 _10187_ sky130_fd_sc_hd__or2b_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _05834_ _05800_ _07520_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__or3_1
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17553_ _10114_ _10118_ vssd1 vssd1 vccd1 vccd1 _10119_ sky130_fd_sc_hd__and2b_1
X_14765_ _07497_ _07498_ _05952_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__mux2_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _04225_ _04749_ _04750_ _04751_ _04208_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o221a_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ _09145_ _09147_ vssd1 vssd1 vccd1 vccd1 _09148_ sky130_fd_sc_hd__xor2_1
XFILLER_205_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13716_ _06441_ _06451_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__and2_1
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10928_ rbzero.tex_b1\[27\] rbzero.tex_b1\[28\] _03806_ vssd1 vssd1 vccd1 vccd1 _03811_
+ sky130_fd_sc_hd__mux2_1
X_17484_ _09938_ _09950_ _10049_ vssd1 vssd1 vccd1 vccd1 _10050_ sky130_fd_sc_hd__a21o_1
XFILLER_177_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14696_ _07375_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19223_ rbzero.spi_registers.got_new_vshift _02708_ vssd1 vssd1 vccd1 vccd1 _02761_
+ sky130_fd_sc_hd__and2_1
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16435_ _09066_ _09079_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__xor2_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _05824_ _05940_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__or2_1
X_10859_ rbzero.tex_b1\[60\] rbzero.tex_b1\[61\] _03773_ vssd1 vssd1 vccd1 vccd1 _03775_
+ sky130_fd_sc_hd__mux2_1
XFILLER_160_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19154_ rbzero.otherx\[3\] _02710_ _02717_ _02714_ vssd1 vssd1 vccd1 vccd1 _00732_
+ sky130_fd_sc_hd__o211a_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16366_ _08360_ _09009_ _09010_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__a21o_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _06101_ _06310_ _06311_ _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o22a_1
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18105_ _01698_ _01732_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__nand2_1
X_15317_ _07933_ _07530_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__o21ai_2
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19085_ rbzero.pov.spi_buffer\[73\] rbzero.pov.ready_buffer\[73\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
X_12529_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__clkbuf_4
X_16297_ _08764_ _08807_ _08941_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18036_ _08242_ _01737_ _10238_ _09552_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__or4_1
X_15248_ _07893_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__clkbuf_4
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15179_ _07820_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _07833_
+ sky130_fd_sc_hd__nor2_1
XFILLER_113_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19987_ rbzero.pov.ready_buffer\[13\] _03252_ _03253_ rbzero.debug_overlay.vplaneX\[-7\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__o221a_1
XFILLER_98_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18938_ _02598_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__clkbuf_1
.ends

