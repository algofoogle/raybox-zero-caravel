// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_outs_enb,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_spare_0,
    i_spare_1,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_outs_enb;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_spare_0;
 input i_spare_1;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire net93;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net94;
 wire net109;
 wire net110;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net127;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net111;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire _00000_;
 wire _00001_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire clknet_0__03506_;
 wire clknet_0__03507_;
 wire clknet_0__03508_;
 wire clknet_0__03509_;
 wire clknet_0__03510_;
 wire clknet_0__03511_;
 wire clknet_0__03512_;
 wire clknet_0__03513_;
 wire clknet_0__03514_;
 wire clknet_0__03840_;
 wire clknet_0__03841_;
 wire clknet_0__03842_;
 wire clknet_0__03843_;
 wire clknet_0__03844_;
 wire clknet_0__03845_;
 wire clknet_0__03846_;
 wire clknet_0__03847_;
 wire clknet_0__03848_;
 wire clknet_0__03849_;
 wire clknet_0__03850_;
 wire clknet_0__03851_;
 wire clknet_0__03852_;
 wire clknet_0__03853_;
 wire clknet_0__03854_;
 wire clknet_0__03855_;
 wire clknet_0__03856_;
 wire clknet_0__03857_;
 wire clknet_0__03858_;
 wire clknet_0__03859_;
 wire clknet_0__03860_;
 wire clknet_0__03861_;
 wire clknet_0__03862_;
 wire clknet_0__03863_;
 wire clknet_0__03864_;
 wire clknet_0__03865_;
 wire clknet_0__03866_;
 wire clknet_0__03867_;
 wire clknet_0__03868_;
 wire clknet_0__03869_;
 wire clknet_0__03870_;
 wire clknet_0__03871_;
 wire clknet_0__03872_;
 wire clknet_0__05645_;
 wire clknet_0__05688_;
 wire clknet_0__05742_;
 wire clknet_0__05794_;
 wire clknet_0__05847_;
 wire clknet_0__05898_;
 wire clknet_0__05946_;
 wire clknet_0_i_clk;
 wire clknet_1_0__leaf__03506_;
 wire clknet_1_0__leaf__03507_;
 wire clknet_1_0__leaf__03508_;
 wire clknet_1_0__leaf__03509_;
 wire clknet_1_0__leaf__03510_;
 wire clknet_1_0__leaf__03511_;
 wire clknet_1_0__leaf__03512_;
 wire clknet_1_0__leaf__03513_;
 wire clknet_1_0__leaf__03514_;
 wire clknet_1_0__leaf__03840_;
 wire clknet_1_0__leaf__03841_;
 wire clknet_1_0__leaf__03842_;
 wire clknet_1_0__leaf__03843_;
 wire clknet_1_0__leaf__03844_;
 wire clknet_1_0__leaf__03845_;
 wire clknet_1_0__leaf__03846_;
 wire clknet_1_0__leaf__03847_;
 wire clknet_1_0__leaf__03848_;
 wire clknet_1_0__leaf__03849_;
 wire clknet_1_0__leaf__03850_;
 wire clknet_1_0__leaf__03851_;
 wire clknet_1_0__leaf__03852_;
 wire clknet_1_0__leaf__03853_;
 wire clknet_1_0__leaf__03854_;
 wire clknet_1_0__leaf__03855_;
 wire clknet_1_0__leaf__03856_;
 wire clknet_1_0__leaf__03857_;
 wire clknet_1_0__leaf__03858_;
 wire clknet_1_0__leaf__03859_;
 wire clknet_1_0__leaf__03860_;
 wire clknet_1_0__leaf__03861_;
 wire clknet_1_0__leaf__03862_;
 wire clknet_1_0__leaf__03863_;
 wire clknet_1_0__leaf__03864_;
 wire clknet_1_0__leaf__03865_;
 wire clknet_1_0__leaf__03866_;
 wire clknet_1_0__leaf__03867_;
 wire clknet_1_0__leaf__03868_;
 wire clknet_1_0__leaf__03869_;
 wire clknet_1_0__leaf__03870_;
 wire clknet_1_0__leaf__03871_;
 wire clknet_1_0__leaf__03872_;
 wire clknet_1_0__leaf__05645_;
 wire clknet_1_0__leaf__05688_;
 wire clknet_1_0__leaf__05742_;
 wire clknet_1_0__leaf__05794_;
 wire clknet_1_0__leaf__05847_;
 wire clknet_1_0__leaf__05898_;
 wire clknet_1_0__leaf__05946_;
 wire clknet_1_1__leaf__03506_;
 wire clknet_1_1__leaf__03507_;
 wire clknet_1_1__leaf__03508_;
 wire clknet_1_1__leaf__03509_;
 wire clknet_1_1__leaf__03510_;
 wire clknet_1_1__leaf__03511_;
 wire clknet_1_1__leaf__03512_;
 wire clknet_1_1__leaf__03513_;
 wire clknet_1_1__leaf__03514_;
 wire clknet_1_1__leaf__03840_;
 wire clknet_1_1__leaf__03841_;
 wire clknet_1_1__leaf__03842_;
 wire clknet_1_1__leaf__03843_;
 wire clknet_1_1__leaf__03844_;
 wire clknet_1_1__leaf__03845_;
 wire clknet_1_1__leaf__03846_;
 wire clknet_1_1__leaf__03847_;
 wire clknet_1_1__leaf__03848_;
 wire clknet_1_1__leaf__03849_;
 wire clknet_1_1__leaf__03850_;
 wire clknet_1_1__leaf__03851_;
 wire clknet_1_1__leaf__03852_;
 wire clknet_1_1__leaf__03853_;
 wire clknet_1_1__leaf__03854_;
 wire clknet_1_1__leaf__03855_;
 wire clknet_1_1__leaf__03856_;
 wire clknet_1_1__leaf__03857_;
 wire clknet_1_1__leaf__03858_;
 wire clknet_1_1__leaf__03859_;
 wire clknet_1_1__leaf__03860_;
 wire clknet_1_1__leaf__03861_;
 wire clknet_1_1__leaf__03862_;
 wire clknet_1_1__leaf__03863_;
 wire clknet_1_1__leaf__03864_;
 wire clknet_1_1__leaf__03865_;
 wire clknet_1_1__leaf__03866_;
 wire clknet_1_1__leaf__03867_;
 wire clknet_1_1__leaf__03868_;
 wire clknet_1_1__leaf__03869_;
 wire clknet_1_1__leaf__03870_;
 wire clknet_1_1__leaf__03871_;
 wire clknet_1_1__leaf__03872_;
 wire clknet_1_1__leaf__05645_;
 wire clknet_1_1__leaf__05688_;
 wire clknet_1_1__leaf__05742_;
 wire clknet_1_1__leaf__05794_;
 wire clknet_1_1__leaf__05847_;
 wire clknet_1_1__leaf__05898_;
 wire clknet_1_1__leaf__05946_;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_4_0__leaf_i_clk;
 wire clknet_4_10__leaf_i_clk;
 wire clknet_4_11__leaf_i_clk;
 wire clknet_4_12__leaf_i_clk;
 wire clknet_4_13__leaf_i_clk;
 wire clknet_4_14__leaf_i_clk;
 wire clknet_4_15__leaf_i_clk;
 wire clknet_4_1__leaf_i_clk;
 wire clknet_4_2__leaf_i_clk;
 wire clknet_4_3__leaf_i_clk;
 wire clknet_4_4__leaf_i_clk;
 wire clknet_4_5__leaf_i_clk;
 wire clknet_4_6__leaf_i_clk;
 wire clknet_4_7__leaf_i_clk;
 wire clknet_4_8__leaf_i_clk;
 wire clknet_4_9__leaf_i_clk;
 wire clknet_leaf_0_i_clk;
 wire clknet_leaf_100_i_clk;
 wire clknet_leaf_101_i_clk;
 wire clknet_leaf_102_i_clk;
 wire clknet_leaf_103_i_clk;
 wire clknet_leaf_104_i_clk;
 wire clknet_leaf_105_i_clk;
 wire clknet_leaf_106_i_clk;
 wire clknet_leaf_107_i_clk;
 wire clknet_leaf_108_i_clk;
 wire clknet_leaf_109_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_110_i_clk;
 wire clknet_leaf_111_i_clk;
 wire clknet_leaf_112_i_clk;
 wire clknet_leaf_113_i_clk;
 wire clknet_leaf_114_i_clk;
 wire clknet_leaf_115_i_clk;
 wire clknet_leaf_116_i_clk;
 wire clknet_leaf_117_i_clk;
 wire clknet_leaf_118_i_clk;
 wire clknet_leaf_119_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_120_i_clk;
 wire clknet_leaf_121_i_clk;
 wire clknet_leaf_122_i_clk;
 wire clknet_leaf_123_i_clk;
 wire clknet_leaf_124_i_clk;
 wire clknet_leaf_125_i_clk;
 wire clknet_leaf_126_i_clk;
 wire clknet_leaf_127_i_clk;
 wire clknet_leaf_128_i_clk;
 wire clknet_leaf_129_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_130_i_clk;
 wire clknet_leaf_131_i_clk;
 wire clknet_leaf_132_i_clk;
 wire clknet_leaf_133_i_clk;
 wire clknet_leaf_134_i_clk;
 wire clknet_leaf_135_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_9_i_clk;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net1;
 wire net10;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net247;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net249;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net254;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net256;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net259;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net26;
 wire net260;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net263;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net264;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net268;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net269;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net274;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net297;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net298;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net303;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net304;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net305;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net306;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net31;
 wire net310;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net311;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net315;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net317;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net324;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net325;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net329;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net33;
 wire net330;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net332;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net336;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net339;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net342;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net344;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net345;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net346;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net354;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net355;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net356;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net357;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net358;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net359;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net360;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net361;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net362;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net363;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net364;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net365;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net366;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net367;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net368;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net369;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net37;
 wire net370;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net371;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net372;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net373;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net374;
 wire net3740;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net375;
 wire net3750;
 wire net3751;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3759;
 wire net376;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net377;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net378;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net379;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net38;
 wire net380;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net381;
 wire net3810;
 wire net3811;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net382;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3828;
 wire net3829;
 wire net383;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net384;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net385;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net386;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net387;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net388;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net389;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net39;
 wire net390;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net391;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net392;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net393;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net394;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net395;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net396;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net397;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net398;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net399;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4;
 wire net40;
 wire net400;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net401;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net402;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net403;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net404;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net405;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net406;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net407;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net408;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net409;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net41;
 wire net410;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net411;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net412;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net413;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net414;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net415;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net416;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net417;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net418;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net419;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net42;
 wire net420;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net421;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net422;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net423;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net424;
 wire net4240;
 wire net4241;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net425;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net426;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net427;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net428;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4288;
 wire net4289;
 wire net429;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net43;
 wire net430;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net431;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4319;
 wire net432;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net433;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net434;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net435;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net436;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net437;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net438;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net439;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net44;
 wire net440;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net441;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net442;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net443;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net444;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net445;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net446;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net447;
 wire net4470;
 wire net4471;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net448;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net449;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net45;
 wire net450;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net451;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net452;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net453;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net454;
 wire net4540;
 wire net4541;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net455;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net456;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net457;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net458;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net459;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net46;
 wire net460;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net461;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net462;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net463;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net464;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net465;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net466;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net467;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4679;
 wire net468;
 wire net4680;
 wire net4681;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net469;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net47;
 wire net470;
 wire net4700;
 wire net4701;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net471;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net472;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net473;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net474;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net475;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net476;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net477;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net478;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net479;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net48;
 wire net480;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net481;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net482;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net483;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net484;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net485;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net486;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net487;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net488;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net489;
 wire net4890;
 wire net4891;
 wire net4893;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net49;
 wire net490;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net491;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net492;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net493;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net494;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net495;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net496;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net497;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net498;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net499;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5;
 wire net50;
 wire net500;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net501;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net502;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net503;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net504;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net505;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net506;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net507;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net508;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net509;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net51;
 wire net510;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net511;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net512;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net513;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net514;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net515;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net516;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net517;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net518;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net519;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net52;
 wire net520;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net521;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net522;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net523;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net524;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net525;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net526;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net527;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net528;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net529;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net53;
 wire net530;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net531;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net532;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net533;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net534;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net535;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net536;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net537;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net538;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net539;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net54;
 wire net540;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net541;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net542;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net543;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net544;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net545;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net546;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net547;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net548;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net549;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net55;
 wire net550;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net551;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net552;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net553;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net554;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net555;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net556;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net557;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net558;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net559;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net56;
 wire net560;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net561;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net562;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net563;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net564;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net565;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net566;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net567;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net568;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net569;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net57;
 wire net570;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net571;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net572;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net573;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net574;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net575;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net576;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net577;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net578;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net579;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net58;
 wire net580;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5808;
 wire net5809;
 wire net581;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net582;
 wire net5820;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net583;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net584;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net585;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net586;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net587;
 wire net5870;
 wire net5871;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net588;
 wire net5880;
 wire net5881;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net589;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net59;
 wire net590;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net591;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net592;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net593;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net594;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net595;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net596;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net597;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net598;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net599;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6;
 wire net60;
 wire net600;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net601;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net602;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net603;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net604;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net605;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net606;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net607;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net608;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net609;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net61;
 wire net610;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net611;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net612;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net613;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net614;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net615;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net616;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net617;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net618;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net619;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net62;
 wire net620;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net621;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net622;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net623;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net624;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net625;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net626;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net627;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net628;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net629;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net63;
 wire net630;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net631;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net632;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net633;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net634;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net635;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net636;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net637;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net638;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net639;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net64;
 wire net640;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net641;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net642;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net643;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net644;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net645;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net646;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net647;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net648;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net649;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net65;
 wire net650;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net651;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net652;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net653;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net654;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net655;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net656;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net657;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net658;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net659;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net66;
 wire net660;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net661;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net662;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net663;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net664;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net665;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net666;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net667;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net668;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net669;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net67;
 wire net670;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net671;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net672;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net673;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net674;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net675;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net676;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net677;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net678;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net679;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net68;
 wire net680;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net681;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net682;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net683;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net684;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net685;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net686;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net687;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net688;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net689;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net69;
 wire net690;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net691;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net692;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net693;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net694;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net695;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net696;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net697;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net698;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net6988;
 wire net6989;
 wire net699;
 wire net6990;
 wire net6991;
 wire net6992;
 wire net6993;
 wire net6994;
 wire net6995;
 wire net6996;
 wire net6997;
 wire net6998;
 wire net6999;
 wire net7;
 wire net70;
 wire net700;
 wire net7000;
 wire net7001;
 wire net7002;
 wire net7003;
 wire net7004;
 wire net7005;
 wire net7006;
 wire net7007;
 wire net7008;
 wire net7009;
 wire net701;
 wire net7010;
 wire net7011;
 wire net7012;
 wire net7013;
 wire net7014;
 wire net7015;
 wire net7016;
 wire net7017;
 wire net7018;
 wire net7019;
 wire net702;
 wire net7020;
 wire net7021;
 wire net7022;
 wire net7023;
 wire net7024;
 wire net7025;
 wire net7026;
 wire net7027;
 wire net7028;
 wire net7029;
 wire net703;
 wire net7030;
 wire net7031;
 wire net7032;
 wire net7033;
 wire net7034;
 wire net7035;
 wire net7036;
 wire net7037;
 wire net7038;
 wire net7039;
 wire net704;
 wire net7040;
 wire net7041;
 wire net7042;
 wire net7043;
 wire net7044;
 wire net7045;
 wire net7046;
 wire net7047;
 wire net7048;
 wire net7049;
 wire net705;
 wire net7050;
 wire net7051;
 wire net7052;
 wire net7053;
 wire net7054;
 wire net7055;
 wire net7056;
 wire net7057;
 wire net7058;
 wire net7059;
 wire net706;
 wire net7060;
 wire net7061;
 wire net7062;
 wire net7063;
 wire net7064;
 wire net7065;
 wire net7066;
 wire net7067;
 wire net7068;
 wire net7069;
 wire net707;
 wire net7070;
 wire net7071;
 wire net7072;
 wire net7073;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7077;
 wire net7078;
 wire net7079;
 wire net708;
 wire net7080;
 wire net7081;
 wire net7082;
 wire net7083;
 wire net7084;
 wire net7085;
 wire net7086;
 wire net7087;
 wire net7088;
 wire net7089;
 wire net709;
 wire net7090;
 wire net7091;
 wire net7092;
 wire net7093;
 wire net7094;
 wire net7095;
 wire net7096;
 wire net7097;
 wire net7098;
 wire net7099;
 wire net71;
 wire net710;
 wire net7100;
 wire net7101;
 wire net7102;
 wire net7103;
 wire net7104;
 wire net7105;
 wire net7106;
 wire net7107;
 wire net7108;
 wire net7109;
 wire net711;
 wire net7110;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7115;
 wire net7116;
 wire net7117;
 wire net7118;
 wire net7119;
 wire net712;
 wire net7120;
 wire net7121;
 wire net7122;
 wire net7123;
 wire net7124;
 wire net7125;
 wire net7126;
 wire net7127;
 wire net7128;
 wire net7129;
 wire net713;
 wire net7130;
 wire net7131;
 wire net7132;
 wire net7133;
 wire net7134;
 wire net7135;
 wire net7136;
 wire net7137;
 wire net7138;
 wire net7139;
 wire net714;
 wire net7140;
 wire net7141;
 wire net7142;
 wire net7143;
 wire net7144;
 wire net7145;
 wire net7146;
 wire net7147;
 wire net7148;
 wire net7149;
 wire net715;
 wire net7150;
 wire net7151;
 wire net7152;
 wire net7153;
 wire net7154;
 wire net7155;
 wire net7156;
 wire net7157;
 wire net7158;
 wire net7159;
 wire net716;
 wire net7160;
 wire net7161;
 wire net7162;
 wire net7163;
 wire net7164;
 wire net7165;
 wire net7166;
 wire net7167;
 wire net7168;
 wire net7169;
 wire net717;
 wire net7170;
 wire net7171;
 wire net7172;
 wire net7173;
 wire net7174;
 wire net7175;
 wire net7176;
 wire net7177;
 wire net7178;
 wire net7179;
 wire net718;
 wire net7180;
 wire net7181;
 wire net7182;
 wire net7183;
 wire net7184;
 wire net7185;
 wire net7186;
 wire net7187;
 wire net7188;
 wire net7189;
 wire net719;
 wire net7190;
 wire net7191;
 wire net7192;
 wire net7193;
 wire net7194;
 wire net7195;
 wire net7196;
 wire net7197;
 wire net7198;
 wire net7199;
 wire net72;
 wire net720;
 wire net7200;
 wire net7201;
 wire net7202;
 wire net7203;
 wire net7204;
 wire net7205;
 wire net7206;
 wire net7207;
 wire net7208;
 wire net7209;
 wire net721;
 wire net7210;
 wire net7211;
 wire net7212;
 wire net7213;
 wire net7214;
 wire net7215;
 wire net7216;
 wire net7217;
 wire net7218;
 wire net7219;
 wire net722;
 wire net7220;
 wire net7221;
 wire net7222;
 wire net7223;
 wire net7224;
 wire net7225;
 wire net7226;
 wire net7227;
 wire net7228;
 wire net7229;
 wire net723;
 wire net7230;
 wire net7231;
 wire net7232;
 wire net7233;
 wire net7234;
 wire net7235;
 wire net7236;
 wire net7237;
 wire net7238;
 wire net7239;
 wire net724;
 wire net7240;
 wire net7241;
 wire net7242;
 wire net7243;
 wire net7244;
 wire net7245;
 wire net7246;
 wire net7247;
 wire net7248;
 wire net7249;
 wire net725;
 wire net7250;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7254;
 wire net7255;
 wire net7256;
 wire net7257;
 wire net7258;
 wire net7259;
 wire net726;
 wire net7260;
 wire net7261;
 wire net7262;
 wire net7263;
 wire net7264;
 wire net7265;
 wire net7266;
 wire net7267;
 wire net7268;
 wire net7269;
 wire net727;
 wire net7270;
 wire net7271;
 wire net7272;
 wire net7273;
 wire net7274;
 wire net7275;
 wire net7276;
 wire net7277;
 wire net7278;
 wire net7279;
 wire net728;
 wire net7280;
 wire net7281;
 wire net7282;
 wire net7283;
 wire net7284;
 wire net7285;
 wire net7286;
 wire net7287;
 wire net7288;
 wire net7289;
 wire net729;
 wire net7290;
 wire net7291;
 wire net7292;
 wire net7293;
 wire net7294;
 wire net7295;
 wire net7296;
 wire net7297;
 wire net7298;
 wire net7299;
 wire net73;
 wire net730;
 wire net7300;
 wire net7301;
 wire net7302;
 wire net7303;
 wire net7304;
 wire net7305;
 wire net7306;
 wire net7307;
 wire net7308;
 wire net7309;
 wire net731;
 wire net7310;
 wire net7311;
 wire net7312;
 wire net7313;
 wire net7314;
 wire net7315;
 wire net7316;
 wire net7317;
 wire net7318;
 wire net7319;
 wire net732;
 wire net7320;
 wire net7321;
 wire net7322;
 wire net7323;
 wire net7324;
 wire net7325;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net733;
 wire net7330;
 wire net7331;
 wire net7332;
 wire net7333;
 wire net7334;
 wire net7335;
 wire net7336;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net734;
 wire net7340;
 wire net7341;
 wire net7342;
 wire net7343;
 wire net7344;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7348;
 wire net7349;
 wire net735;
 wire net7350;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net736;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net737;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net738;
 wire net7380;
 wire net7381;
 wire net7382;
 wire net7383;
 wire net7384;
 wire net7385;
 wire net7386;
 wire net7387;
 wire net7388;
 wire net7389;
 wire net739;
 wire net7390;
 wire net7391;
 wire net7392;
 wire net7393;
 wire net7394;
 wire net7395;
 wire net7396;
 wire net7397;
 wire net7398;
 wire net7399;
 wire net74;
 wire net740;
 wire net7400;
 wire net7401;
 wire net7402;
 wire net7403;
 wire net7404;
 wire net7405;
 wire net7406;
 wire net7407;
 wire net7408;
 wire net7409;
 wire net741;
 wire net7410;
 wire net7411;
 wire net7412;
 wire net7413;
 wire net7414;
 wire net7415;
 wire net7416;
 wire net7417;
 wire net7418;
 wire net7419;
 wire net742;
 wire net7420;
 wire net7421;
 wire net7422;
 wire net7423;
 wire net7424;
 wire net7425;
 wire net7426;
 wire net7427;
 wire net7428;
 wire net7429;
 wire net743;
 wire net7430;
 wire net7431;
 wire net7432;
 wire net7433;
 wire net7434;
 wire net7435;
 wire net7436;
 wire net7437;
 wire net7438;
 wire net7439;
 wire net744;
 wire net7440;
 wire net7441;
 wire net7442;
 wire net7443;
 wire net7444;
 wire net7445;
 wire net7446;
 wire net7447;
 wire net7448;
 wire net7449;
 wire net745;
 wire net7450;
 wire net7451;
 wire net7452;
 wire net7453;
 wire net7454;
 wire net7455;
 wire net7456;
 wire net7457;
 wire net7458;
 wire net7459;
 wire net746;
 wire net7460;
 wire net7461;
 wire net7462;
 wire net7463;
 wire net7464;
 wire net7465;
 wire net7466;
 wire net7467;
 wire net7468;
 wire net7469;
 wire net747;
 wire net7470;
 wire net7471;
 wire net7472;
 wire net7473;
 wire net7474;
 wire net7475;
 wire net7476;
 wire net7477;
 wire net7478;
 wire net7479;
 wire net748;
 wire net7480;
 wire net7481;
 wire net7482;
 wire net7483;
 wire net7484;
 wire net7485;
 wire net7486;
 wire net7487;
 wire net7488;
 wire net7489;
 wire net749;
 wire net7490;
 wire net7491;
 wire net7492;
 wire net7493;
 wire net7494;
 wire net7495;
 wire net7496;
 wire net7497;
 wire net7498;
 wire net7499;
 wire net75;
 wire net750;
 wire net7500;
 wire net7501;
 wire net7502;
 wire net7503;
 wire net7504;
 wire net7505;
 wire net7506;
 wire net7507;
 wire net7508;
 wire net7509;
 wire net751;
 wire net7510;
 wire net7511;
 wire net7512;
 wire net7513;
 wire net7514;
 wire net7515;
 wire net7516;
 wire net7517;
 wire net7518;
 wire net7519;
 wire net752;
 wire net7520;
 wire net7521;
 wire net7522;
 wire net7523;
 wire net7524;
 wire net7525;
 wire net7526;
 wire net7527;
 wire net7528;
 wire net7529;
 wire net753;
 wire net7530;
 wire net7531;
 wire net7532;
 wire net7533;
 wire net7534;
 wire net7535;
 wire net7536;
 wire net7537;
 wire net7538;
 wire net7539;
 wire net754;
 wire net7540;
 wire net7541;
 wire net7542;
 wire net7543;
 wire net7544;
 wire net7545;
 wire net7546;
 wire net7547;
 wire net7548;
 wire net7549;
 wire net755;
 wire net7550;
 wire net7551;
 wire net7552;
 wire net7553;
 wire net7554;
 wire net7555;
 wire net7556;
 wire net7557;
 wire net7558;
 wire net7559;
 wire net756;
 wire net7560;
 wire net7561;
 wire net7562;
 wire net7563;
 wire net7564;
 wire net7565;
 wire net7566;
 wire net7567;
 wire net7568;
 wire net7569;
 wire net757;
 wire net7570;
 wire net7571;
 wire net7572;
 wire net7573;
 wire net7574;
 wire net7575;
 wire net7576;
 wire net7577;
 wire net7578;
 wire net7579;
 wire net758;
 wire net7580;
 wire net7581;
 wire net7582;
 wire net7583;
 wire net7584;
 wire net7585;
 wire net7586;
 wire net7587;
 wire net7588;
 wire net7589;
 wire net759;
 wire net7590;
 wire net7591;
 wire net7592;
 wire net7593;
 wire net7594;
 wire net7595;
 wire net7596;
 wire net7597;
 wire net7598;
 wire net7599;
 wire net76;
 wire net760;
 wire net7600;
 wire net7601;
 wire net7602;
 wire net7603;
 wire net7604;
 wire net7605;
 wire net7606;
 wire net7607;
 wire net7608;
 wire net7609;
 wire net761;
 wire net7610;
 wire net7611;
 wire net7612;
 wire net7613;
 wire net7614;
 wire net7615;
 wire net7616;
 wire net7617;
 wire net7618;
 wire net7619;
 wire net762;
 wire net7620;
 wire net7621;
 wire net7623;
 wire net7624;
 wire net7626;
 wire net7627;
 wire net7628;
 wire net7629;
 wire net763;
 wire net7630;
 wire net7631;
 wire net7632;
 wire net7633;
 wire net7634;
 wire net7635;
 wire net7636;
 wire net7637;
 wire net7639;
 wire net764;
 wire net7640;
 wire net7642;
 wire net7643;
 wire net7645;
 wire net7646;
 wire net7647;
 wire net7648;
 wire net7649;
 wire net765;
 wire net7650;
 wire net7652;
 wire net7653;
 wire net7654;
 wire net7655;
 wire net7656;
 wire net7657;
 wire net7659;
 wire net766;
 wire net7660;
 wire net7662;
 wire net7663;
 wire net7664;
 wire net7665;
 wire net7666;
 wire net7667;
 wire net7668;
 wire net7669;
 wire net767;
 wire net7670;
 wire net7671;
 wire net7672;
 wire net7673;
 wire net7674;
 wire net7675;
 wire net7676;
 wire net7677;
 wire net7678;
 wire net7679;
 wire net768;
 wire net7680;
 wire net7681;
 wire net7682;
 wire net7683;
 wire net7684;
 wire net7685;
 wire net7686;
 wire net7687;
 wire net7688;
 wire net7689;
 wire net769;
 wire net7690;
 wire net7691;
 wire net7692;
 wire net7693;
 wire net7694;
 wire net7695;
 wire net7696;
 wire net7697;
 wire net7698;
 wire net7699;
 wire net77;
 wire net770;
 wire net7700;
 wire net7701;
 wire net7702;
 wire net7703;
 wire net7704;
 wire net7705;
 wire net7706;
 wire net7707;
 wire net7708;
 wire net7709;
 wire net771;
 wire net7710;
 wire net7711;
 wire net7712;
 wire net7713;
 wire net7714;
 wire net7715;
 wire net7716;
 wire net7717;
 wire net7718;
 wire net7719;
 wire net772;
 wire net7720;
 wire net7721;
 wire net7722;
 wire net7723;
 wire net7724;
 wire net7725;
 wire net7726;
 wire net7727;
 wire net7728;
 wire net7729;
 wire net773;
 wire net7730;
 wire net7731;
 wire net7732;
 wire net7733;
 wire net7734;
 wire net7735;
 wire net7736;
 wire net7737;
 wire net7738;
 wire net7739;
 wire net774;
 wire net7741;
 wire net7742;
 wire net7743;
 wire net7744;
 wire net7745;
 wire net7746;
 wire net7747;
 wire net7748;
 wire net7749;
 wire net775;
 wire net7750;
 wire net7751;
 wire net7752;
 wire net776;
 wire net7763;
 wire net7764;
 wire net7765;
 wire net7766;
 wire net7767;
 wire net7768;
 wire net7769;
 wire net777;
 wire net7770;
 wire net7771;
 wire net7772;
 wire net7775;
 wire net7776;
 wire net7777;
 wire net7778;
 wire net7779;
 wire net778;
 wire net7780;
 wire net7781;
 wire net7783;
 wire net7784;
 wire net7785;
 wire net7786;
 wire net7787;
 wire net7788;
 wire net7789;
 wire net779;
 wire net7793;
 wire net7794;
 wire net7795;
 wire net7796;
 wire net7797;
 wire net7798;
 wire net7799;
 wire net78;
 wire net780;
 wire net7805;
 wire net7806;
 wire net7807;
 wire net7808;
 wire net7809;
 wire net781;
 wire net7810;
 wire net7811;
 wire net7812;
 wire net7813;
 wire net7814;
 wire net7815;
 wire net7816;
 wire net7817;
 wire net7818;
 wire net782;
 wire net7821;
 wire net7823;
 wire net7824;
 wire net7825;
 wire net7826;
 wire net7827;
 wire net783;
 wire net7830;
 wire net7831;
 wire net7832;
 wire net7833;
 wire net7835;
 wire net7836;
 wire net7837;
 wire net7839;
 wire net784;
 wire net7840;
 wire net7841;
 wire net7842;
 wire net7843;
 wire net7845;
 wire net7846;
 wire net7847;
 wire net7848;
 wire net785;
 wire net7850;
 wire net7851;
 wire net7852;
 wire net7853;
 wire net7854;
 wire net7855;
 wire net7856;
 wire net7857;
 wire net7858;
 wire net786;
 wire net7861;
 wire net7862;
 wire net7863;
 wire net7866;
 wire net7867;
 wire net7868;
 wire net7869;
 wire net787;
 wire net7870;
 wire net7871;
 wire net7872;
 wire net7873;
 wire net7874;
 wire net7875;
 wire net7876;
 wire net7877;
 wire net7878;
 wire net7879;
 wire net788;
 wire net7880;
 wire net7881;
 wire net7882;
 wire net7883;
 wire net7884;
 wire net7885;
 wire net7886;
 wire net7887;
 wire net7888;
 wire net7889;
 wire net789;
 wire net7890;
 wire net7891;
 wire net7892;
 wire net7893;
 wire net7894;
 wire net7895;
 wire net7896;
 wire net7897;
 wire net7898;
 wire net7899;
 wire net79;
 wire net790;
 wire net7900;
 wire net7901;
 wire net7902;
 wire net7903;
 wire net7904;
 wire net7905;
 wire net7906;
 wire net7907;
 wire net7908;
 wire net7909;
 wire net791;
 wire net7910;
 wire net7912;
 wire net7913;
 wire net7914;
 wire net7915;
 wire net7916;
 wire net7917;
 wire net7918;
 wire net7919;
 wire net792;
 wire net7921;
 wire net7922;
 wire net7923;
 wire net7925;
 wire net7926;
 wire net7927;
 wire net7928;
 wire net7929;
 wire net793;
 wire net7930;
 wire net7931;
 wire net7933;
 wire net7934;
 wire net7935;
 wire net7936;
 wire net7937;
 wire net7938;
 wire net7939;
 wire net794;
 wire net7940;
 wire net7941;
 wire net7942;
 wire net7945;
 wire net7946;
 wire net7947;
 wire net7948;
 wire net7949;
 wire net795;
 wire net7950;
 wire net7951;
 wire net7952;
 wire net7953;
 wire net7954;
 wire net7955;
 wire net7956;
 wire net7957;
 wire net7958;
 wire net7959;
 wire net796;
 wire net7960;
 wire net7961;
 wire net7962;
 wire net7963;
 wire net7964;
 wire net7965;
 wire net7966;
 wire net7967;
 wire net7968;
 wire net7969;
 wire net797;
 wire net7970;
 wire net7971;
 wire net7972;
 wire net7973;
 wire net7974;
 wire net7975;
 wire net7976;
 wire net7977;
 wire net7978;
 wire net7979;
 wire net798;
 wire net7980;
 wire net7981;
 wire net7982;
 wire net7983;
 wire net7984;
 wire net7985;
 wire net7986;
 wire net7987;
 wire net7988;
 wire net7989;
 wire net799;
 wire net7990;
 wire net7991;
 wire net7992;
 wire net7993;
 wire net7994;
 wire net7995;
 wire net7996;
 wire net7997;
 wire net7998;
 wire net7999;
 wire net8;
 wire net80;
 wire net800;
 wire net8000;
 wire net8001;
 wire net8002;
 wire net8003;
 wire net8004;
 wire net8005;
 wire net8006;
 wire net8007;
 wire net8008;
 wire net8009;
 wire net801;
 wire net8010;
 wire net8011;
 wire net8012;
 wire net8013;
 wire net8014;
 wire net8015;
 wire net8016;
 wire net8017;
 wire net8018;
 wire net8019;
 wire net802;
 wire net8020;
 wire net8021;
 wire net8022;
 wire net8023;
 wire net8025;
 wire net8026;
 wire net8027;
 wire net8028;
 wire net8029;
 wire net803;
 wire net8030;
 wire net8031;
 wire net8033;
 wire net8034;
 wire net8035;
 wire net8036;
 wire net8037;
 wire net8038;
 wire net8039;
 wire net804;
 wire net8041;
 wire net8042;
 wire net8044;
 wire net8045;
 wire net8047;
 wire net8048;
 wire net8049;
 wire net805;
 wire net8050;
 wire net8051;
 wire net8052;
 wire net8053;
 wire net8055;
 wire net8056;
 wire net8057;
 wire net8058;
 wire net806;
 wire net8060;
 wire net8061;
 wire net8062;
 wire net8063;
 wire net8065;
 wire net8066;
 wire net8067;
 wire net8068;
 wire net8069;
 wire net807;
 wire net8070;
 wire net8071;
 wire net8072;
 wire net8074;
 wire net8075;
 wire net8076;
 wire net8077;
 wire net8078;
 wire net8079;
 wire net808;
 wire net8080;
 wire net8081;
 wire net8082;
 wire net8084;
 wire net8085;
 wire net8086;
 wire net8087;
 wire net8088;
 wire net8089;
 wire net809;
 wire net8090;
 wire net8092;
 wire net8093;
 wire net8094;
 wire net8095;
 wire net8096;
 wire net8097;
 wire net8098;
 wire net8099;
 wire net81;
 wire net810;
 wire net8100;
 wire net8101;
 wire net8102;
 wire net8103;
 wire net8104;
 wire net8105;
 wire net8106;
 wire net8108;
 wire net8109;
 wire net811;
 wire net8110;
 wire net8112;
 wire net8113;
 wire net8114;
 wire net8115;
 wire net8116;
 wire net8117;
 wire net8118;
 wire net8119;
 wire net812;
 wire net8120;
 wire net8121;
 wire net8122;
 wire net8123;
 wire net8124;
 wire net8125;
 wire net8126;
 wire net8127;
 wire net8128;
 wire net8129;
 wire net813;
 wire net8130;
 wire net8131;
 wire net8132;
 wire net8133;
 wire net8134;
 wire net8135;
 wire net8136;
 wire net8137;
 wire net8138;
 wire net8139;
 wire net814;
 wire net8140;
 wire net8141;
 wire net8142;
 wire net8143;
 wire net8144;
 wire net8145;
 wire net8146;
 wire net8147;
 wire net8148;
 wire net8149;
 wire net815;
 wire net8150;
 wire net8151;
 wire net8152;
 wire net8153;
 wire net8154;
 wire net8155;
 wire net8156;
 wire net8157;
 wire net8158;
 wire net8159;
 wire net816;
 wire net8160;
 wire net8161;
 wire net8162;
 wire net8163;
 wire net8164;
 wire net8165;
 wire net8166;
 wire net8167;
 wire net8168;
 wire net8169;
 wire net817;
 wire net8170;
 wire net8171;
 wire net8172;
 wire net8173;
 wire net8174;
 wire net8175;
 wire net8177;
 wire net8179;
 wire net818;
 wire net8180;
 wire net8181;
 wire net8182;
 wire net8184;
 wire net8186;
 wire net8188;
 wire net819;
 wire net8190;
 wire net8191;
 wire net8192;
 wire net8193;
 wire net8194;
 wire net8195;
 wire net8196;
 wire net8197;
 wire net8198;
 wire net8199;
 wire net82;
 wire net820;
 wire net8200;
 wire net8202;
 wire net8203;
 wire net8205;
 wire net8206;
 wire net8207;
 wire net8208;
 wire net8209;
 wire net821;
 wire net8210;
 wire net8212;
 wire net8213;
 wire net8214;
 wire net8215;
 wire net8216;
 wire net8217;
 wire net8218;
 wire net8219;
 wire net822;
 wire net8220;
 wire net8221;
 wire net8222;
 wire net8223;
 wire net8224;
 wire net8225;
 wire net8226;
 wire net8227;
 wire net8228;
 wire net8229;
 wire net823;
 wire net8230;
 wire net8231;
 wire net8232;
 wire net8233;
 wire net8234;
 wire net8235;
 wire net8236;
 wire net8238;
 wire net824;
 wire net8240;
 wire net8241;
 wire net8242;
 wire net8243;
 wire net8244;
 wire net8245;
 wire net8246;
 wire net8247;
 wire net8248;
 wire net8249;
 wire net825;
 wire net8250;
 wire net8251;
 wire net8252;
 wire net8253;
 wire net8254;
 wire net8255;
 wire net8257;
 wire net8258;
 wire net8259;
 wire net826;
 wire net8260;
 wire net8261;
 wire net8262;
 wire net8263;
 wire net8264;
 wire net8265;
 wire net8266;
 wire net8267;
 wire net8268;
 wire net8269;
 wire net827;
 wire net8270;
 wire net8272;
 wire net8273;
 wire net8274;
 wire net8275;
 wire net8276;
 wire net828;
 wire net829;
 wire net8296;
 wire net8297;
 wire net8298;
 wire net83;
 wire net830;
 wire net8301;
 wire net8302;
 wire net8303;
 wire net8306;
 wire net8307;
 wire net8308;
 wire net8309;
 wire net831;
 wire net8310;
 wire net8311;
 wire net8312;
 wire net8313;
 wire net8314;
 wire net8315;
 wire net8316;
 wire net8317;
 wire net8318;
 wire net8319;
 wire net832;
 wire net8320;
 wire net8321;
 wire net8322;
 wire net8323;
 wire net8324;
 wire net8325;
 wire net8326;
 wire net8327;
 wire net8328;
 wire net8329;
 wire net833;
 wire net8330;
 wire net8331;
 wire net8332;
 wire net8333;
 wire net8334;
 wire net8335;
 wire net8336;
 wire net8337;
 wire net8338;
 wire net8339;
 wire net834;
 wire net8340;
 wire net8341;
 wire net8342;
 wire net8343;
 wire net8344;
 wire net8345;
 wire net8346;
 wire net8347;
 wire net8348;
 wire net8349;
 wire net835;
 wire net8350;
 wire net8351;
 wire net8352;
 wire net8353;
 wire net8354;
 wire net8355;
 wire net8356;
 wire net8357;
 wire net8358;
 wire net8359;
 wire net836;
 wire net8361;
 wire net8362;
 wire net8364;
 wire net8365;
 wire net8366;
 wire net8367;
 wire net8369;
 wire net837;
 wire net8370;
 wire net8372;
 wire net8373;
 wire net8374;
 wire net8375;
 wire net8377;
 wire net8378;
 wire net8379;
 wire net838;
 wire net8380;
 wire net8381;
 wire net8382;
 wire net8383;
 wire net839;
 wire net8390;
 wire net8391;
 wire net8393;
 wire net8394;
 wire net8395;
 wire net8397;
 wire net8399;
 wire net84;
 wire net840;
 wire net8400;
 wire net8402;
 wire net8403;
 wire net8404;
 wire net8405;
 wire net8409;
 wire net841;
 wire net8410;
 wire net8411;
 wire net8412;
 wire net8413;
 wire net8414;
 wire net8415;
 wire net8416;
 wire net8418;
 wire net842;
 wire net8420;
 wire net8422;
 wire net8423;
 wire net8425;
 wire net843;
 wire net8434;
 wire net8436;
 wire net844;
 wire net8441;
 wire net8442;
 wire net8443;
 wire net8444;
 wire net8446;
 wire net8447;
 wire net845;
 wire net8457;
 wire net846;
 wire net8467;
 wire net847;
 wire net848;
 wire net849;
 wire net8491;
 wire net8497;
 wire net8498;
 wire net85;
 wire net850;
 wire net8500;
 wire net8501;
 wire net851;
 wire net8519;
 wire net852;
 wire net8520;
 wire net853;
 wire net8535;
 wire net854;
 wire net8541;
 wire net8542;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdx[5] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_mapdy[5] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.side_hot ;
 wire \rbzero.spi_registers.got_new_floor ;
 wire \rbzero.spi_registers.got_new_leak ;
 wire \rbzero.spi_registers.got_new_mapd ;
 wire \rbzero.spi_registers.got_new_other ;
 wire \rbzero.spi_registers.got_new_sky ;
 wire \rbzero.spi_registers.got_new_texadd[0] ;
 wire \rbzero.spi_registers.got_new_texadd[1] ;
 wire \rbzero.spi_registers.got_new_texadd[2] ;
 wire \rbzero.spi_registers.got_new_texadd[3] ;
 wire \rbzero.spi_registers.got_new_vinf ;
 wire \rbzero.spi_registers.got_new_vshift ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.new_floor[0] ;
 wire \rbzero.spi_registers.new_floor[1] ;
 wire \rbzero.spi_registers.new_floor[2] ;
 wire \rbzero.spi_registers.new_floor[3] ;
 wire \rbzero.spi_registers.new_floor[4] ;
 wire \rbzero.spi_registers.new_floor[5] ;
 wire \rbzero.spi_registers.new_leak[0] ;
 wire \rbzero.spi_registers.new_leak[1] ;
 wire \rbzero.spi_registers.new_leak[2] ;
 wire \rbzero.spi_registers.new_leak[3] ;
 wire \rbzero.spi_registers.new_leak[4] ;
 wire \rbzero.spi_registers.new_leak[5] ;
 wire \rbzero.spi_registers.new_mapd[0] ;
 wire \rbzero.spi_registers.new_mapd[10] ;
 wire \rbzero.spi_registers.new_mapd[11] ;
 wire \rbzero.spi_registers.new_mapd[12] ;
 wire \rbzero.spi_registers.new_mapd[13] ;
 wire \rbzero.spi_registers.new_mapd[14] ;
 wire \rbzero.spi_registers.new_mapd[15] ;
 wire \rbzero.spi_registers.new_mapd[1] ;
 wire \rbzero.spi_registers.new_mapd[2] ;
 wire \rbzero.spi_registers.new_mapd[3] ;
 wire \rbzero.spi_registers.new_mapd[4] ;
 wire \rbzero.spi_registers.new_mapd[5] ;
 wire \rbzero.spi_registers.new_mapd[6] ;
 wire \rbzero.spi_registers.new_mapd[7] ;
 wire \rbzero.spi_registers.new_mapd[8] ;
 wire \rbzero.spi_registers.new_mapd[9] ;
 wire \rbzero.spi_registers.new_other[0] ;
 wire \rbzero.spi_registers.new_other[10] ;
 wire \rbzero.spi_registers.new_other[1] ;
 wire \rbzero.spi_registers.new_other[2] ;
 wire \rbzero.spi_registers.new_other[3] ;
 wire \rbzero.spi_registers.new_other[4] ;
 wire \rbzero.spi_registers.new_other[6] ;
 wire \rbzero.spi_registers.new_other[7] ;
 wire \rbzero.spi_registers.new_other[8] ;
 wire \rbzero.spi_registers.new_other[9] ;
 wire \rbzero.spi_registers.new_sky[0] ;
 wire \rbzero.spi_registers.new_sky[1] ;
 wire \rbzero.spi_registers.new_sky[2] ;
 wire \rbzero.spi_registers.new_sky[3] ;
 wire \rbzero.spi_registers.new_sky[4] ;
 wire \rbzero.spi_registers.new_sky[5] ;
 wire \rbzero.spi_registers.new_texadd[0][0] ;
 wire \rbzero.spi_registers.new_texadd[0][10] ;
 wire \rbzero.spi_registers.new_texadd[0][11] ;
 wire \rbzero.spi_registers.new_texadd[0][12] ;
 wire \rbzero.spi_registers.new_texadd[0][13] ;
 wire \rbzero.spi_registers.new_texadd[0][14] ;
 wire \rbzero.spi_registers.new_texadd[0][15] ;
 wire \rbzero.spi_registers.new_texadd[0][16] ;
 wire \rbzero.spi_registers.new_texadd[0][17] ;
 wire \rbzero.spi_registers.new_texadd[0][18] ;
 wire \rbzero.spi_registers.new_texadd[0][19] ;
 wire \rbzero.spi_registers.new_texadd[0][1] ;
 wire \rbzero.spi_registers.new_texadd[0][20] ;
 wire \rbzero.spi_registers.new_texadd[0][21] ;
 wire \rbzero.spi_registers.new_texadd[0][22] ;
 wire \rbzero.spi_registers.new_texadd[0][23] ;
 wire \rbzero.spi_registers.new_texadd[0][2] ;
 wire \rbzero.spi_registers.new_texadd[0][3] ;
 wire \rbzero.spi_registers.new_texadd[0][4] ;
 wire \rbzero.spi_registers.new_texadd[0][5] ;
 wire \rbzero.spi_registers.new_texadd[0][6] ;
 wire \rbzero.spi_registers.new_texadd[0][7] ;
 wire \rbzero.spi_registers.new_texadd[0][8] ;
 wire \rbzero.spi_registers.new_texadd[0][9] ;
 wire \rbzero.spi_registers.new_texadd[1][0] ;
 wire \rbzero.spi_registers.new_texadd[1][10] ;
 wire \rbzero.spi_registers.new_texadd[1][11] ;
 wire \rbzero.spi_registers.new_texadd[1][12] ;
 wire \rbzero.spi_registers.new_texadd[1][13] ;
 wire \rbzero.spi_registers.new_texadd[1][14] ;
 wire \rbzero.spi_registers.new_texadd[1][15] ;
 wire \rbzero.spi_registers.new_texadd[1][16] ;
 wire \rbzero.spi_registers.new_texadd[1][17] ;
 wire \rbzero.spi_registers.new_texadd[1][18] ;
 wire \rbzero.spi_registers.new_texadd[1][19] ;
 wire \rbzero.spi_registers.new_texadd[1][1] ;
 wire \rbzero.spi_registers.new_texadd[1][20] ;
 wire \rbzero.spi_registers.new_texadd[1][21] ;
 wire \rbzero.spi_registers.new_texadd[1][22] ;
 wire \rbzero.spi_registers.new_texadd[1][23] ;
 wire \rbzero.spi_registers.new_texadd[1][2] ;
 wire \rbzero.spi_registers.new_texadd[1][3] ;
 wire \rbzero.spi_registers.new_texadd[1][4] ;
 wire \rbzero.spi_registers.new_texadd[1][5] ;
 wire \rbzero.spi_registers.new_texadd[1][6] ;
 wire \rbzero.spi_registers.new_texadd[1][7] ;
 wire \rbzero.spi_registers.new_texadd[1][8] ;
 wire \rbzero.spi_registers.new_texadd[1][9] ;
 wire \rbzero.spi_registers.new_texadd[2][0] ;
 wire \rbzero.spi_registers.new_texadd[2][10] ;
 wire \rbzero.spi_registers.new_texadd[2][11] ;
 wire \rbzero.spi_registers.new_texadd[2][12] ;
 wire \rbzero.spi_registers.new_texadd[2][13] ;
 wire \rbzero.spi_registers.new_texadd[2][14] ;
 wire \rbzero.spi_registers.new_texadd[2][15] ;
 wire \rbzero.spi_registers.new_texadd[2][16] ;
 wire \rbzero.spi_registers.new_texadd[2][17] ;
 wire \rbzero.spi_registers.new_texadd[2][18] ;
 wire \rbzero.spi_registers.new_texadd[2][19] ;
 wire \rbzero.spi_registers.new_texadd[2][1] ;
 wire \rbzero.spi_registers.new_texadd[2][20] ;
 wire \rbzero.spi_registers.new_texadd[2][21] ;
 wire \rbzero.spi_registers.new_texadd[2][22] ;
 wire \rbzero.spi_registers.new_texadd[2][23] ;
 wire \rbzero.spi_registers.new_texadd[2][2] ;
 wire \rbzero.spi_registers.new_texadd[2][3] ;
 wire \rbzero.spi_registers.new_texadd[2][4] ;
 wire \rbzero.spi_registers.new_texadd[2][5] ;
 wire \rbzero.spi_registers.new_texadd[2][6] ;
 wire \rbzero.spi_registers.new_texadd[2][7] ;
 wire \rbzero.spi_registers.new_texadd[2][8] ;
 wire \rbzero.spi_registers.new_texadd[2][9] ;
 wire \rbzero.spi_registers.new_texadd[3][0] ;
 wire \rbzero.spi_registers.new_texadd[3][10] ;
 wire \rbzero.spi_registers.new_texadd[3][11] ;
 wire \rbzero.spi_registers.new_texadd[3][12] ;
 wire \rbzero.spi_registers.new_texadd[3][13] ;
 wire \rbzero.spi_registers.new_texadd[3][14] ;
 wire \rbzero.spi_registers.new_texadd[3][15] ;
 wire \rbzero.spi_registers.new_texadd[3][16] ;
 wire \rbzero.spi_registers.new_texadd[3][17] ;
 wire \rbzero.spi_registers.new_texadd[3][18] ;
 wire \rbzero.spi_registers.new_texadd[3][19] ;
 wire \rbzero.spi_registers.new_texadd[3][1] ;
 wire \rbzero.spi_registers.new_texadd[3][20] ;
 wire \rbzero.spi_registers.new_texadd[3][21] ;
 wire \rbzero.spi_registers.new_texadd[3][22] ;
 wire \rbzero.spi_registers.new_texadd[3][23] ;
 wire \rbzero.spi_registers.new_texadd[3][2] ;
 wire \rbzero.spi_registers.new_texadd[3][3] ;
 wire \rbzero.spi_registers.new_texadd[3][4] ;
 wire \rbzero.spi_registers.new_texadd[3][5] ;
 wire \rbzero.spi_registers.new_texadd[3][6] ;
 wire \rbzero.spi_registers.new_texadd[3][7] ;
 wire \rbzero.spi_registers.new_texadd[3][8] ;
 wire \rbzero.spi_registers.new_texadd[3][9] ;
 wire \rbzero.spi_registers.new_vinf ;
 wire \rbzero.spi_registers.new_vshift[0] ;
 wire \rbzero.spi_registers.new_vshift[1] ;
 wire \rbzero.spi_registers.new_vshift[2] ;
 wire \rbzero.spi_registers.new_vshift[3] ;
 wire \rbzero.spi_registers.new_vshift[4] ;
 wire \rbzero.spi_registers.new_vshift[5] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[16] ;
 wire \rbzero.spi_registers.spi_buffer[17] ;
 wire \rbzero.spi_registers.spi_buffer[18] ;
 wire \rbzero.spi_registers.spi_buffer[19] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[20] ;
 wire \rbzero.spi_registers.spi_buffer[21] ;
 wire \rbzero.spi_registers.spi_buffer[22] ;
 wire \rbzero.spi_registers.spi_buffer[23] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.texadd0[0] ;
 wire \rbzero.spi_registers.texadd0[10] ;
 wire \rbzero.spi_registers.texadd0[11] ;
 wire \rbzero.spi_registers.texadd0[12] ;
 wire \rbzero.spi_registers.texadd0[13] ;
 wire \rbzero.spi_registers.texadd0[14] ;
 wire \rbzero.spi_registers.texadd0[15] ;
 wire \rbzero.spi_registers.texadd0[16] ;
 wire \rbzero.spi_registers.texadd0[17] ;
 wire \rbzero.spi_registers.texadd0[18] ;
 wire \rbzero.spi_registers.texadd0[19] ;
 wire \rbzero.spi_registers.texadd0[1] ;
 wire \rbzero.spi_registers.texadd0[20] ;
 wire \rbzero.spi_registers.texadd0[21] ;
 wire \rbzero.spi_registers.texadd0[22] ;
 wire \rbzero.spi_registers.texadd0[23] ;
 wire \rbzero.spi_registers.texadd0[2] ;
 wire \rbzero.spi_registers.texadd0[3] ;
 wire \rbzero.spi_registers.texadd0[4] ;
 wire \rbzero.spi_registers.texadd0[5] ;
 wire \rbzero.spi_registers.texadd0[6] ;
 wire \rbzero.spi_registers.texadd0[7] ;
 wire \rbzero.spi_registers.texadd0[8] ;
 wire \rbzero.spi_registers.texadd0[9] ;
 wire \rbzero.spi_registers.texadd1[0] ;
 wire \rbzero.spi_registers.texadd1[10] ;
 wire \rbzero.spi_registers.texadd1[11] ;
 wire \rbzero.spi_registers.texadd1[12] ;
 wire \rbzero.spi_registers.texadd1[13] ;
 wire \rbzero.spi_registers.texadd1[14] ;
 wire \rbzero.spi_registers.texadd1[15] ;
 wire \rbzero.spi_registers.texadd1[16] ;
 wire \rbzero.spi_registers.texadd1[17] ;
 wire \rbzero.spi_registers.texadd1[18] ;
 wire \rbzero.spi_registers.texadd1[19] ;
 wire \rbzero.spi_registers.texadd1[1] ;
 wire \rbzero.spi_registers.texadd1[20] ;
 wire \rbzero.spi_registers.texadd1[21] ;
 wire \rbzero.spi_registers.texadd1[22] ;
 wire \rbzero.spi_registers.texadd1[23] ;
 wire \rbzero.spi_registers.texadd1[2] ;
 wire \rbzero.spi_registers.texadd1[3] ;
 wire \rbzero.spi_registers.texadd1[4] ;
 wire \rbzero.spi_registers.texadd1[5] ;
 wire \rbzero.spi_registers.texadd1[6] ;
 wire \rbzero.spi_registers.texadd1[7] ;
 wire \rbzero.spi_registers.texadd1[8] ;
 wire \rbzero.spi_registers.texadd1[9] ;
 wire \rbzero.spi_registers.texadd2[0] ;
 wire \rbzero.spi_registers.texadd2[10] ;
 wire \rbzero.spi_registers.texadd2[11] ;
 wire \rbzero.spi_registers.texadd2[12] ;
 wire \rbzero.spi_registers.texadd2[13] ;
 wire \rbzero.spi_registers.texadd2[14] ;
 wire \rbzero.spi_registers.texadd2[15] ;
 wire \rbzero.spi_registers.texadd2[16] ;
 wire \rbzero.spi_registers.texadd2[17] ;
 wire \rbzero.spi_registers.texadd2[18] ;
 wire \rbzero.spi_registers.texadd2[19] ;
 wire \rbzero.spi_registers.texadd2[1] ;
 wire \rbzero.spi_registers.texadd2[20] ;
 wire \rbzero.spi_registers.texadd2[21] ;
 wire \rbzero.spi_registers.texadd2[22] ;
 wire \rbzero.spi_registers.texadd2[23] ;
 wire \rbzero.spi_registers.texadd2[2] ;
 wire \rbzero.spi_registers.texadd2[3] ;
 wire \rbzero.spi_registers.texadd2[4] ;
 wire \rbzero.spi_registers.texadd2[5] ;
 wire \rbzero.spi_registers.texadd2[6] ;
 wire \rbzero.spi_registers.texadd2[7] ;
 wire \rbzero.spi_registers.texadd2[8] ;
 wire \rbzero.spi_registers.texadd2[9] ;
 wire \rbzero.spi_registers.texadd3[0] ;
 wire \rbzero.spi_registers.texadd3[10] ;
 wire \rbzero.spi_registers.texadd3[11] ;
 wire \rbzero.spi_registers.texadd3[12] ;
 wire \rbzero.spi_registers.texadd3[13] ;
 wire \rbzero.spi_registers.texadd3[14] ;
 wire \rbzero.spi_registers.texadd3[15] ;
 wire \rbzero.spi_registers.texadd3[16] ;
 wire \rbzero.spi_registers.texadd3[17] ;
 wire \rbzero.spi_registers.texadd3[18] ;
 wire \rbzero.spi_registers.texadd3[19] ;
 wire \rbzero.spi_registers.texadd3[1] ;
 wire \rbzero.spi_registers.texadd3[20] ;
 wire \rbzero.spi_registers.texadd3[21] ;
 wire \rbzero.spi_registers.texadd3[22] ;
 wire \rbzero.spi_registers.texadd3[23] ;
 wire \rbzero.spi_registers.texadd3[2] ;
 wire \rbzero.spi_registers.texadd3[3] ;
 wire \rbzero.spi_registers.texadd3[4] ;
 wire \rbzero.spi_registers.texadd3[5] ;
 wire \rbzero.spi_registers.texadd3[6] ;
 wire \rbzero.spi_registers.texadd3[7] ;
 wire \rbzero.spi_registers.texadd3[8] ;
 wire \rbzero.spi_registers.texadd3[9] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.texu_hot[0] ;
 wire \rbzero.texu_hot[1] ;
 wire \rbzero.texu_hot[2] ;
 wire \rbzero.texu_hot[3] ;
 wire \rbzero.texu_hot[4] ;
 wire \rbzero.texu_hot[5] ;
 wire \rbzero.trace_state[0] ;
 wire \rbzero.trace_state[1] ;
 wire \rbzero.trace_state[2] ;
 wire \rbzero.trace_state[3] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_hot[0] ;
 wire \rbzero.wall_hot[1] ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \reg_gpout[0] ;
 wire \reg_gpout[1] ;
 wire \reg_gpout[2] ;
 wire \reg_gpout[3] ;
 wire \reg_gpout[4] ;
 wire \reg_gpout[5] ;
 wire reg_hsync;
 wire \reg_rgb[14] ;
 wire \reg_rgb[15] ;
 wire \reg_rgb[22] ;
 wire \reg_rgb[23] ;
 wire \reg_rgb[6] ;
 wire \reg_rgb[7] ;
 wire reg_vsync;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_04597_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net4705));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_06057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_07903_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_07903_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_08295_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_09094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_04612_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net3469));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net3592));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net4173));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net4490));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_05055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net4490));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net4694));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net4751));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net6143));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net6714));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net8002));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net8467));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_03202_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_04829_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_05680_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_08038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net2094));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net2094));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_05795_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net4293));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net4912));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net8002));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net8012));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net8264));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net8270));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net49));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1067 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_993 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_8 _10439_ (.A(net6038),
    .X(_04020_));
 sky130_fd_sc_hd__clkbuf_8 _10440_ (.A(net6039),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_4 _10441_ (.A(net7710),
    .X(_04022_));
 sky130_fd_sc_hd__buf_4 _10442_ (.A(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__clkbuf_1 _10443_ (.A(net4132),
    .X(_04024_));
 sky130_fd_sc_hd__clkbuf_1 _10444_ (.A(net4145),
    .X(_04025_));
 sky130_fd_sc_hd__and2b_1 _10445_ (.A_N(net4133),
    .B(net4089),
    .X(_04026_));
 sky130_fd_sc_hd__and2_1 _10446_ (.A(_04023_),
    .B(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__xor2_4 _10447_ (.A(net47),
    .B(net48),
    .X(_04028_));
 sky130_fd_sc_hd__and3_2 _10448_ (.A(_04021_),
    .B(_04027_),
    .C(net92),
    .X(_04029_));
 sky130_fd_sc_hd__buf_4 _10449_ (.A(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__clkbuf_4 _10450_ (.A(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__mux2_1 _10451_ (.A0(net3067),
    .A1(net49),
    .S(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__clkbuf_1 _10452_ (.A(net2394),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(net7121),
    .A1(net3067),
    .S(_04031_),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_1 _10454_ (.A(net3068),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _10455_ (.A0(net6940),
    .A1(net7121),
    .S(_04031_),
    .X(_04034_));
 sky130_fd_sc_hd__clkbuf_1 _10456_ (.A(net2549),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(net6581),
    .A1(net6940),
    .S(_04031_),
    .X(_04035_));
 sky130_fd_sc_hd__clkbuf_1 _10458_ (.A(net2027),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(net2348),
    .A1(net6581),
    .S(_04031_),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_1 _10460_ (.A(net6583),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(net6888),
    .A1(net6902),
    .S(_04031_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _10462_ (.A(net2349),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(net6836),
    .A1(net6888),
    .S(_04031_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _10464_ (.A(net2298),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(net2851),
    .A1(net6836),
    .S(_04031_),
    .X(_04039_));
 sky130_fd_sc_hd__clkbuf_1 _10466_ (.A(net6838),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(net6689),
    .A1(net7236),
    .S(_04031_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_1 _10468_ (.A(net2852),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(net2131),
    .A1(net6689),
    .S(_04031_),
    .X(_04041_));
 sky130_fd_sc_hd__clkbuf_1 _10470_ (.A(net6691),
    .X(_01588_));
 sky130_fd_sc_hd__clkbuf_4 _10471_ (.A(_04030_),
    .X(_04042_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(net2780),
    .A1(net6758),
    .S(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_1 _10473_ (.A(net6760),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _10474_ (.A0(net7123),
    .A1(net7365),
    .S(_04042_),
    .X(_04044_));
 sky130_fd_sc_hd__clkbuf_1 _10475_ (.A(net2781),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(net6952),
    .A1(net7123),
    .S(_04042_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _10477_ (.A(net2689),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _10478_ (.A0(net6140),
    .A1(net6952),
    .S(_04042_),
    .X(_04046_));
 sky130_fd_sc_hd__clkbuf_1 _10479_ (.A(net2497),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(net2438),
    .A1(net6140),
    .S(_04042_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_1 _10481_ (.A(net6142),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _10482_ (.A0(net3128),
    .A1(net7328),
    .S(_04042_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_1 _10483_ (.A(net7330),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(net7268),
    .A1(net7359),
    .S(_04042_),
    .X(_04049_));
 sky130_fd_sc_hd__clkbuf_1 _10485_ (.A(net3129),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _10486_ (.A0(net6880),
    .A1(net7268),
    .S(_04042_),
    .X(_04050_));
 sky130_fd_sc_hd__clkbuf_1 _10487_ (.A(net2985),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(net2229),
    .A1(net6880),
    .S(_04042_),
    .X(_04051_));
 sky130_fd_sc_hd__clkbuf_1 _10489_ (.A(net6882),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(net2499),
    .A1(net6975),
    .S(_04042_),
    .X(_04052_));
 sky130_fd_sc_hd__clkbuf_1 _10491_ (.A(net6977),
    .X(_01578_));
 sky130_fd_sc_hd__clkbuf_4 _10492_ (.A(_04030_),
    .X(_04053_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(net7161),
    .A1(net7165),
    .S(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_1 _10494_ (.A(net2500),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(net2657),
    .A1(net7161),
    .S(_04053_),
    .X(_04055_));
 sky130_fd_sc_hd__clkbuf_1 _10496_ (.A(net7163),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(net7063),
    .A1(net2657),
    .S(_04053_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_1 _10498_ (.A(net7065),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _10499_ (.A0(net5788),
    .A1(net7063),
    .S(_04053_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_1 _10500_ (.A(net2260),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(net3240),
    .A1(net5788),
    .S(_04053_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(net5790),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _10503_ (.A0(net5677),
    .A1(net3240),
    .S(_04053_),
    .X(_04059_));
 sky130_fd_sc_hd__clkbuf_1 _10504_ (.A(net5679),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(net2790),
    .A1(net5598),
    .S(_04053_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _10506_ (.A(net5600),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(net6999),
    .A1(net2790),
    .S(_04053_),
    .X(_04061_));
 sky130_fd_sc_hd__clkbuf_1 _10508_ (.A(net2791),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(net6259),
    .A1(net6999),
    .S(_04053_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_1 _10510_ (.A(net2561),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(net2774),
    .A1(net6259),
    .S(_04053_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _10512_ (.A(net6261),
    .X(_01568_));
 sky130_fd_sc_hd__clkbuf_4 _10513_ (.A(_04030_),
    .X(_04064_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(net5645),
    .A1(net7295),
    .S(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__clkbuf_1 _10515_ (.A(net2775),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(net5637),
    .A1(net5645),
    .S(_04064_),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _10517_ (.A(net5647),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(net2373),
    .A1(net5637),
    .S(_04064_),
    .X(_04067_));
 sky130_fd_sc_hd__clkbuf_1 _10519_ (.A(net5639),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _10520_ (.A0(net2797),
    .A1(net7457),
    .S(_04064_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_1 _10521_ (.A(net2798),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(net5696),
    .A1(net2797),
    .S(_04064_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _10523_ (.A(net976),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _10524_ (.A0(net5547),
    .A1(net5696),
    .S(_04064_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_1 _10525_ (.A(net5698),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(net2152),
    .A1(net5547),
    .S(_04064_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _10527_ (.A(net5549),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(net7087),
    .A1(net7439),
    .S(_04064_),
    .X(_04072_));
 sky130_fd_sc_hd__clkbuf_1 _10529_ (.A(net2982),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(net2719),
    .A1(net7087),
    .S(_04064_),
    .X(_04073_));
 sky130_fd_sc_hd__clkbuf_1 _10531_ (.A(net1939),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(net7192),
    .A1(net2719),
    .S(_04064_),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _10533_ (.A(net2720),
    .X(_01558_));
 sky130_fd_sc_hd__clkbuf_4 _10534_ (.A(_04030_),
    .X(_04075_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(net6985),
    .A1(net7192),
    .S(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__clkbuf_1 _10536_ (.A(net2466),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(net6754),
    .A1(net6985),
    .S(_04075_),
    .X(_04077_));
 sky130_fd_sc_hd__clkbuf_1 _10538_ (.A(net2174),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(net6752),
    .A1(net6754),
    .S(_04075_),
    .X(_04078_));
 sky130_fd_sc_hd__clkbuf_1 _10540_ (.A(net1992),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(net6088),
    .A1(net6752),
    .S(_04075_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _10542_ (.A(net1913),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(net1839),
    .A1(net6088),
    .S(_04075_),
    .X(_04080_));
 sky130_fd_sc_hd__clkbuf_1 _10544_ (.A(net6090),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _10545_ (.A0(net2641),
    .A1(net6715),
    .S(_04075_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_1 _10546_ (.A(net6717),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _10547_ (.A0(net6872),
    .A1(net7055),
    .S(_04075_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _10548_ (.A(net2642),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _10549_ (.A0(net5730),
    .A1(net6872),
    .S(_04075_),
    .X(_04083_));
 sky130_fd_sc_hd__clkbuf_1 _10550_ (.A(net2021),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(net5659),
    .A1(net5730),
    .S(_04075_),
    .X(_04084_));
 sky130_fd_sc_hd__clkbuf_1 _10552_ (.A(net5732),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(net2342),
    .A1(net5659),
    .S(_04075_),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _10554_ (.A(net5661),
    .X(_01548_));
 sky130_fd_sc_hd__clkbuf_4 _10555_ (.A(_04030_),
    .X(_04086_));
 sky130_fd_sc_hd__mux2_1 _10556_ (.A0(net2880),
    .A1(net7226),
    .S(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__clkbuf_1 _10557_ (.A(net2768),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(net6922),
    .A1(net2880),
    .S(_04086_),
    .X(_04088_));
 sky130_fd_sc_hd__clkbuf_1 _10559_ (.A(net2881),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(net6195),
    .A1(net6922),
    .S(_04086_),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_1 _10561_ (.A(net2272),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(net6144),
    .A1(net6195),
    .S(_04086_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_1 _10563_ (.A(net1116),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(net2370),
    .A1(net6144),
    .S(_04086_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _10565_ (.A(net6146),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(net7266),
    .A1(net7324),
    .S(_04086_),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _10567_ (.A(net2371),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(net6607),
    .A1(net7266),
    .S(_04086_),
    .X(_04093_));
 sky130_fd_sc_hd__clkbuf_1 _10569_ (.A(net2525),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(net2336),
    .A1(net6607),
    .S(_04086_),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _10571_ (.A(net6609),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(net2324),
    .A1(net6898),
    .S(_04086_),
    .X(_04095_));
 sky130_fd_sc_hd__clkbuf_1 _10573_ (.A(net6900),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(net6554),
    .A1(net6967),
    .S(_04086_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _10575_ (.A(net2325),
    .X(_01538_));
 sky130_fd_sc_hd__clkbuf_4 _10576_ (.A(_04030_),
    .X(_04097_));
 sky130_fd_sc_hd__mux2_1 _10577_ (.A0(net1958),
    .A1(net6554),
    .S(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _10578_ (.A(net6556),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(net1529),
    .A1(net6928),
    .S(_04097_),
    .X(_04099_));
 sky130_fd_sc_hd__clkbuf_1 _10580_ (.A(net6930),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(net5550),
    .A1(net1529),
    .S(_04097_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _10582_ (.A(net5552),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(net5558),
    .A1(net5550),
    .S(_04097_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_1 _10584_ (.A(net5560),
    .X(_01534_));
 sky130_fd_sc_hd__inv_6 _10585_ (.A(_04028_),
    .Y(_04102_));
 sky130_fd_sc_hd__or3b_4 _10586_ (.A(_04102_),
    .B(_04021_),
    .C_N(_04027_),
    .X(_04103_));
 sky130_fd_sc_hd__buf_4 _10587_ (.A(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_4 _10588_ (.A(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(net49),
    .A1(net2947),
    .S(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _10590_ (.A(net2948),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10591_ (.A0(net2947),
    .A1(net7287),
    .S(_04105_),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _10592_ (.A(net2304),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10593_ (.A0(net7287),
    .A1(net2914),
    .S(_04105_),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_1 _10594_ (.A(net7289),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10595_ (.A0(net7415),
    .A1(net7103),
    .S(_04105_),
    .X(_04109_));
 sky130_fd_sc_hd__clkbuf_1 _10596_ (.A(net2915),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(net7103),
    .A1(net6983),
    .S(_04105_),
    .X(_04110_));
 sky130_fd_sc_hd__clkbuf_1 _10598_ (.A(net1843),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(net6983),
    .A1(net6906),
    .S(_04105_),
    .X(_04111_));
 sky130_fd_sc_hd__clkbuf_1 _10600_ (.A(net2531),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(net6906),
    .A1(net2201),
    .S(_04105_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(net6908),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(net7135),
    .A1(net7067),
    .S(_04105_),
    .X(_04113_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(net2202),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(net7067),
    .A1(net2384),
    .S(_04105_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(net7069),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(net7141),
    .A1(net6187),
    .S(_04105_),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(net2385),
    .X(_01524_));
 sky130_fd_sc_hd__clkbuf_4 _10609_ (.A(_04104_),
    .X(_04116_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(net6187),
    .A1(net2247),
    .S(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _10611_ (.A(net6189),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(net7009),
    .A1(net2959),
    .S(_04116_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _10613_ (.A(net7011),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10614_ (.A0(net7403),
    .A1(net7200),
    .S(_04116_),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _10615_ (.A(net2960),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(net7200),
    .A1(net7184),
    .S(_04116_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _10617_ (.A(net2445),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(net7184),
    .A1(net5706),
    .S(_04116_),
    .X(_04121_));
 sky130_fd_sc_hd__clkbuf_1 _10619_ (.A(net2677),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(net5706),
    .A1(net5577),
    .S(_04116_),
    .X(_04122_));
 sky130_fd_sc_hd__buf_1 _10621_ (.A(net5708),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(net5577),
    .A1(net2581),
    .S(_04116_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(net5579),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(net7369),
    .A1(net2610),
    .S(_04116_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(net7371),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(net7469),
    .A1(net2817),
    .S(_04116_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(net2818),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(net2817),
    .A1(net6172),
    .S(_04116_),
    .X(_04126_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(net1895),
    .X(_01514_));
 sky130_fd_sc_hd__clkbuf_4 _10630_ (.A(_04104_),
    .X(_04127_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(net6172),
    .A1(net2993),
    .S(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _10632_ (.A(net6174),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _10633_ (.A0(net7441),
    .A1(net6669),
    .S(_04127_),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_1 _10634_ (.A(net2994),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(net6669),
    .A1(net2423),
    .S(_04127_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _10636_ (.A(net6671),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(net6914),
    .A1(net2043),
    .S(_04127_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _10638_ (.A(net6916),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _10639_ (.A0(net7019),
    .A1(net6822),
    .S(_04127_),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _10640_ (.A(net2044),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(net6822),
    .A1(net1517),
    .S(_04127_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _10642_ (.A(net6824),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(net6826),
    .A1(net2950),
    .S(_04127_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(net6828),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(net7326),
    .A1(net7238),
    .S(_04127_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(net2951),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(net7238),
    .A1(net6735),
    .S(_04127_),
    .X(_04136_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(net2756),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(net6735),
    .A1(net2094),
    .S(_04127_),
    .X(_04137_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(net6737),
    .X(_01504_));
 sky130_fd_sc_hd__clkbuf_4 _10651_ (.A(_04104_),
    .X(_04138_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(net7017),
    .A1(net6651),
    .S(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _10653_ (.A(net2095),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(net6651),
    .A1(net2405),
    .S(_04138_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_1 _10655_ (.A(net6653),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(net6918),
    .A1(net2155),
    .S(_04138_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _10657_ (.A(net6920),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(net7299),
    .A1(net7224),
    .S(_04138_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _10659_ (.A(net2156),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(net7224),
    .A1(net6277),
    .S(_04138_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _10661_ (.A(net2391),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(net6277),
    .A1(net2140),
    .S(_04138_),
    .X(_04144_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(net6279),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(net6860),
    .A1(net6840),
    .S(_04138_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(net2141),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(net6840),
    .A1(net2625),
    .S(_04138_),
    .X(_04146_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(net6842),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(net7222),
    .A1(net6703),
    .S(_04138_),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(net2626),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(net6703),
    .A1(net6084),
    .S(_04138_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(net2092),
    .X(_01494_));
 sky130_fd_sc_hd__clkbuf_4 _10672_ (.A(_04104_),
    .X(_04149_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(net6084),
    .A1(net2294),
    .S(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _10674_ (.A(net6086),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(net7149),
    .A1(net2635),
    .S(_04149_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _10676_ (.A(net7151),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10677_ (.A0(net7220),
    .A1(net7129),
    .S(_04149_),
    .X(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _10678_ (.A(net2636),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(net7129),
    .A1(net6989),
    .S(_04149_),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_1 _10680_ (.A(net2033),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(net6989),
    .A1(net6488),
    .S(_04149_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _10682_ (.A(net2620),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10683_ (.A0(net6488),
    .A1(net2450),
    .S(_04149_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _10684_ (.A(net6490),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(net7208),
    .A1(net6979),
    .S(_04149_),
    .X(_04156_));
 sky130_fd_sc_hd__clkbuf_1 _10686_ (.A(net2451),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(net6979),
    .A1(net2728),
    .S(_04149_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _10688_ (.A(net6981),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(net7348),
    .A1(net7095),
    .S(_04149_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _10690_ (.A(net2729),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(net7095),
    .A1(net6152),
    .S(_04149_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _10692_ (.A(net2188),
    .X(_01484_));
 sky130_fd_sc_hd__clkbuf_4 _10693_ (.A(_04104_),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(net6152),
    .A1(net3356),
    .S(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(net6154),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(net7518),
    .A1(net6834),
    .S(_04160_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10697_ (.A(net3357),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(net6834),
    .A1(net5688),
    .S(_04160_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _10699_ (.A(net1927),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(net5688),
    .A1(net5544),
    .S(_04160_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _10701_ (.A(net5690),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(net5544),
    .A1(net2122),
    .S(_04160_),
    .X(_04165_));
 sky130_fd_sc_hd__clkbuf_1 _10703_ (.A(net5546),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(net6963),
    .A1(net2143),
    .S(_04160_),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_1 _10705_ (.A(net6965),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(net7285),
    .A1(net2661),
    .S(_04160_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(net2662),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(net2661),
    .A1(net7035),
    .S(_04160_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(net2319),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(net7035),
    .A1(net2592),
    .S(_04160_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(net7037),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(net7252),
    .A1(net5991),
    .S(_04160_),
    .X(_04170_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(net2593),
    .X(_01474_));
 sky130_fd_sc_hd__clkbuf_4 _10714_ (.A(_04104_),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(net5991),
    .A1(net5630),
    .S(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _10716_ (.A(net591),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(net5630),
    .A1(net5601),
    .S(_04171_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _10718_ (.A(net5632),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(net5601),
    .A1(net2793),
    .S(_04171_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _10720_ (.A(net5603),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(net2793),
    .A1(net6359),
    .S(_04171_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _10722_ (.A(net6361),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(net2907),
    .A1(net50),
    .S(_04097_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _10724_ (.A(net2908),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(net7117),
    .A1(net2907),
    .S(_04097_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(net2811),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(net6818),
    .A1(net7117),
    .S(_04097_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(net2748),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10729_ (.A0(net2049),
    .A1(net6818),
    .S(_04097_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(net6820),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10731_ (.A0(net6796),
    .A1(net2049),
    .S(_04097_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _10732_ (.A(net6798),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(net6227),
    .A1(net6796),
    .S(_04097_),
    .X(_04181_));
 sky130_fd_sc_hd__clkbuf_1 _10734_ (.A(net1995),
    .X(_01464_));
 sky130_fd_sc_hd__clkbuf_4 _10735_ (.A(_04030_),
    .X(_04182_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(net2244),
    .A1(net6227),
    .S(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(net6229),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(net6910),
    .A1(net2244),
    .S(_04182_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(net6912),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(net6615),
    .A1(net6910),
    .S(_04182_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_1 _10741_ (.A(net2701),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(net2417),
    .A1(net6615),
    .S(_04182_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _10743_ (.A(net6617),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(net2999),
    .A1(net7029),
    .S(_04182_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _10745_ (.A(net7031),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(net7262),
    .A1(net7427),
    .S(_04182_),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _10747_ (.A(net3000),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(net2518),
    .A1(net7262),
    .S(_04182_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _10749_ (.A(net7264),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(net6466),
    .A1(net7275),
    .S(_04182_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _10751_ (.A(net2519),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(net2008),
    .A1(net6466),
    .S(_04182_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(net6468),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(net6203),
    .A1(net6772),
    .S(_04182_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _10755_ (.A(net2009),
    .X(_01454_));
 sky130_fd_sc_hd__buf_4 _10756_ (.A(_04029_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_4 _10757_ (.A(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(net2288),
    .A1(net6203),
    .S(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(net6205),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(net6243),
    .A1(net7015),
    .S(_04194_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(net2289),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(net2750),
    .A1(net6243),
    .S(_04194_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(net6245),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(net2376),
    .A1(net7079),
    .S(_04194_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(net7081),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(net7137),
    .A1(net2376),
    .S(_04194_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(net7139),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(net7091),
    .A1(net7137),
    .S(_04194_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(net2552),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(net6812),
    .A1(net7091),
    .S(_04194_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _10771_ (.A(net2433),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(net2533),
    .A1(net6812),
    .S(_04194_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _10773_ (.A(net6814),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(net7105),
    .A1(net7381),
    .S(_04194_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _10775_ (.A(net2534),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(net6114),
    .A1(net7105),
    .S(_04194_),
    .X(_04204_));
 sky130_fd_sc_hd__clkbuf_1 _10777_ (.A(net2177),
    .X(_01444_));
 sky130_fd_sc_hd__clkbuf_4 _10778_ (.A(_04193_),
    .X(_04205_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(net2429),
    .A1(net6114),
    .S(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(net6116),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(net2569),
    .A1(net6719),
    .S(_04205_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(net6721),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(net2471),
    .A1(net7180),
    .S(_04205_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(net7182),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(net7210),
    .A1(net7399),
    .S(_04205_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(net2472),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(net6456),
    .A1(net7210),
    .S(_04205_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(net2460),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(net2408),
    .A1(net6456),
    .S(_04205_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(net6458),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(net6991),
    .A1(net2408),
    .S(_04205_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(net6993),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(net7001),
    .A1(net6991),
    .S(_04205_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _10794_ (.A(net2567),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(net7373),
    .A1(net7001),
    .S(_04205_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(net2971),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(net6168),
    .A1(net7373),
    .S(_04205_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _10798_ (.A(net3170),
    .X(_01434_));
 sky130_fd_sc_hd__clkbuf_4 _10799_ (.A(_04193_),
    .X(_04216_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(net1985),
    .A1(net6168),
    .S(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _10801_ (.A(net6170),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(net2515),
    .A1(net6784),
    .S(_04216_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(net6786),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(net6643),
    .A1(net7153),
    .S(_04216_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(net2516),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(net2996),
    .A1(net6643),
    .S(_04216_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(net6645),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(net7250),
    .A1(net7429),
    .S(_04216_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _10809_ (.A(net2997),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(net7171),
    .A1(net7250),
    .S(_04216_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(net2652),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(net2521),
    .A1(net7171),
    .S(_04216_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(net7173),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(net6808),
    .A1(net7336),
    .S(_04216_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _10815_ (.A(net2522),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(net2638),
    .A1(net6808),
    .S(_04216_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(net6810),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(net6478),
    .A1(net7293),
    .S(_04216_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _10819_ (.A(net2639),
    .X(_01424_));
 sky130_fd_sc_hd__clkbuf_4 _10820_ (.A(_04193_),
    .X(_04227_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(net2783),
    .A1(net6478),
    .S(_04227_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(net6480),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(net6774),
    .A1(net7340),
    .S(_04227_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(net2784),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(net6750),
    .A1(net6774),
    .S(_04227_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(net2086),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(net6211),
    .A1(net6750),
    .S(_04227_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _10828_ (.A(net2030),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(net3249),
    .A1(net6211),
    .S(_04227_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(net6213),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(net7492),
    .A1(net7514),
    .S(_04227_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(net3250),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(net2848),
    .A1(net7492),
    .S(_04227_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(net7494),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(net7005),
    .A1(net2848),
    .S(_04227_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(net7007),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(net7043),
    .A1(net7005),
    .S(_04227_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(net2739),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(net6034),
    .A1(net7043),
    .S(_04227_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(net2966),
    .X(_01414_));
 sky130_fd_sc_hd__clkbuf_4 _10841_ (.A(_04193_),
    .X(_04238_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(net2023),
    .A1(net6034),
    .S(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _10843_ (.A(net6036),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(net7049),
    .A1(net7111),
    .S(_04238_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _10845_ (.A(net2024),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10846_ (.A0(net6223),
    .A1(net7049),
    .S(_04238_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _10847_ (.A(net2400),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10848_ (.A0(net2595),
    .A1(net6223),
    .S(_04238_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _10849_ (.A(net6225),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10850_ (.A0(net7351),
    .A1(net2595),
    .S(_04238_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _10851_ (.A(net7353),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(net5662),
    .A1(net2462),
    .S(_04238_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _10853_ (.A(net5664),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(net3104),
    .A1(net5700),
    .S(_04238_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _10855_ (.A(net5702),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10856_ (.A0(net6293),
    .A1(net3104),
    .S(_04238_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _10857_ (.A(net6295),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10858_ (.A0(net50),
    .A1(net2503),
    .S(_04171_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _10859_ (.A(net2504),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10860_ (.A0(net2503),
    .A1(net6587),
    .S(_04171_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _10861_ (.A(net2477),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(net6587),
    .A1(net2826),
    .S(_04171_),
    .X(_04249_));
 sky130_fd_sc_hd__buf_1 _10863_ (.A(net6589),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(net7431),
    .A1(net7145),
    .S(_04171_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _10865_ (.A(net2827),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(net7145),
    .A1(net7131),
    .S(_04171_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(net2292),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(net7131),
    .A1(net2685),
    .S(_04171_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(net7133),
    .X(_01400_));
 sky130_fd_sc_hd__clkbuf_4 _10870_ (.A(_04104_),
    .X(_04253_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(net7216),
    .A1(net6593),
    .S(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _10872_ (.A(net2686),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _10873_ (.A0(net6593),
    .A1(net2886),
    .S(_04253_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _10874_ (.A(net6595),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(net2886),
    .A1(net7355),
    .S(_04253_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _10876_ (.A(net7357),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(net7355),
    .A1(net7186),
    .S(_04253_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _10878_ (.A(net2924),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(net7186),
    .A1(net6756),
    .S(_04253_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _10880_ (.A(net2692),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(net6756),
    .A1(net6092),
    .S(_04253_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _10882_ (.A(net2053),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(net6092),
    .A1(net2575),
    .S(_04253_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _10884_ (.A(net6094),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(net7291),
    .A1(net6884),
    .S(_04253_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(net2576),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(net6884),
    .A1(net1964),
    .S(_04253_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(net6886),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(net7051),
    .A1(net2900),
    .S(_04253_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(net7053),
    .X(_01390_));
 sky130_fd_sc_hd__clkbuf_4 _10891_ (.A(_04103_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_4 _10892_ (.A(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(net7477),
    .A1(net3202),
    .S(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(net7479),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(net7500),
    .A1(net6924),
    .S(_04265_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(net3203),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(net6924),
    .A1(net2589),
    .S(_04265_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(net6926),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(net7279),
    .A1(net7057),
    .S(_04265_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(net2590),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(net7057),
    .A1(net7033),
    .S(_04265_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(net2236),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(net7033),
    .A1(net6164),
    .S(_04265_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(net2454),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(net6164),
    .A1(net2282),
    .S(_04265_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(net6166),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(net7167),
    .A1(net3070),
    .S(_04265_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(net7169),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(net7397),
    .A1(net6762),
    .S(_04265_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(net3071),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(net6762),
    .A1(net6235),
    .S(_04265_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(net1901),
    .X(_01380_));
 sky130_fd_sc_hd__clkbuf_4 _10913_ (.A(_04264_),
    .X(_04276_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(net6235),
    .A1(net2604),
    .S(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _10915_ (.A(net6237),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(net7423),
    .A1(net6854),
    .S(_04276_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _10917_ (.A(net2605),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(net6854),
    .A1(net3176),
    .S(_04276_),
    .X(_04279_));
 sky130_fd_sc_hd__buf_1 _10919_ (.A(net6856),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(net7437),
    .A1(net7234),
    .S(_04276_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _10921_ (.A(net3177),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(net7234),
    .A1(net7190),
    .S(_04276_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(net2732),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(net7190),
    .A1(net6072),
    .S(_04276_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(net2617),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(net6072),
    .A1(net3107),
    .S(_04276_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(net6074),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(net7486),
    .A1(net3246),
    .S(_04276_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(net7488),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(net7532),
    .A1(net7433),
    .S(_04276_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _10931_ (.A(net3247),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(net7433),
    .A1(net3263),
    .S(_04276_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _10933_ (.A(net7435),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_4 _10934_ (.A(_04264_),
    .X(_04287_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(net7484),
    .A1(net7232),
    .S(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _10936_ (.A(net3264),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(net7232),
    .A1(net6723),
    .S(_04287_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _10938_ (.A(net2723),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _10939_ (.A0(net6723),
    .A1(net2217),
    .S(_04287_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _10940_ (.A(net6725),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(net7071),
    .A1(net2300),
    .S(_04287_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _10942_ (.A(net7073),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(net7316),
    .A1(net2482),
    .S(_04287_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(net7318),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(net7361),
    .A1(net6107),
    .S(_04287_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(net2483),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(net6107),
    .A1(net2110),
    .S(_04287_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(net6109),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(net6711),
    .A1(net2265),
    .S(_04287_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(net6713),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(net6936),
    .A1(net6591),
    .S(_04287_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _10952_ (.A(net2266),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _10953_ (.A0(net6591),
    .A1(net6506),
    .S(_04287_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _10954_ (.A(net1740),
    .X(_01360_));
 sky130_fd_sc_hd__clkbuf_4 _10955_ (.A(_04264_),
    .X(_04298_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(net6506),
    .A1(net1920),
    .S(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _10957_ (.A(net6508),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(net6776),
    .A1(net2017),
    .S(_04298_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _10959_ (.A(net6778),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(net7228),
    .A1(net3029),
    .S(_04298_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _10961_ (.A(net7230),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(net7473),
    .A1(net7194),
    .S(_04298_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _10963_ (.A(net3030),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(net7194),
    .A1(net6705),
    .S(_04298_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _10965_ (.A(net2492),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(net6705),
    .A1(net6197),
    .S(_04298_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _10967_ (.A(net1873),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(net6197),
    .A1(net1715),
    .S(_04298_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(net6199),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(net6641),
    .A1(net6500),
    .S(_04298_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(net1716),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(net6500),
    .A1(net2670),
    .S(_04298_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(net6502),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(net7254),
    .A1(net2715),
    .S(_04298_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _10975_ (.A(net7256),
    .X(_01350_));
 sky130_fd_sc_hd__buf_4 _10976_ (.A(_04264_),
    .X(_04309_));
 sky130_fd_sc_hd__mux2_1 _10977_ (.A0(net7314),
    .A1(net7013),
    .S(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _10978_ (.A(net2716),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(net7013),
    .A1(net6655),
    .S(_04309_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _10980_ (.A(net2355),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(net6655),
    .A1(net6633),
    .S(_04309_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _10982_ (.A(net1974),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10983_ (.A0(net6633),
    .A1(net2116),
    .S(_04309_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _10984_ (.A(net6635),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(net6874),
    .A1(net2857),
    .S(_04309_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _10986_ (.A(net6876),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(net2857),
    .A1(net7212),
    .S(_04309_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _10988_ (.A(net7214),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(net655),
    .A1(net5640),
    .S(_04309_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _10990_ (.A(net5642),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(net5640),
    .A1(net5714),
    .S(_04309_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _10992_ (.A(net5716),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(net2845),
    .A1(net51),
    .S(_04238_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _10994_ (.A(net2846),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(net6345),
    .A1(net2845),
    .S(_04238_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _10996_ (.A(net2683),
    .X(_01340_));
 sky130_fd_sc_hd__clkbuf_4 _10997_ (.A(_04193_),
    .X(_04320_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(net5653),
    .A1(net6345),
    .S(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_1 _10999_ (.A(net1299),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(net5574),
    .A1(net5653),
    .S(_04320_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _11001_ (.A(net5655),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(net2285),
    .A1(net5574),
    .S(_04320_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _11003_ (.A(net5576),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _11004_ (.A0(net3163),
    .A1(net7389),
    .S(_04320_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _11005_ (.A(net2867),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _11006_ (.A0(net7101),
    .A1(net3163),
    .S(_04320_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _11007_ (.A(net3164),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _11008_ (.A0(net6548),
    .A1(net7101),
    .S(_04320_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _11009_ (.A(net2114),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _11010_ (.A0(net2253),
    .A1(net6548),
    .S(_04320_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _11011_ (.A(net6550),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(net7157),
    .A1(net7240),
    .S(_04320_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _11013_ (.A(net2254),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(net2545),
    .A1(net7157),
    .S(_04320_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _11015_ (.A(net7159),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(net6249),
    .A1(net7338),
    .S(_04320_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _11017_ (.A(net2546),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_4 _11018_ (.A(_04193_),
    .X(_04331_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(net2063),
    .A1(net6249),
    .S(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_1 _11020_ (.A(net6251),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(net2667),
    .A1(net6894),
    .S(_04331_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _11022_ (.A(net6896),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(net5718),
    .A1(net7451),
    .S(_04331_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _11024_ (.A(net2668),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _11025_ (.A0(net5669),
    .A1(net5718),
    .S(_04331_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _11026_ (.A(net5720),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(net2735),
    .A1(net5669),
    .S(_04331_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _11028_ (.A(net5671),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(net6118),
    .A1(net2735),
    .S(_04331_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _11030_ (.A(net2736),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(net2000),
    .A1(net6118),
    .S(_04331_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _11032_ (.A(net6120),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(net6442),
    .A1(net6764),
    .S(_04331_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _11034_ (.A(net2001),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(net2937),
    .A1(net6442),
    .S(_04331_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _11036_ (.A(net6444),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(net7196),
    .A1(net7344),
    .S(_04331_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _11038_ (.A(net2938),
    .X(_01320_));
 sky130_fd_sc_hd__clkbuf_4 _11039_ (.A(_04193_),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(net2777),
    .A1(net7196),
    .S(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _11041_ (.A(net7198),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _11042_ (.A0(net7039),
    .A1(net7218),
    .S(_04342_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _11043_ (.A(net2778),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _11044_ (.A0(net2333),
    .A1(net7039),
    .S(_04342_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _11045_ (.A(net7041),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _11046_ (.A0(net7346),
    .A1(net7401),
    .S(_04342_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _11047_ (.A(net2334),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _11048_ (.A0(net7099),
    .A1(net7346),
    .S(_04342_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _11049_ (.A(net2707),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _11050_ (.A0(net6219),
    .A1(net7099),
    .S(_04342_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _11051_ (.A(net2358),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(net1408),
    .A1(net6219),
    .S(_04342_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _11053_ (.A(net6221),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(net1955),
    .A1(net6524),
    .S(_04342_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(net6526),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(net5634),
    .A1(net6766),
    .S(_04342_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _11057_ (.A(net1956),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(net5589),
    .A1(net5634),
    .S(_04342_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _11059_ (.A(net5636),
    .X(_01310_));
 sky130_fd_sc_hd__clkbuf_4 _11060_ (.A(_04193_),
    .X(_04353_));
 sky130_fd_sc_hd__mux2_1 _11061_ (.A0(net2632),
    .A1(net5589),
    .S(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _11062_ (.A(net5591),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _11063_ (.A0(net6866),
    .A1(net2632),
    .S(_04353_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _11064_ (.A(net2633),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _11065_ (.A0(net5649),
    .A1(net6866),
    .S(_04353_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _11066_ (.A(net1889),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _11067_ (.A0(net5592),
    .A1(net5649),
    .S(_04353_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _11068_ (.A(net5651),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _11069_ (.A0(net2239),
    .A1(net5592),
    .S(_04353_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _11070_ (.A(net5594),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _11071_ (.A0(net6128),
    .A1(net2239),
    .S(_04353_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _11072_ (.A(net2240),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(net1797),
    .A1(net6128),
    .S(_04353_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _11074_ (.A(net6130),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(net1660),
    .A1(net6657),
    .S(_04353_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _11076_ (.A(net6659),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(net2274),
    .A1(net6699),
    .S(_04353_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _11078_ (.A(net6701),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(net3092),
    .A1(net6948),
    .S(_04353_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _11080_ (.A(net6950),
    .X(_01300_));
 sky130_fd_sc_hd__clkbuf_4 _11081_ (.A(_04193_),
    .X(_04364_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(net6846),
    .A1(net7322),
    .S(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _11083_ (.A(net3093),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(net3243),
    .A1(net6846),
    .S(_04364_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _11085_ (.A(net6848),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(net7306),
    .A1(net7530),
    .S(_04364_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _11087_ (.A(net3244),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(net2557),
    .A1(net7306),
    .S(_04364_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _11089_ (.A(net7308),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(net2367),
    .A1(net7383),
    .S(_04364_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _11091_ (.A(net7385),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(net6184),
    .A1(net7407),
    .S(_04364_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_1 _11093_ (.A(net2368),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(net5673),
    .A1(net6184),
    .S(_04364_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(net1070),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(net5586),
    .A1(net5673),
    .S(_04364_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(net5675),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(net2978),
    .A1(net5586),
    .S(_04364_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(net5588),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(net6271),
    .A1(net2978),
    .S(_04364_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(net2979),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_4 _11102_ (.A(_04029_),
    .X(_04375_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(net2664),
    .A1(net6271),
    .S(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _11104_ (.A(net6273),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _11105_ (.A0(net2601),
    .A1(net7075),
    .S(_04375_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _11106_ (.A(net7077),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _11107_ (.A0(net6637),
    .A1(net7097),
    .S(_04375_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _11108_ (.A(net2602),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(net2578),
    .A1(net6637),
    .S(_04375_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _11110_ (.A(net6639),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(net6890),
    .A1(net2578),
    .S(_04375_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _11112_ (.A(net6892),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(net6052),
    .A1(net6890),
    .S(_04375_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _11114_ (.A(net2537),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(net2149),
    .A1(net6052),
    .S(_04375_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(net6054),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(net2930),
    .A1(net6956),
    .S(_04375_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(net6958),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(net5684),
    .A1(net7342),
    .S(_04375_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _11120_ (.A(net2931),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(net5680),
    .A1(net5684),
    .S(_04375_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _11122_ (.A(net5686),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _11123_ (.A0(net2351),
    .A1(net5680),
    .S(_04030_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _11124_ (.A(net5682),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(net6267),
    .A1(net2351),
    .S(_04030_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _11126_ (.A(net6269),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(net51),
    .A1(net6904),
    .S(_04309_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _11128_ (.A(net1968),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(net6904),
    .A1(net6946),
    .S(_04309_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(net2083),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_4 _11131_ (.A(_04264_),
    .X(_04390_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(net6946),
    .A1(net2648),
    .S(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _11133_ (.A(net2361),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(net2648),
    .A1(net6026),
    .S(_04390_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _11135_ (.A(net2649),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(net6026),
    .A1(net2279),
    .S(_04390_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _11137_ (.A(net6028),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _11138_ (.A0(net6973),
    .A1(net6746),
    .S(_04390_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _11139_ (.A(net2280),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _11140_ (.A0(net6746),
    .A1(net1819),
    .S(_04390_),
    .X(_04395_));
 sky130_fd_sc_hd__clkbuf_1 _11141_ (.A(net6748),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(net6804),
    .A1(net2512),
    .S(_04390_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(net6806),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _11144_ (.A0(net7242),
    .A1(net6534),
    .S(_04390_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _11145_ (.A(net2513),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(net6534),
    .A1(net2987),
    .S(_04390_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _11147_ (.A(net6536),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(net7405),
    .A1(net6995),
    .S(_04390_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _11149_ (.A(net2988),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(net6995),
    .A1(net2387),
    .S(_04390_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _11151_ (.A(net6997),
    .X(_01074_));
 sky130_fd_sc_hd__clkbuf_4 _11152_ (.A(_04264_),
    .X(_04401_));
 sky130_fd_sc_hd__mux2_1 _11153_ (.A0(net7204),
    .A1(net2539),
    .S(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _11154_ (.A(net7206),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _11155_ (.A0(net7363),
    .A1(net6103),
    .S(_04401_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _11156_ (.A(net2540),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _11157_ (.A0(net6103),
    .A1(net2572),
    .S(_04401_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _11158_ (.A(net6105),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(net7244),
    .A1(net2488),
    .S(_04401_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _11160_ (.A(net7246),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(net7377),
    .A1(net3117),
    .S(_04401_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _11162_ (.A(net7379),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(net7504),
    .A1(net6460),
    .S(_04401_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(net3118),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(net6460),
    .A1(net1982),
    .S(_04401_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _11166_ (.A(net6462),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(net6788),
    .A1(net2804),
    .S(_04401_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _11168_ (.A(net6790),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(net7447),
    .A1(net7417),
    .S(_04401_),
    .X(_04410_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(net2805),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(net7417),
    .A1(net7393),
    .S(_04401_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(net2655),
    .X(_01064_));
 sky130_fd_sc_hd__clkbuf_4 _11173_ (.A(_04264_),
    .X(_04412_));
 sky130_fd_sc_hd__mux2_1 _11174_ (.A0(net7393),
    .A1(net7391),
    .S(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _11175_ (.A(net2814),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _11176_ (.A0(net7391),
    .A1(net6156),
    .S(_04412_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _11177_ (.A(net2674),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _11178_ (.A0(net6156),
    .A1(net1929),
    .S(_04412_),
    .X(_04415_));
 sky130_fd_sc_hd__clkbuf_1 _11179_ (.A(net6158),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _11180_ (.A0(net7025),
    .A1(net2381),
    .S(_04412_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _11181_ (.A(net7027),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _11182_ (.A0(net7248),
    .A1(net7059),
    .S(_04412_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _11183_ (.A(net2382),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(net7059),
    .A1(net2841),
    .S(_04412_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(net7061),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(net7147),
    .A1(net7089),
    .S(_04412_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _11187_ (.A(net2842),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(net7089),
    .A1(net6538),
    .S(_04412_),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(net2726),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(net6538),
    .A1(net1773),
    .S(_04412_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_1 _11191_ (.A(net6540),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(net6942),
    .A1(net2744),
    .S(_04412_),
    .X(_04422_));
 sky130_fd_sc_hd__clkbuf_1 _11193_ (.A(net6944),
    .X(_01054_));
 sky130_fd_sc_hd__clkbuf_4 _11194_ (.A(_04264_),
    .X(_04423_));
 sky130_fd_sc_hd__mux2_1 _11195_ (.A0(net7270),
    .A1(net6987),
    .S(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _11196_ (.A(net2745),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _11197_ (.A0(net6987),
    .A1(net6096),
    .S(_04423_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _11198_ (.A(net2457),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _11199_ (.A0(net6096),
    .A1(net1897),
    .S(_04423_),
    .X(_04426_));
 sky130_fd_sc_hd__clkbuf_1 _11200_ (.A(net6098),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _11201_ (.A0(net6830),
    .A1(net2527),
    .S(_04423_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _11202_ (.A(net6832),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(net7107),
    .A1(net2962),
    .S(_04423_),
    .X(_04428_));
 sky130_fd_sc_hd__clkbuf_1 _11204_ (.A(net7109),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(net7459),
    .A1(net7202),
    .S(_04423_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _11206_ (.A(net2963),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(net7202),
    .A1(net6673),
    .S(_04423_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(net2608),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(net6673),
    .A1(net1758),
    .S(_04423_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(net6675),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(net6850),
    .A1(net2854),
    .S(_04423_),
    .X(_04432_));
 sky130_fd_sc_hd__clkbuf_1 _11212_ (.A(net6852),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(net7301),
    .A1(net7297),
    .S(_04423_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _11214_ (.A(net2855),
    .X(_01044_));
 sky130_fd_sc_hd__clkbuf_4 _11215_ (.A(_04264_),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_1 _11216_ (.A0(net7297),
    .A1(net6802),
    .S(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _11217_ (.A(net2480),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _11218_ (.A0(net6802),
    .A1(net6030),
    .S(_04434_),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_1 _11219_ (.A(net1825),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _11220_ (.A0(net6030),
    .A1(net2679),
    .S(_04434_),
    .X(_04437_));
 sky130_fd_sc_hd__clkbuf_1 _11221_ (.A(net6032),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _11222_ (.A0(net7125),
    .A1(net2917),
    .S(_04434_),
    .X(_04438_));
 sky130_fd_sc_hd__clkbuf_1 _11223_ (.A(net7127),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _11224_ (.A0(net7387),
    .A1(net6768),
    .S(_04434_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _11225_ (.A(net2918),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(net6768),
    .A1(net2345),
    .S(_04434_),
    .X(_04440_));
 sky130_fd_sc_hd__clkbuf_1 _11227_ (.A(net6770),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(net7332),
    .A1(net6780),
    .S(_04434_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _11229_ (.A(net2346),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _11230_ (.A0(net6780),
    .A1(net2170),
    .S(_04434_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _11231_ (.A(net6782),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(net7119),
    .A1(net6868),
    .S(_04434_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _11233_ (.A(net2171),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(net6868),
    .A1(net2911),
    .S(_04434_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_1 _11235_ (.A(net6870),
    .X(_01034_));
 sky130_fd_sc_hd__clkbuf_4 _11236_ (.A(_04103_),
    .X(_04445_));
 sky130_fd_sc_hd__mux2_1 _11237_ (.A0(net7281),
    .A1(net2892),
    .S(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _11238_ (.A(net7283),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _11239_ (.A0(net7320),
    .A1(net6215),
    .S(_04445_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _11240_ (.A(net2893),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(net6215),
    .A1(net2072),
    .S(_04445_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _11242_ (.A(net6217),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _11243_ (.A0(net6932),
    .A1(net2832),
    .S(_04445_),
    .X(_04449_));
 sky130_fd_sc_hd__clkbuf_1 _11244_ (.A(net6934),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _11245_ (.A0(net7258),
    .A1(net3005),
    .S(_04445_),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _11246_ (.A(net7260),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _11247_ (.A0(net7413),
    .A1(net7023),
    .S(_04445_),
    .X(_04451_));
 sky130_fd_sc_hd__clkbuf_1 _11248_ (.A(net3006),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(net7023),
    .A1(net6969),
    .S(_04445_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _11250_ (.A(net2316),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(net6969),
    .A1(net2164),
    .S(_04445_),
    .X(_04453_));
 sky130_fd_sc_hd__clkbuf_1 _11252_ (.A(net6971),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _11253_ (.A0(net7113),
    .A1(net2895),
    .S(_04445_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _11254_ (.A(net7115),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(net7375),
    .A1(net5626),
    .S(_04445_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_1 _11256_ (.A(net2896),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _11257_ (.A0(net5626),
    .A1(net5566),
    .S(_04104_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _11258_ (.A(net5628),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(net5566),
    .A1(net1836),
    .S(_04104_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _11260_ (.A(net5568),
    .X(_01022_));
 sky130_fd_sc_hd__clkbuf_8 _11261_ (.A(_04102_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_8 _11262_ (.A(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__buf_8 _11263_ (.A(_04459_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 _11264_ (.A(net5911),
    .X(_04460_));
 sky130_fd_sc_hd__buf_4 _11265_ (.A(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__clkbuf_4 _11266_ (.A(net5946),
    .X(_04462_));
 sky130_fd_sc_hd__inv_2 _11267_ (.A(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__clkbuf_4 _11268_ (.A(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__clkinv_4 _11269_ (.A(net4057),
    .Y(_04465_));
 sky130_fd_sc_hd__nor2_2 _11270_ (.A(_04464_),
    .B(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__clkbuf_4 _11271_ (.A(net5205),
    .X(_04467_));
 sky130_fd_sc_hd__buf_4 _11272_ (.A(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__o21a_1 _11273_ (.A1(_04461_),
    .A2(_04466_),
    .B1(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__a21bo_1 _11274_ (.A1(_04461_),
    .A2(_04466_),
    .B1_N(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__or4b_1 _11275_ (.A(_04023_),
    .B(_04470_),
    .C(net4133),
    .D_N(net4089),
    .X(_04471_));
 sky130_fd_sc_hd__buf_8 _11276_ (.A(_04471_),
    .X(net71));
 sky130_fd_sc_hd__inv_2 _11277_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .Y(_04472_));
 sky130_fd_sc_hd__clkbuf_1 _11278_ (.A(net5922),
    .X(_04473_));
 sky130_fd_sc_hd__buf_1 _11279_ (.A(net3975),
    .X(_04474_));
 sky130_fd_sc_hd__or2_1 _11280_ (.A(net4083),
    .B(net4862),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_2 _11281_ (.A(net4863),
    .X(_04476_));
 sky130_fd_sc_hd__inv_2 _11282_ (.A(net4186),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_2 _11283_ (.A(net3337),
    .B(net92),
    .Y(_04478_));
 sky130_fd_sc_hd__inv_2 _11284_ (.A(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__clkbuf_4 _11285_ (.A(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__buf_4 _11286_ (.A(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__buf_4 _11287_ (.A(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__o31ai_2 _11288_ (.A1(net3871),
    .A2(net3976),
    .A3(_04476_),
    .B1(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__inv_2 _11289_ (.A(net4083),
    .Y(_04484_));
 sky130_fd_sc_hd__buf_2 _11290_ (.A(net4862),
    .X(_04485_));
 sky130_fd_sc_hd__or4b_2 _11291_ (.A(net3871),
    .B(net3976),
    .C(net3774),
    .D_N(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__or4bb_1 _11292_ (.A(net3976),
    .B(net4083),
    .C_N(_04485_),
    .D_N(net3871),
    .X(_04487_));
 sky130_fd_sc_hd__nand2_1 _11293_ (.A(_04486_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__buf_4 _11294_ (.A(_04478_),
    .X(_04489_));
 sky130_fd_sc_hd__buf_4 _11295_ (.A(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__o32ai_1 _11296_ (.A1(net8051),
    .A2(_04483_),
    .A3(_04488_),
    .B1(_04490_),
    .B2(_04486_),
    .Y(_00001_));
 sky130_fd_sc_hd__o21ai_4 _11297_ (.A1(_04023_),
    .A2(_04469_),
    .B1(_04026_),
    .Y(net70));
 sky130_fd_sc_hd__clkbuf_4 _11298_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _11299_ (.A(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__a31o_1 _11300_ (.A1(net8217),
    .A2(_04486_),
    .A3(_04487_),
    .B1(_04483_),
    .X(_00000_));
 sky130_fd_sc_hd__inv_2 _11301_ (.A(net71),
    .Y(_04493_));
 sky130_fd_sc_hd__buf_6 _11302_ (.A(net7678),
    .X(_04494_));
 sky130_fd_sc_hd__clkbuf_8 _11303_ (.A(net7708),
    .X(_04495_));
 sky130_fd_sc_hd__buf_4 _11304_ (.A(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__or3_1 _11305_ (.A(net3954),
    .B(_04495_),
    .C(net3641),
    .X(_04497_));
 sky130_fd_sc_hd__o21ai_1 _11306_ (.A1(_04494_),
    .A2(_04496_),
    .B1(_04021_),
    .Y(_04498_));
 sky130_fd_sc_hd__a22o_1 _11307_ (.A1(_04494_),
    .A2(_04496_),
    .B1(_04497_),
    .B2(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__buf_4 _11308_ (.A(_04462_),
    .X(_04500_));
 sky130_fd_sc_hd__clkinv_4 _11309_ (.A(net5205),
    .Y(_04501_));
 sky130_fd_sc_hd__inv_2 _11310_ (.A(net3641),
    .Y(_04502_));
 sky130_fd_sc_hd__clkbuf_4 _11311_ (.A(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__buf_4 _11312_ (.A(net7747),
    .X(_04504_));
 sky130_fd_sc_hd__buf_4 _11313_ (.A(net7748),
    .X(_04505_));
 sky130_fd_sc_hd__and2_2 _11314_ (.A(_04504_),
    .B(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__nor3b_1 _11315_ (.A(_04504_),
    .B(_04505_),
    .C_N(\rbzero.spi_registers.texadd3[14] ),
    .Y(_04507_));
 sky130_fd_sc_hd__mux2_1 _11316_ (.A0(\rbzero.spi_registers.texadd3[13] ),
    .A1(\rbzero.spi_registers.texadd1[13] ),
    .S(_04504_),
    .X(_04508_));
 sky130_fd_sc_hd__or2b_1 _11317_ (.A(_04505_),
    .B_N(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__clkbuf_2 _11318_ (.A(net4180),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_8 _11319_ (.A(net4181),
    .X(_04511_));
 sky130_fd_sc_hd__mux4_2 _11320_ (.A0(\rbzero.spi_registers.texadd3[12] ),
    .A1(\rbzero.spi_registers.texadd1[12] ),
    .A2(\rbzero.spi_registers.texadd0[12] ),
    .A3(\rbzero.spi_registers.texadd2[12] ),
    .S0(_04504_),
    .S1(_04505_),
    .X(_04512_));
 sky130_fd_sc_hd__and2_1 _11321_ (.A(_04511_),
    .B(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__mux4_2 _11322_ (.A0(\rbzero.spi_registers.texadd3[11] ),
    .A1(\rbzero.spi_registers.texadd1[11] ),
    .A2(\rbzero.spi_registers.texadd0[11] ),
    .A3(\rbzero.spi_registers.texadd2[11] ),
    .S0(_04504_),
    .S1(_04505_),
    .X(_04514_));
 sky130_fd_sc_hd__nand2_1 _11323_ (.A(\rbzero.texu_hot[5] ),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__mux4_2 _11324_ (.A0(\rbzero.spi_registers.texadd3[10] ),
    .A1(\rbzero.spi_registers.texadd1[10] ),
    .A2(\rbzero.spi_registers.texadd0[10] ),
    .A3(\rbzero.spi_registers.texadd2[10] ),
    .S0(_04504_),
    .S1(_04505_),
    .X(_04516_));
 sky130_fd_sc_hd__nand2_1 _11325_ (.A(\rbzero.texu_hot[4] ),
    .B(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__mux4_2 _11326_ (.A0(\rbzero.spi_registers.texadd3[9] ),
    .A1(\rbzero.spi_registers.texadd1[9] ),
    .A2(\rbzero.spi_registers.texadd0[9] ),
    .A3(\rbzero.spi_registers.texadd2[9] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _11327_ (.A(\rbzero.texu_hot[3] ),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__mux4_2 _11328_ (.A0(\rbzero.spi_registers.texadd3[8] ),
    .A1(\rbzero.spi_registers.texadd1[8] ),
    .A2(\rbzero.spi_registers.texadd0[8] ),
    .A3(\rbzero.spi_registers.texadd2[8] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04520_));
 sky130_fd_sc_hd__nand2_1 _11329_ (.A(\rbzero.texu_hot[2] ),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__mux4_2 _11330_ (.A0(\rbzero.spi_registers.texadd3[7] ),
    .A1(\rbzero.spi_registers.texadd1[7] ),
    .A2(\rbzero.spi_registers.texadd0[7] ),
    .A3(\rbzero.spi_registers.texadd2[7] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04522_));
 sky130_fd_sc_hd__nand2_1 _11331_ (.A(\rbzero.texu_hot[1] ),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__mux4_2 _11332_ (.A0(\rbzero.spi_registers.texadd3[6] ),
    .A1(\rbzero.spi_registers.texadd1[6] ),
    .A2(\rbzero.spi_registers.texadd0[6] ),
    .A3(\rbzero.spi_registers.texadd2[6] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04524_));
 sky130_fd_sc_hd__nand2_1 _11333_ (.A(\rbzero.texu_hot[0] ),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__or2_1 _11334_ (.A(\rbzero.texu_hot[1] ),
    .B(_04522_),
    .X(_04526_));
 sky130_fd_sc_hd__nand2_1 _11335_ (.A(_04523_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__or2_1 _11336_ (.A(_04525_),
    .B(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__or2_1 _11337_ (.A(\rbzero.texu_hot[2] ),
    .B(_04520_),
    .X(_04529_));
 sky130_fd_sc_hd__nand2_1 _11338_ (.A(_04521_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__a21o_1 _11339_ (.A1(_04523_),
    .A2(_04528_),
    .B1(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__or2_1 _11340_ (.A(\rbzero.texu_hot[3] ),
    .B(_04518_),
    .X(_04532_));
 sky130_fd_sc_hd__nand2_1 _11341_ (.A(_04519_),
    .B(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__a21o_1 _11342_ (.A1(_04521_),
    .A2(_04531_),
    .B1(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__or2_1 _11343_ (.A(\rbzero.texu_hot[4] ),
    .B(_04516_),
    .X(_04535_));
 sky130_fd_sc_hd__nand2_1 _11344_ (.A(_04517_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__a21o_1 _11345_ (.A1(_04519_),
    .A2(_04534_),
    .B1(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__or2_1 _11346_ (.A(\rbzero.texu_hot[5] ),
    .B(_04514_),
    .X(_04538_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(_04515_),
    .B(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__a21o_1 _11348_ (.A1(_04517_),
    .A2(_04537_),
    .B1(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__nor2_1 _11349_ (.A(_04511_),
    .B(_04512_),
    .Y(_04541_));
 sky130_fd_sc_hd__or2_1 _11350_ (.A(_04513_),
    .B(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__a21oi_1 _11351_ (.A1(_04515_),
    .A2(_04540_),
    .B1(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__inv_2 _11352_ (.A(_04506_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2b_2 _11353_ (.A_N(_04504_),
    .B(_04505_),
    .Y(_04545_));
 sky130_fd_sc_hd__o221a_1 _11354_ (.A1(\rbzero.spi_registers.texadd2[13] ),
    .A2(_04544_),
    .B1(_04545_),
    .B2(\rbzero.spi_registers.texadd0[13] ),
    .C1(_04509_),
    .X(_04546_));
 sky130_fd_sc_hd__o21ai_1 _11355_ (.A1(_04513_),
    .A2(_04543_),
    .B1(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__and2b_2 _11356_ (.A_N(_04505_),
    .B(_04504_),
    .X(_04548_));
 sky130_fd_sc_hd__inv_2 _11357_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .Y(_04549_));
 sky130_fd_sc_hd__a2bb2o_1 _11358_ (.A1_N(\rbzero.spi_registers.texadd0[14] ),
    .A2_N(_04545_),
    .B1(_04548_),
    .B2(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__a211o_1 _11359_ (.A1(\rbzero.spi_registers.texadd2[14] ),
    .A2(_04506_),
    .B1(_04507_),
    .C1(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__a21oi_1 _11360_ (.A1(_04509_),
    .A2(_04547_),
    .B1(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a211o_1 _11361_ (.A1(\rbzero.spi_registers.texadd2[14] ),
    .A2(_04506_),
    .B1(_04507_),
    .C1(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__buf_4 _11362_ (.A(_04504_),
    .X(_04554_));
 sky130_fd_sc_hd__buf_4 _11363_ (.A(_04505_),
    .X(_04555_));
 sky130_fd_sc_hd__mux4_2 _11364_ (.A0(\rbzero.spi_registers.texadd3[15] ),
    .A1(\rbzero.spi_registers.texadd1[15] ),
    .A2(\rbzero.spi_registers.texadd0[15] ),
    .A3(\rbzero.spi_registers.texadd2[15] ),
    .S0(_04554_),
    .S1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__mux4_2 _11365_ (.A0(\rbzero.spi_registers.texadd3[16] ),
    .A1(\rbzero.spi_registers.texadd1[16] ),
    .A2(\rbzero.spi_registers.texadd0[16] ),
    .A3(\rbzero.spi_registers.texadd2[16] ),
    .S0(_04504_),
    .S1(_04505_),
    .X(_04557_));
 sky130_fd_sc_hd__and3_1 _11366_ (.A(_04553_),
    .B(_04556_),
    .C(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__mux4_2 _11367_ (.A0(\rbzero.spi_registers.texadd3[17] ),
    .A1(\rbzero.spi_registers.texadd1[17] ),
    .A2(\rbzero.spi_registers.texadd0[17] ),
    .A3(\rbzero.spi_registers.texadd2[17] ),
    .S0(_04554_),
    .S1(_04555_),
    .X(_04559_));
 sky130_fd_sc_hd__mux4_2 _11368_ (.A0(\rbzero.spi_registers.texadd3[18] ),
    .A1(\rbzero.spi_registers.texadd1[18] ),
    .A2(\rbzero.spi_registers.texadd0[18] ),
    .A3(\rbzero.spi_registers.texadd2[18] ),
    .S0(_04554_),
    .S1(_04555_),
    .X(_04560_));
 sky130_fd_sc_hd__and3_1 _11369_ (.A(_04558_),
    .B(_04559_),
    .C(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__mux4_2 _11370_ (.A0(\rbzero.spi_registers.texadd3[19] ),
    .A1(\rbzero.spi_registers.texadd1[19] ),
    .A2(\rbzero.spi_registers.texadd0[19] ),
    .A3(\rbzero.spi_registers.texadd2[19] ),
    .S0(_04554_),
    .S1(_04555_),
    .X(_04562_));
 sky130_fd_sc_hd__mux4_1 _11371_ (.A0(\rbzero.spi_registers.texadd3[20] ),
    .A1(\rbzero.spi_registers.texadd1[20] ),
    .A2(\rbzero.spi_registers.texadd0[20] ),
    .A3(\rbzero.spi_registers.texadd2[20] ),
    .S0(_04554_),
    .S1(_04555_),
    .X(_04563_));
 sky130_fd_sc_hd__and3_1 _11372_ (.A(_04561_),
    .B(_04562_),
    .C(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__a21oi_1 _11373_ (.A1(_04561_),
    .A2(_04562_),
    .B1(_04563_),
    .Y(_04565_));
 sky130_fd_sc_hd__buf_4 _11374_ (.A(_04554_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_4 _11375_ (.A(_04555_),
    .X(_04567_));
 sky130_fd_sc_hd__mux4_1 _11376_ (.A0(\rbzero.spi_registers.texadd3[21] ),
    .A1(\rbzero.spi_registers.texadd1[21] ),
    .A2(\rbzero.spi_registers.texadd0[21] ),
    .A3(\rbzero.spi_registers.texadd2[21] ),
    .S0(_04566_),
    .S1(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__nand2_1 _11377_ (.A(_04564_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__or2_1 _11378_ (.A(_04564_),
    .B(_04568_),
    .X(_04570_));
 sky130_fd_sc_hd__nand3_1 _11379_ (.A(_04503_),
    .B(_04569_),
    .C(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__o311a_1 _11380_ (.A1(_04503_),
    .A2(_04564_),
    .A3(_04565_),
    .B1(_04571_),
    .C1(_04496_),
    .X(_04572_));
 sky130_fd_sc_hd__o21ba_1 _11381_ (.A1(\rbzero.spi_registers.texadd3[22] ),
    .A2(_04567_),
    .B1_N(_04554_),
    .X(_04573_));
 sky130_fd_sc_hd__a221o_1 _11382_ (.A1(\rbzero.spi_registers.texadd2[22] ),
    .A2(_04567_),
    .B1(_04548_),
    .B2(\rbzero.spi_registers.texadd1[22] ),
    .C1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__o21ai_1 _11383_ (.A1(\rbzero.spi_registers.texadd0[22] ),
    .A2(_04545_),
    .B1(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__and3_1 _11384_ (.A(_04021_),
    .B(_04569_),
    .C(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__or2_1 _11385_ (.A(_04569_),
    .B(_04575_),
    .X(_04577_));
 sky130_fd_sc_hd__inv_2 _11386_ (.A(\rbzero.spi_registers.texadd0[23] ),
    .Y(_04578_));
 sky130_fd_sc_hd__and2b_1 _11387_ (.A_N(_04566_),
    .B(\rbzero.spi_registers.texadd3[23] ),
    .X(_04579_));
 sky130_fd_sc_hd__a221o_1 _11388_ (.A1(\rbzero.spi_registers.texadd2[23] ),
    .A2(_04506_),
    .B1(_04548_),
    .B2(\rbzero.spi_registers.texadd1[23] ),
    .C1(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__nand2_1 _11389_ (.A(_04545_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__o211a_1 _11390_ (.A1(_04578_),
    .A2(_04545_),
    .B1(_04581_),
    .C1(_04503_),
    .X(_04582_));
 sky130_fd_sc_hd__xnor2_1 _11391_ (.A(_04577_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__clkinv_4 _11392_ (.A(net3857),
    .Y(_04584_));
 sky130_fd_sc_hd__o21a_1 _11393_ (.A1(_04576_),
    .A2(_04583_),
    .B1(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__a21oi_1 _11394_ (.A1(_04558_),
    .A2(_04559_),
    .B1(_04560_),
    .Y(_04586_));
 sky130_fd_sc_hd__nand2_1 _11395_ (.A(_04561_),
    .B(_04562_),
    .Y(_04587_));
 sky130_fd_sc_hd__or2_1 _11396_ (.A(_04561_),
    .B(_04562_),
    .X(_04588_));
 sky130_fd_sc_hd__nand3_1 _11397_ (.A(_04503_),
    .B(_04587_),
    .C(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__o311a_1 _11398_ (.A1(_04503_),
    .A2(_04561_),
    .A3(_04586_),
    .B1(_04589_),
    .C1(_04584_),
    .X(_04590_));
 sky130_fd_sc_hd__and2_1 _11399_ (.A(_04553_),
    .B(_04556_),
    .X(_04591_));
 sky130_fd_sc_hd__nor2_1 _11400_ (.A(_04591_),
    .B(_04557_),
    .Y(_04592_));
 sky130_fd_sc_hd__nor2_1 _11401_ (.A(_04558_),
    .B(_04559_),
    .Y(_04593_));
 sky130_fd_sc_hd__nand2_1 _11402_ (.A(_04558_),
    .B(_04559_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _11403_ (.A(_04503_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__o32a_1 _11404_ (.A1(_04503_),
    .A2(_04558_),
    .A3(_04592_),
    .B1(_04593_),
    .B2(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__inv_2 _11405_ (.A(net3954),
    .Y(_04597_));
 sky130_fd_sc_hd__a21o_1 _11406_ (.A1(_04496_),
    .A2(_04596_),
    .B1(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__o32a_2 _11407_ (.A1(_04494_),
    .A2(_04572_),
    .A3(_04585_),
    .B1(_04590_),
    .B2(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__clkbuf_4 _11408_ (.A(net7562),
    .X(_04600_));
 sky130_fd_sc_hd__nor2_2 _11409_ (.A(_04462_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__o32a_1 _11410_ (.A1(_04500_),
    .A2(_04501_),
    .A3(_04599_),
    .B1(_04601_),
    .B2(_04466_),
    .X(_04602_));
 sky130_fd_sc_hd__nor2_1 _11411_ (.A(net71),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__and3_1 _11412_ (.A(_04509_),
    .B(_04547_),
    .C(_04551_),
    .X(_04604_));
 sky130_fd_sc_hd__and3_1 _11413_ (.A(_04542_),
    .B(_04515_),
    .C(_04540_),
    .X(_04605_));
 sky130_fd_sc_hd__or3_1 _11414_ (.A(_04584_),
    .B(_04543_),
    .C(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__o31a_1 _11415_ (.A1(_04496_),
    .A2(_04552_),
    .A3(_04604_),
    .B1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__or2_1 _11416_ (.A(_04553_),
    .B(_04556_),
    .X(_04608_));
 sky130_fd_sc_hd__or3b_1 _11417_ (.A(_04496_),
    .B(_04591_),
    .C_N(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__or3_1 _11418_ (.A(_04513_),
    .B(_04543_),
    .C(_04546_),
    .X(_04610_));
 sky130_fd_sc_hd__a31oi_1 _11419_ (.A1(_04496_),
    .A2(_04547_),
    .A3(_04610_),
    .B1(_04021_),
    .Y(_04611_));
 sky130_fd_sc_hd__a221o_2 _11420_ (.A1(_04021_),
    .A2(_04607_),
    .B1(_04609_),
    .B2(_04611_),
    .C1(_04494_),
    .X(_04612_));
 sky130_fd_sc_hd__nand3_1 _11421_ (.A(_04536_),
    .B(_04519_),
    .C(_04534_),
    .Y(_04613_));
 sky130_fd_sc_hd__and2_1 _11422_ (.A(_04537_),
    .B(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__nand3_1 _11423_ (.A(_04539_),
    .B(_04517_),
    .C(_04537_),
    .Y(_04615_));
 sky130_fd_sc_hd__and2_1 _11424_ (.A(_04540_),
    .B(_04615_),
    .X(_04616_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(_04614_),
    .A1(_04616_),
    .S(_04503_),
    .X(_04617_));
 sky130_fd_sc_hd__nand3_1 _11426_ (.A(_04521_),
    .B(_04531_),
    .C(_04533_),
    .Y(_04618_));
 sky130_fd_sc_hd__and3_1 _11427_ (.A(_04503_),
    .B(_04534_),
    .C(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__nand3_1 _11428_ (.A(_04530_),
    .B(_04523_),
    .C(_04528_),
    .Y(_04620_));
 sky130_fd_sc_hd__a31o_1 _11429_ (.A1(_04021_),
    .A2(_04531_),
    .A3(_04620_),
    .B1(_04584_),
    .X(_04621_));
 sky130_fd_sc_hd__o221ai_4 _11430_ (.A1(_04496_),
    .A2(_04617_),
    .B1(_04619_),
    .B2(_04621_),
    .C1(_04494_),
    .Y(_04622_));
 sky130_fd_sc_hd__or2_1 _11431_ (.A(\rbzero.texu_hot[0] ),
    .B(_04524_),
    .X(_04623_));
 sky130_fd_sc_hd__and2_1 _11432_ (.A(_04525_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__nand2_1 _11433_ (.A(_04525_),
    .B(_04527_),
    .Y(_04625_));
 sky130_fd_sc_hd__and2_1 _11434_ (.A(_04528_),
    .B(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__mux4_1 _11435_ (.A0(\rbzero.spi_registers.texadd3[4] ),
    .A1(\rbzero.spi_registers.texadd1[4] ),
    .A2(\rbzero.spi_registers.texadd0[4] ),
    .A3(\rbzero.spi_registers.texadd2[4] ),
    .S0(_04566_),
    .S1(_04567_),
    .X(_04627_));
 sky130_fd_sc_hd__mux4_1 _11436_ (.A0(\rbzero.spi_registers.texadd3[5] ),
    .A1(\rbzero.spi_registers.texadd1[5] ),
    .A2(\rbzero.spi_registers.texadd0[5] ),
    .A3(\rbzero.spi_registers.texadd2[5] ),
    .S0(_04566_),
    .S1(_04567_),
    .X(_04628_));
 sky130_fd_sc_hd__mux4_1 _11437_ (.A0(_04624_),
    .A1(_04626_),
    .A2(_04627_),
    .A3(_04628_),
    .S0(_04503_),
    .S1(_04496_),
    .X(_04629_));
 sky130_fd_sc_hd__mux2_1 _11438_ (.A0(\rbzero.spi_registers.texadd0[3] ),
    .A1(\rbzero.spi_registers.texadd0[2] ),
    .S(_04020_),
    .X(_04630_));
 sky130_fd_sc_hd__mux2_1 _11439_ (.A0(\rbzero.spi_registers.texadd0[1] ),
    .A1(\rbzero.spi_registers.texadd0[0] ),
    .S(_04020_),
    .X(_04631_));
 sky130_fd_sc_hd__or3b_1 _11440_ (.A(_04554_),
    .B(_04555_),
    .C_N(\rbzero.spi_registers.texadd3[2] ),
    .X(_04632_));
 sky130_fd_sc_hd__a21bo_1 _11441_ (.A1(\rbzero.spi_registers.texadd2[2] ),
    .A2(_04506_),
    .B1_N(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__and2_1 _11442_ (.A(\rbzero.spi_registers.texadd1[2] ),
    .B(_04548_),
    .X(_04634_));
 sky130_fd_sc_hd__a31o_1 _11443_ (.A1(\rbzero.spi_registers.texadd2[3] ),
    .A2(_04566_),
    .A3(_04567_),
    .B1(_04020_),
    .X(_04635_));
 sky130_fd_sc_hd__or3b_1 _11444_ (.A(_04554_),
    .B(_04555_),
    .C_N(\rbzero.spi_registers.texadd3[3] ),
    .X(_04636_));
 sky130_fd_sc_hd__a21bo_1 _11445_ (.A1(\rbzero.spi_registers.texadd1[3] ),
    .A2(_04548_),
    .B1_N(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__o32a_1 _11446_ (.A1(_04502_),
    .A2(_04633_),
    .A3(_04634_),
    .B1(_04635_),
    .B2(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__and3_1 _11447_ (.A(\rbzero.spi_registers.texadd2[0] ),
    .B(_04566_),
    .C(_04567_),
    .X(_04639_));
 sky130_fd_sc_hd__or3b_1 _11448_ (.A(_04554_),
    .B(_04555_),
    .C_N(\rbzero.spi_registers.texadd3[0] ),
    .X(_04640_));
 sky130_fd_sc_hd__a21bo_1 _11449_ (.A1(\rbzero.spi_registers.texadd1[0] ),
    .A2(_04548_),
    .B1_N(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__a31o_1 _11450_ (.A1(\rbzero.spi_registers.texadd2[1] ),
    .A2(_04566_),
    .A3(_04567_),
    .B1(_04020_),
    .X(_04642_));
 sky130_fd_sc_hd__or3b_1 _11451_ (.A(_04566_),
    .B(_04555_),
    .C_N(\rbzero.spi_registers.texadd3[1] ),
    .X(_04643_));
 sky130_fd_sc_hd__a21bo_1 _11452_ (.A1(\rbzero.spi_registers.texadd1[1] ),
    .A2(_04548_),
    .B1_N(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__o32a_1 _11453_ (.A1(_04502_),
    .A2(_04639_),
    .A3(_04641_),
    .B1(_04642_),
    .B2(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__mux4_1 _11454_ (.A0(_04630_),
    .A1(_04631_),
    .A2(_04638_),
    .A3(_04645_),
    .S0(_04495_),
    .S1(_04545_),
    .X(_04646_));
 sky130_fd_sc_hd__mux2_1 _11455_ (.A0(_04629_),
    .A1(_04646_),
    .S(_04494_),
    .X(_04647_));
 sky130_fd_sc_hd__buf_4 _11456_ (.A(_04600_),
    .X(_04648_));
 sky130_fd_sc_hd__a31o_1 _11457_ (.A1(_04500_),
    .A2(_04461_),
    .A3(_04648_),
    .B1(_04468_),
    .X(_04649_));
 sky130_fd_sc_hd__o21ai_1 _11458_ (.A1(_04500_),
    .A2(_04647_),
    .B1(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__a31oi_1 _11459_ (.A1(_04465_),
    .A2(_04612_),
    .A3(_04622_),
    .B1(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__or3_1 _11460_ (.A(_04466_),
    .B(_04601_),
    .C(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__a32o_4 _11461_ (.A1(_04466_),
    .A2(_04493_),
    .A3(_04499_),
    .B1(_04603_),
    .B2(_04652_),
    .X(net72));
 sky130_fd_sc_hd__inv_2 _11462__1 (.A(clknet_4_9__leaf_i_clk),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _11463_ (.A(net2),
    .Y(_04653_));
 sky130_fd_sc_hd__nand2_1 _11464_ (.A(net3871),
    .B(net3975),
    .Y(_04654_));
 sky130_fd_sc_hd__nand2_1 _11465_ (.A(net4083),
    .B(net4862),
    .Y(_04655_));
 sky130_fd_sc_hd__o21a_1 _11466_ (.A1(net3452),
    .A2(net3628),
    .B1(net2),
    .X(_04656_));
 sky130_fd_sc_hd__inv_2 _11467_ (.A(net4176),
    .Y(_04657_));
 sky130_fd_sc_hd__nor2_2 _11468_ (.A(net4126),
    .B(net4160),
    .Y(_04658_));
 sky130_fd_sc_hd__nand2_2 _11469_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__nor3_2 _11470_ (.A(net4110),
    .B(net4023),
    .C(net4102),
    .Y(_04660_));
 sky130_fd_sc_hd__or2b_1 _11471_ (.A(_04659_),
    .B_N(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__or4b_1 _11472_ (.A(net3995),
    .B(net4065),
    .C(net4091),
    .D_N(net3),
    .X(_04662_));
 sky130_fd_sc_hd__nand2_1 _11473_ (.A(net3857),
    .B(net3641),
    .Y(_04663_));
 sky130_fd_sc_hd__nor2_2 _11474_ (.A(net3955),
    .B(net3858),
    .Y(_04664_));
 sky130_fd_sc_hd__and2_1 _11475_ (.A(net5946),
    .B(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__or2_2 _11476_ (.A(net7562),
    .B(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__o211a_1 _11477_ (.A1(net4105),
    .A2(_04666_),
    .B1(net4115),
    .C1(net3516),
    .X(_04667_));
 sky130_fd_sc_hd__a21oi_1 _11478_ (.A1(net4132),
    .A2(_04667_),
    .B1(net4145),
    .Y(_04668_));
 sky130_fd_sc_hd__a211oi_1 _11479_ (.A1(net4138),
    .A2(_04661_),
    .B1(_04662_),
    .C1(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__buf_2 _11480_ (.A(net4176),
    .X(_04670_));
 sky130_fd_sc_hd__xnor2_1 _11481_ (.A(net4177),
    .B(net4436),
    .Y(_04671_));
 sky130_fd_sc_hd__clkbuf_1 _11482_ (.A(net4160),
    .X(_04672_));
 sky130_fd_sc_hd__xnor2_1 _11483_ (.A(net4095),
    .B(net3326),
    .Y(_04673_));
 sky130_fd_sc_hd__inv_2 _11484_ (.A(net3473),
    .Y(_04674_));
 sky130_fd_sc_hd__xnor2_1 _11485_ (.A(net4126),
    .B(net4748),
    .Y(_04675_));
 sky130_fd_sc_hd__o221a_1 _11486_ (.A1(net4138),
    .A2(_04674_),
    .B1(net3443),
    .B2(_04464_),
    .C1(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__a22o_1 _11487_ (.A1(net3443),
    .A2(_04464_),
    .B1(_04501_),
    .B2(net3431),
    .X(_04677_));
 sky130_fd_sc_hd__inv_2 _11488_ (.A(net3990),
    .Y(_04678_));
 sky130_fd_sc_hd__inv_2 _11489_ (.A(net4091),
    .Y(_04679_));
 sky130_fd_sc_hd__o22a_1 _11490_ (.A1(_04679_),
    .A2(net3552),
    .B1(net3990),
    .B2(_04465_),
    .X(_04680_));
 sky130_fd_sc_hd__o221a_1 _11491_ (.A1(net3431),
    .A2(_04501_),
    .B1(_04600_),
    .B2(net3991),
    .C1(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__inv_2 _11492_ (.A(net4138),
    .Y(_04682_));
 sky130_fd_sc_hd__inv_2 _11493_ (.A(net4105),
    .Y(_04683_));
 sky130_fd_sc_hd__buf_4 _11494_ (.A(net4106),
    .X(_04684_));
 sky130_fd_sc_hd__inv_2 _11495_ (.A(net3552),
    .Y(_04685_));
 sky130_fd_sc_hd__inv_2 _11496_ (.A(net5915),
    .Y(_04686_));
 sky130_fd_sc_hd__o22a_1 _11497_ (.A1(net4091),
    .A2(net3553),
    .B1(_04686_),
    .B2(_04460_),
    .X(_04687_));
 sky130_fd_sc_hd__o221a_1 _11498_ (.A1(_04682_),
    .A2(net3473),
    .B1(net3389),
    .B2(_04684_),
    .C1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__xnor2_1 _11499_ (.A(net3682),
    .B(_04022_),
    .Y(_04689_));
 sky130_fd_sc_hd__and4b_1 _11500_ (.A_N(_04677_),
    .B(_04681_),
    .C(_04688_),
    .D(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__and4_1 _11501_ (.A(_04671_),
    .B(_04673_),
    .C(_04676_),
    .D(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__inv_2 _11502_ (.A(net8207),
    .Y(_04692_));
 sky130_fd_sc_hd__xnor2_1 _11503_ (.A(net5981),
    .B(net3445),
    .Y(_04693_));
 sky130_fd_sc_hd__o221a_1 _11504_ (.A1(net4102),
    .A2(_04692_),
    .B1(net8193),
    .B2(net3955),
    .C1(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__inv_2 _11505_ (.A(net3461),
    .Y(_04695_));
 sky130_fd_sc_hd__xor2_1 _11506_ (.A(net4110),
    .B(net4188),
    .X(_04696_));
 sky130_fd_sc_hd__a221o_1 _11507_ (.A1(net4102),
    .A2(_04692_),
    .B1(_04695_),
    .B2(_04495_),
    .C1(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__xor2_1 _11508_ (.A(net3457),
    .B(net3641),
    .X(_04698_));
 sky130_fd_sc_hd__a221o_1 _11509_ (.A1(net2898),
    .A2(net3955),
    .B1(_04584_),
    .B2(net3461),
    .C1(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__nor2_1 _11510_ (.A(_04697_),
    .B(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__or2_1 _11511_ (.A(_04022_),
    .B(_04467_),
    .X(_04701_));
 sky130_fd_sc_hd__or3b_1 _11512_ (.A(_04701_),
    .B(_04460_),
    .C_N(_04601_),
    .X(_04702_));
 sky130_fd_sc_hd__or2_1 _11513_ (.A(net3642),
    .B(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__or3_1 _11514_ (.A(net4091),
    .B(net4138),
    .C(_04661_),
    .X(_04704_));
 sky130_fd_sc_hd__or3b_1 _11515_ (.A(net6044),
    .B(net4145),
    .C_N(net1),
    .X(_04705_));
 sky130_fd_sc_hd__a221o_2 _11516_ (.A1(net4132),
    .A2(_04703_),
    .B1(_04704_),
    .B2(net5965),
    .C1(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__a31o_1 _11517_ (.A1(_04691_),
    .A2(_04694_),
    .A3(_04700_),
    .B1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__xor2_1 _11518_ (.A(net4095),
    .B(net1817),
    .X(_04708_));
 sky130_fd_sc_hd__or2_1 _11519_ (.A(net4176),
    .B(net4324),
    .X(_04709_));
 sky130_fd_sc_hd__nand2_1 _11520_ (.A(_04670_),
    .B(net4324),
    .Y(_04710_));
 sky130_fd_sc_hd__or2_1 _11521_ (.A(net4126),
    .B(net2038),
    .X(_04711_));
 sky130_fd_sc_hd__buf_1 _11522_ (.A(net4126),
    .X(_04712_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(net4127),
    .B(net2038),
    .Y(_04713_));
 sky130_fd_sc_hd__a2bb2o_1 _11524_ (.A1_N(_04464_),
    .A2_N(net4152),
    .B1(net4306),
    .B2(_04682_),
    .X(_04714_));
 sky130_fd_sc_hd__a221o_1 _11525_ (.A1(_04709_),
    .A2(_04710_),
    .B1(_04711_),
    .B2(_04713_),
    .C1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__xor2_1 _11526_ (.A(net2185),
    .B(_04022_),
    .X(_04716_));
 sky130_fd_sc_hd__a221o_1 _11527_ (.A1(net4152),
    .A2(_04464_),
    .B1(_04501_),
    .B2(net8170),
    .C1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__inv_2 _11528_ (.A(net4309),
    .Y(_04718_));
 sky130_fd_sc_hd__o22a_1 _11529_ (.A1(_04679_),
    .A2(net1803),
    .B1(net4309),
    .B2(_04465_),
    .X(_04719_));
 sky130_fd_sc_hd__o221a_1 _11530_ (.A1(net4347),
    .A2(_04501_),
    .B1(_04600_),
    .B2(_04718_),
    .C1(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__inv_2 _11531_ (.A(net1803),
    .Y(_04721_));
 sky130_fd_sc_hd__inv_2 _11532_ (.A(net4315),
    .Y(_04722_));
 sky130_fd_sc_hd__o22a_1 _11533_ (.A1(net4091),
    .A2(_04721_),
    .B1(_04722_),
    .B2(_04460_),
    .X(_04723_));
 sky130_fd_sc_hd__o221a_1 _11534_ (.A1(_04682_),
    .A2(net4306),
    .B1(net4315),
    .B2(_04684_),
    .C1(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__nand2_1 _11535_ (.A(_04720_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__or4_1 _11536_ (.A(_04708_),
    .B(_04715_),
    .C(net4153),
    .D(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__a22o_1 _11537_ (.A1(_04679_),
    .A2(net4357),
    .B1(net4393),
    .B2(_04657_),
    .X(_04727_));
 sky130_fd_sc_hd__inv_2 _11538_ (.A(net4384),
    .Y(_04728_));
 sky130_fd_sc_hd__xnor2_1 _11539_ (.A(net4127),
    .B(net4366),
    .Y(_04729_));
 sky130_fd_sc_hd__o221a_1 _11540_ (.A1(net4138),
    .A2(_04728_),
    .B1(net4393),
    .B2(_04657_),
    .C1(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__inv_2 _11541_ (.A(net2587),
    .Y(_04731_));
 sky130_fd_sc_hd__or4_1 _11542_ (.A(net4384),
    .B(net4393),
    .C(net4366),
    .D(net2587),
    .X(_04732_));
 sky130_fd_sc_hd__o21a_1 _11543_ (.A1(net1163),
    .A2(_04732_),
    .B1(_04679_),
    .X(_04733_));
 sky130_fd_sc_hd__o2bb2a_1 _11544_ (.A1_N(_04731_),
    .A2_N(net4095),
    .B1(_04682_),
    .B2(net4384),
    .X(_04734_));
 sky130_fd_sc_hd__o221a_1 _11545_ (.A1(net4095),
    .A2(_04731_),
    .B1(_04733_),
    .B2(net4357),
    .C1(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__and3b_1 _11546_ (.A_N(_04727_),
    .B(_04730_),
    .C(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__inv_2 _11547_ (.A(net3982),
    .Y(_04737_));
 sky130_fd_sc_hd__inv_2 _11548_ (.A(net4369),
    .Y(_04738_));
 sky130_fd_sc_hd__a22o_1 _11549_ (.A1(net3983),
    .A2(_04022_),
    .B1(_04600_),
    .B2(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__xor2_1 _11550_ (.A(net4420),
    .B(_04460_),
    .X(_04740_));
 sky130_fd_sc_hd__a221o_1 _11551_ (.A1(net4354),
    .A2(_04464_),
    .B1(_04465_),
    .B2(net4369),
    .C1(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__inv_2 _11552_ (.A(net4431),
    .Y(_04742_));
 sky130_fd_sc_hd__or4_1 _11553_ (.A(net4431),
    .B(net4420),
    .C(net4369),
    .D(net4354),
    .X(_04743_));
 sky130_fd_sc_hd__o21a_1 _11554_ (.A1(net1024),
    .A2(_04743_),
    .B1(net3983),
    .X(_04744_));
 sky130_fd_sc_hd__o22a_1 _11555_ (.A1(net4354),
    .A2(_04464_),
    .B1(_04501_),
    .B2(net4431),
    .X(_04745_));
 sky130_fd_sc_hd__o221a_1 _11556_ (.A1(_04742_),
    .A2(_04467_),
    .B1(_04744_),
    .B2(_04022_),
    .C1(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__or3b_1 _11557_ (.A(_04739_),
    .B(_04741_),
    .C_N(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__nand2_1 _11558_ (.A(_04736_),
    .B(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__inv_2 _11559_ (.A(net3642),
    .Y(_04749_));
 sky130_fd_sc_hd__or2_1 _11560_ (.A(_04749_),
    .B(_04660_),
    .X(_04750_));
 sky130_fd_sc_hd__or2_1 _11561_ (.A(_04691_),
    .B(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__a21oi_1 _11562_ (.A1(net4154),
    .A2(_04748_),
    .B1(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _11563_ (.A(net1079),
    .B(net1228),
    .Y(_04753_));
 sky130_fd_sc_hd__xnor2_1 _11564_ (.A(net941),
    .B(net1918),
    .Y(_04754_));
 sky130_fd_sc_hd__xnor2_2 _11565_ (.A(_04753_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__or2_1 _11566_ (.A(net1079),
    .B(net1228),
    .X(_04756_));
 sky130_fd_sc_hd__nand2_1 _11567_ (.A(_04753_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__or2_1 _11568_ (.A(net1138),
    .B(net1122),
    .X(_04758_));
 sky130_fd_sc_hd__nand2_1 _11569_ (.A(net1138),
    .B(net1122),
    .Y(_04759_));
 sky130_fd_sc_hd__a21boi_1 _11570_ (.A1(net3189),
    .A2(_04758_),
    .B1_N(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_1 _11571_ (.A(net1105),
    .B(net1156),
    .Y(_04761_));
 sky130_fd_sc_hd__or2_1 _11572_ (.A(net1105),
    .B(net1156),
    .X(_04762_));
 sky130_fd_sc_hd__nand3_1 _11573_ (.A(net2753),
    .B(_04761_),
    .C(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21o_1 _11574_ (.A1(_04761_),
    .A2(_04762_),
    .B1(net2753),
    .X(_04764_));
 sky130_fd_sc_hd__nand2_1 _11575_ (.A(_04763_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _11576_ (.A(net1101),
    .B(net4230),
    .Y(_04766_));
 sky130_fd_sc_hd__or2_1 _11577_ (.A(net1101),
    .B(net4230),
    .X(_04767_));
 sky130_fd_sc_hd__nand3_1 _11578_ (.A(net1284),
    .B(_04766_),
    .C(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand3_1 _11579_ (.A(_04765_),
    .B(_04766_),
    .C(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__a21o_1 _11580_ (.A1(_04766_),
    .A2(_04767_),
    .B1(net1284),
    .X(_04770_));
 sky130_fd_sc_hd__nand2_1 _11581_ (.A(_04768_),
    .B(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__and2_1 _11582_ (.A(net1086),
    .B(net1851),
    .X(_04772_));
 sky130_fd_sc_hd__nor2_1 _11583_ (.A(net1086),
    .B(net1851),
    .Y(_04773_));
 sky130_fd_sc_hd__nor2_1 _11584_ (.A(_04772_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__a21oi_1 _11585_ (.A1(net2494),
    .A2(_04774_),
    .B1(_04772_),
    .Y(_04775_));
 sky130_fd_sc_hd__xnor2_1 _11586_ (.A(_04771_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nand2_1 _11587_ (.A(net1075),
    .B(net1658),
    .Y(_04777_));
 sky130_fd_sc_hd__or2_1 _11588_ (.A(net1075),
    .B(net1658),
    .X(_04778_));
 sky130_fd_sc_hd__nand3_1 _11589_ (.A(net1616),
    .B(_04777_),
    .C(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__xnor2_1 _11590_ (.A(net2494),
    .B(_04774_),
    .Y(_04780_));
 sky130_fd_sc_hd__a21oi_1 _11591_ (.A1(_04777_),
    .A2(_04779_),
    .B1(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__a21o_1 _11592_ (.A1(_04777_),
    .A2(_04778_),
    .B1(net1616),
    .X(_04782_));
 sky130_fd_sc_hd__nand2_1 _11593_ (.A(_04779_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__or2_1 _11594_ (.A(net1023),
    .B(net4312),
    .X(_04784_));
 sky130_fd_sc_hd__nand2_1 _11595_ (.A(net1023),
    .B(net4312),
    .Y(_04785_));
 sky130_fd_sc_hd__a21boi_1 _11596_ (.A1(net2474),
    .A2(_04784_),
    .B1_N(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__nor2_1 _11597_ (.A(_04783_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__nand2_1 _11598_ (.A(_04785_),
    .B(_04784_),
    .Y(_04788_));
 sky130_fd_sc_hd__xor2_1 _11599_ (.A(net2474),
    .B(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__o211a_1 _11600_ (.A1(net1008),
    .A2(net1233),
    .B1(net1046),
    .C1(net647),
    .X(_04790_));
 sky130_fd_sc_hd__a22o_1 _11601_ (.A1(net950),
    .A2(net1217),
    .B1(net1233),
    .B2(net1008),
    .X(_04791_));
 sky130_fd_sc_hd__nor2_1 _11602_ (.A(_04790_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__nor2_1 _11603_ (.A(net950),
    .B(net1217),
    .Y(_04793_));
 sky130_fd_sc_hd__or3_2 _11604_ (.A(_04789_),
    .B(_04792_),
    .C(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__xnor2_1 _11605_ (.A(_04783_),
    .B(_04786_),
    .Y(_04795_));
 sky130_fd_sc_hd__nor2_1 _11606_ (.A(_04794_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__and3_1 _11607_ (.A(_04780_),
    .B(_04777_),
    .C(_04779_),
    .X(_04797_));
 sky130_fd_sc_hd__or2_1 _11608_ (.A(_04781_),
    .B(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__inv_2 _11609_ (.A(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__o21a_1 _11610_ (.A1(_04787_),
    .A2(_04796_),
    .B1(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__nor2_1 _11611_ (.A(_04781_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _11612_ (.A(_04776_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__o21bai_2 _11613_ (.A1(_04771_),
    .A2(_04775_),
    .B1_N(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__a21oi_1 _11614_ (.A1(_04766_),
    .A2(_04768_),
    .B1(_04765_),
    .Y(_04804_));
 sky130_fd_sc_hd__a21o_1 _11615_ (.A1(_04769_),
    .A2(_04803_),
    .B1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__nand2_1 _11616_ (.A(_04758_),
    .B(_04759_),
    .Y(_04806_));
 sky130_fd_sc_hd__xor2_1 _11617_ (.A(net3189),
    .B(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__nand3_1 _11618_ (.A(_04807_),
    .B(_04761_),
    .C(_04763_),
    .Y(_04808_));
 sky130_fd_sc_hd__a21oi_1 _11619_ (.A1(_04761_),
    .A2(_04763_),
    .B1(_04807_),
    .Y(_04809_));
 sky130_fd_sc_hd__a21oi_1 _11620_ (.A1(_04805_),
    .A2(_04808_),
    .B1(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__a21o_1 _11621_ (.A1(_04757_),
    .A2(_04760_),
    .B1(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__o21a_1 _11622_ (.A1(_04757_),
    .A2(_04760_),
    .B1(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__xnor2_4 _11623_ (.A(_04755_),
    .B(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__nor2_4 _11624_ (.A(net4450),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__and2b_1 _11625_ (.A_N(_04804_),
    .B(_04769_),
    .X(_04815_));
 sky130_fd_sc_hd__xnor2_2 _11626_ (.A(_04803_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__or2_4 _11627_ (.A(_04814_),
    .B(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__clkbuf_8 _11628_ (.A(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__and2b_1 _11629_ (.A_N(_04809_),
    .B(_04808_),
    .X(_04819_));
 sky130_fd_sc_hd__xnor2_1 _11630_ (.A(_04805_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__or2_4 _11631_ (.A(_04814_),
    .B(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__and2_1 _11632_ (.A(_04776_),
    .B(_04801_),
    .X(_04822_));
 sky130_fd_sc_hd__or3_1 _11633_ (.A(_04802_),
    .B(_04814_),
    .C(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__clkbuf_8 _11634_ (.A(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__buf_4 _11635_ (.A(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__nor3_1 _11636_ (.A(_04799_),
    .B(_04787_),
    .C(_04796_),
    .Y(_04826_));
 sky130_fd_sc_hd__or3_1 _11637_ (.A(_04800_),
    .B(_04814_),
    .C(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__buf_4 _11638_ (.A(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__clkbuf_8 _11639_ (.A(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__and2_1 _11640_ (.A(_04794_),
    .B(_04795_),
    .X(_04830_));
 sky130_fd_sc_hd__or3_1 _11641_ (.A(_04796_),
    .B(_04814_),
    .C(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__buf_4 _11642_ (.A(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__or2_1 _11643_ (.A(net1136),
    .B(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__o21ai_2 _11644_ (.A1(_04792_),
    .A2(_04793_),
    .B1(_04789_),
    .Y(_04834_));
 sky130_fd_sc_hd__o211ai_4 _11645_ (.A1(net4450),
    .A2(_04813_),
    .B1(_04834_),
    .C1(_04794_),
    .Y(_04835_));
 sky130_fd_sc_hd__buf_4 _11646_ (.A(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__buf_4 _11647_ (.A(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_8 _11648_ (.A(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__a22o_1 _11649_ (.A1(net1209),
    .A2(_04828_),
    .B1(_04832_),
    .B2(net1136),
    .X(_04839_));
 sky130_fd_sc_hd__a31o_1 _11650_ (.A1(net1050),
    .A2(_04833_),
    .A3(_04838_),
    .B1(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__o221a_1 _11651_ (.A1(net1209),
    .A2(_04829_),
    .B1(_04824_),
    .B2(net1255),
    .C1(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__a221o_1 _11652_ (.A1(net1255),
    .A2(_04825_),
    .B1(_04817_),
    .B2(net1550),
    .C1(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__o221a_1 _11653_ (.A1(net5518),
    .A2(_04818_),
    .B1(_04821_),
    .B2(net5509),
    .C1(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__nor2_4 _11654_ (.A(_04814_),
    .B(_04816_),
    .Y(_04844_));
 sky130_fd_sc_hd__a21oi_4 _11655_ (.A1(net4132),
    .A2(_04701_),
    .B1(net4145),
    .Y(_04845_));
 sky130_fd_sc_hd__nor3_1 _11656_ (.A(_04796_),
    .B(_04814_),
    .C(_04830_),
    .Y(_04846_));
 sky130_fd_sc_hd__buf_4 _11657_ (.A(net88),
    .X(_04847_));
 sky130_fd_sc_hd__o211a_1 _11658_ (.A1(net7569),
    .A2(_04813_),
    .B1(_04834_),
    .C1(_04794_),
    .X(_04848_));
 sky130_fd_sc_hd__clkinv_4 _11659_ (.A(_04821_),
    .Y(_04849_));
 sky130_fd_sc_hd__nor3_1 _11660_ (.A(_04800_),
    .B(_04814_),
    .C(_04826_),
    .Y(_04850_));
 sky130_fd_sc_hd__nor3_2 _11661_ (.A(_04802_),
    .B(_04814_),
    .C(_04822_),
    .Y(_04851_));
 sky130_fd_sc_hd__or3_1 _11662_ (.A(net87),
    .B(net88),
    .C(net85),
    .X(_04852_));
 sky130_fd_sc_hd__or4_1 _11663_ (.A(_04847_),
    .B(_04848_),
    .C(_04849_),
    .D(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__inv_2 _11664_ (.A(net3405),
    .Y(_04854_));
 sky130_fd_sc_hd__nor2_1 _11665_ (.A(net3406),
    .B(net1361),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_1 _11666_ (.A(_04854_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__or2_1 _11667_ (.A(net2910),
    .B(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__or3_1 _11668_ (.A(net3151),
    .B(net3488),
    .C(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__and2_1 _11669_ (.A(net3014),
    .B(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__xnor2_1 _11670_ (.A(net3365),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__o21a_1 _11671_ (.A1(net3365),
    .A2(_04859_),
    .B1(net3423),
    .X(_04861_));
 sky130_fd_sc_hd__nor3_1 _11672_ (.A(net3423),
    .B(net3365),
    .C(_04859_),
    .Y(_04862_));
 sky130_fd_sc_hd__nor2_1 _11673_ (.A(_04861_),
    .B(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__nor2_1 _11674_ (.A(net3014),
    .B(_04858_),
    .Y(_04864_));
 sky130_fd_sc_hd__nor2_1 _11675_ (.A(_04859_),
    .B(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__o21ai_1 _11676_ (.A1(net3488),
    .A2(_04857_),
    .B1(net3151),
    .Y(_04866_));
 sky130_fd_sc_hd__nand2_1 _11677_ (.A(_04858_),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__xnor2_1 _11678_ (.A(net3488),
    .B(_04857_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_1 _11679_ (.A(net2910),
    .B(_04856_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(_04857_),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__or2_1 _11681_ (.A(_04462_),
    .B(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__o21a_1 _11682_ (.A1(net3406),
    .A2(net3641),
    .B1(net3857),
    .X(_04872_));
 sky130_fd_sc_hd__and3_1 _11683_ (.A(net3406),
    .B(net1361),
    .C(net3641),
    .X(_04873_));
 sky130_fd_sc_hd__or2_1 _11684_ (.A(_04854_),
    .B(_04855_),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _11685_ (.A(_04856_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__o32a_1 _11686_ (.A1(_04855_),
    .A2(_04872_),
    .A3(_04873_),
    .B1(_04875_),
    .B2(net3954),
    .X(_04876_));
 sky130_fd_sc_hd__a221o_1 _11687_ (.A1(net3405),
    .A2(net3954),
    .B1(_04870_),
    .B2(_04462_),
    .C1(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__a22o_1 _11688_ (.A1(_04871_),
    .A2(_04877_),
    .B1(_04868_),
    .B2(net4057),
    .X(_04878_));
 sky130_fd_sc_hd__o221a_1 _11689_ (.A1(net4057),
    .A2(_04868_),
    .B1(_04867_),
    .B2(net4105),
    .C1(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__a221o_1 _11690_ (.A1(net4105),
    .A2(_04867_),
    .B1(_04865_),
    .B2(_04467_),
    .C1(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__o221a_1 _11691_ (.A1(_04467_),
    .A2(_04865_),
    .B1(_04860_),
    .B2(_04022_),
    .C1(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__a221o_1 _11692_ (.A1(_04022_),
    .A2(_04860_),
    .B1(_04863_),
    .B2(net4132),
    .C1(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__xnor2_1 _11693_ (.A(net3388),
    .B(_04861_),
    .Y(_04883_));
 sky130_fd_sc_hd__or2_1 _11694_ (.A(net4132),
    .B(_04863_),
    .X(_04884_));
 sky130_fd_sc_hd__a31o_1 _11695_ (.A1(_04882_),
    .A2(_04883_),
    .A3(_04884_),
    .B1(net4145),
    .X(_04885_));
 sky130_fd_sc_hd__a21o_1 _11696_ (.A1(net3365),
    .A2(net3014),
    .B1(net3423),
    .X(_04886_));
 sky130_fd_sc_hd__nor2_1 _11697_ (.A(net3388),
    .B(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__nand3_1 _11698_ (.A(net3423),
    .B(net3365),
    .C(net3014),
    .Y(_04888_));
 sky130_fd_sc_hd__and2_1 _11699_ (.A(_04886_),
    .B(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__a211o_1 _11700_ (.A1(net3406),
    .A2(_04584_),
    .B1(_04502_),
    .C1(net1361),
    .X(_04890_));
 sky130_fd_sc_hd__o221a_1 _11701_ (.A1(net3405),
    .A2(net3955),
    .B1(_04584_),
    .B2(net3406),
    .C1(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__a221o_1 _11702_ (.A1(net2910),
    .A2(_04463_),
    .B1(net3955),
    .B2(net3405),
    .C1(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__o221a_1 _11703_ (.A1(net2910),
    .A2(_04464_),
    .B1(_04465_),
    .B2(net3488),
    .C1(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__a221o_1 _11704_ (.A1(net3151),
    .A2(_04684_),
    .B1(_04465_),
    .B2(net3488),
    .C1(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__o2bb2a_1 _11705_ (.A1_N(net3014),
    .A2_N(_04467_),
    .B1(_04684_),
    .B2(net3151),
    .X(_04895_));
 sky130_fd_sc_hd__xnor2_1 _11706_ (.A(net3365),
    .B(net3014),
    .Y(_04896_));
 sky130_fd_sc_hd__o22ai_1 _11707_ (.A1(net3014),
    .A2(_04467_),
    .B1(_04896_),
    .B2(net4115),
    .Y(_04897_));
 sky130_fd_sc_hd__a21oi_1 _11708_ (.A1(_04894_),
    .A2(_04895_),
    .B1(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__a22o_1 _11709_ (.A1(net4132),
    .A2(_04889_),
    .B1(_04896_),
    .B2(net4115),
    .X(_04899_));
 sky130_fd_sc_hd__o22a_1 _11710_ (.A1(net4132),
    .A2(_04889_),
    .B1(_04898_),
    .B2(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__a21oi_1 _11711_ (.A1(net4145),
    .A2(_04887_),
    .B1(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__nor2_1 _11712_ (.A(net4145),
    .B(_04887_),
    .Y(_04902_));
 sky130_fd_sc_hd__a211o_1 _11713_ (.A1(net3388),
    .A2(_04886_),
    .B1(_04901_),
    .C1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__a2111o_2 _11714_ (.A1(_04885_),
    .A2(_04903_),
    .B1(net654),
    .C1(net3388),
    .D1(_04861_),
    .X(_04904_));
 sky130_fd_sc_hd__o31a_1 _11715_ (.A1(_04844_),
    .A2(_04845_),
    .A3(_04853_),
    .B1(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__a2bb2o_1 _11716_ (.A1_N(net7569),
    .A2_N(_04905_),
    .B1(_04821_),
    .B2(net5509),
    .X(_04906_));
 sky130_fd_sc_hd__nor2_1 _11717_ (.A(_04843_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__mux2_1 _11718_ (.A0(net5356),
    .A1(net7730),
    .S(_04845_),
    .X(_04908_));
 sky130_fd_sc_hd__inv_2 _11719_ (.A(net42),
    .Y(_04909_));
 sky130_fd_sc_hd__buf_4 _11720_ (.A(net88),
    .X(_04910_));
 sky130_fd_sc_hd__clkbuf_8 _11721_ (.A(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__buf_4 _11722_ (.A(_04835_),
    .X(_04912_));
 sky130_fd_sc_hd__clkbuf_8 _11723_ (.A(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__mux2_1 _11724_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__buf_4 _11725_ (.A(_04831_),
    .X(_04915_));
 sky130_fd_sc_hd__clkbuf_8 _11726_ (.A(_04835_),
    .X(_04916_));
 sky130_fd_sc_hd__mux2_1 _11727_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__or2_1 _11728_ (.A(_04915_),
    .B(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__buf_4 _11729_ (.A(_04828_),
    .X(_04919_));
 sky130_fd_sc_hd__o211a_1 _11730_ (.A1(_04911_),
    .A2(_04914_),
    .B1(_04918_),
    .C1(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__buf_4 _11731_ (.A(_04832_),
    .X(_04921_));
 sky130_fd_sc_hd__buf_4 _11732_ (.A(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__buf_4 _11733_ (.A(_04836_),
    .X(_04923_));
 sky130_fd_sc_hd__clkbuf_8 _11734_ (.A(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04912_),
    .X(_04926_));
 sky130_fd_sc_hd__or2_1 _11737_ (.A(_04910_),
    .B(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__buf_4 _11738_ (.A(net86),
    .X(_04928_));
 sky130_fd_sc_hd__o211a_1 _11739_ (.A1(_04922_),
    .A2(_04925_),
    .B1(_04927_),
    .C1(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__buf_4 _11740_ (.A(_04832_),
    .X(_04930_));
 sky130_fd_sc_hd__mux2_1 _11741_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_04912_),
    .X(_04931_));
 sky130_fd_sc_hd__or2_1 _11742_ (.A(_04930_),
    .B(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__buf_4 _11743_ (.A(_04836_),
    .X(_04933_));
 sky130_fd_sc_hd__mux2_1 _11744_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__o21a_1 _11745_ (.A1(_04910_),
    .A2(_04934_),
    .B1(_04829_),
    .X(_04935_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04912_),
    .X(_04936_));
 sky130_fd_sc_hd__mux2_1 _11747_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04912_),
    .X(_04937_));
 sky130_fd_sc_hd__buf_4 _11748_ (.A(_04832_),
    .X(_04938_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(_04936_),
    .A1(_04937_),
    .S(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__a221o_1 _11750_ (.A1(_04932_),
    .A2(_04935_),
    .B1(_04939_),
    .B2(_04928_),
    .C1(net84),
    .X(_04940_));
 sky130_fd_sc_hd__o311a_1 _11751_ (.A1(_04825_),
    .A2(_04920_),
    .A3(_04929_),
    .B1(_04940_),
    .C1(_04844_),
    .X(_04941_));
 sky130_fd_sc_hd__buf_4 _11752_ (.A(net84),
    .X(_04942_));
 sky130_fd_sc_hd__buf_4 _11753_ (.A(_04847_),
    .X(_04943_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04924_),
    .X(_04944_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04923_),
    .X(_04945_));
 sky130_fd_sc_hd__or2_1 _11756_ (.A(_04930_),
    .B(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__buf_4 _11757_ (.A(_04829_),
    .X(_04947_));
 sky130_fd_sc_hd__o211a_1 _11758_ (.A1(_04943_),
    .A2(_04944_),
    .B1(_04946_),
    .C1(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__buf_4 _11759_ (.A(_04921_),
    .X(_04949_));
 sky130_fd_sc_hd__buf_4 _11760_ (.A(_04836_),
    .X(_04950_));
 sky130_fd_sc_hd__buf_4 _11761_ (.A(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_1 _11763_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04933_),
    .X(_04953_));
 sky130_fd_sc_hd__or2_1 _11764_ (.A(_04910_),
    .B(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__buf_4 _11765_ (.A(_04850_),
    .X(_04955_));
 sky130_fd_sc_hd__o211a_1 _11766_ (.A1(_04949_),
    .A2(_04952_),
    .B1(_04954_),
    .C1(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04933_),
    .X(_04957_));
 sky130_fd_sc_hd__or2_1 _11768_ (.A(_04921_),
    .B(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04950_),
    .X(_04959_));
 sky130_fd_sc_hd__o21a_1 _11770_ (.A1(_04847_),
    .A2(_04959_),
    .B1(_04829_),
    .X(_04960_));
 sky130_fd_sc_hd__mux2_1 _11771_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04923_),
    .X(_04961_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04923_),
    .X(_04962_));
 sky130_fd_sc_hd__mux2_1 _11773_ (.A0(_04961_),
    .A1(_04962_),
    .S(_04915_),
    .X(_04963_));
 sky130_fd_sc_hd__a221o_1 _11774_ (.A1(_04958_),
    .A2(_04960_),
    .B1(_04963_),
    .B2(_04928_),
    .C1(_04824_),
    .X(_04964_));
 sky130_fd_sc_hd__o311a_1 _11775_ (.A1(_04942_),
    .A2(_04948_),
    .A3(_04956_),
    .B1(_04964_),
    .C1(_04817_),
    .X(_04965_));
 sky130_fd_sc_hd__nor2_1 _11776_ (.A(_04941_),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__buf_4 _11777_ (.A(_04942_),
    .X(_04967_));
 sky130_fd_sc_hd__clkbuf_8 _11778_ (.A(_04836_),
    .X(_04968_));
 sky130_fd_sc_hd__mux2_1 _11779_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04837_),
    .X(_04970_));
 sky130_fd_sc_hd__mux2_1 _11781_ (.A0(_04969_),
    .A1(_04970_),
    .S(_04847_),
    .X(_04971_));
 sky130_fd_sc_hd__mux2_1 _11782_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04968_),
    .X(_04972_));
 sky130_fd_sc_hd__mux2_1 _11783_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04837_),
    .X(_04973_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(_04972_),
    .A1(_04973_),
    .S(_04921_),
    .X(_04974_));
 sky130_fd_sc_hd__mux2_1 _11785_ (.A0(_04971_),
    .A1(_04974_),
    .S(_04955_),
    .X(_04975_));
 sky130_fd_sc_hd__buf_4 _11786_ (.A(_04846_),
    .X(_04976_));
 sky130_fd_sc_hd__buf_4 _11787_ (.A(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__buf_4 _11788_ (.A(_04835_),
    .X(_04978_));
 sky130_fd_sc_hd__buf_4 _11789_ (.A(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__mux2_1 _11790_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__mux2_1 _11791_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_04978_),
    .X(_04981_));
 sky130_fd_sc_hd__or2_1 _11792_ (.A(_04938_),
    .B(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__o211a_1 _11793_ (.A1(_04977_),
    .A2(_04980_),
    .B1(_04982_),
    .C1(_04919_),
    .X(_04983_));
 sky130_fd_sc_hd__clkbuf_8 _11794_ (.A(_04938_),
    .X(_04984_));
 sky130_fd_sc_hd__mux2_1 _11795_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04979_),
    .X(_04985_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04978_),
    .X(_04986_));
 sky130_fd_sc_hd__or2_1 _11797_ (.A(_04976_),
    .B(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__clkbuf_8 _11798_ (.A(net87),
    .X(_04988_));
 sky130_fd_sc_hd__o211a_1 _11799_ (.A1(_04984_),
    .A2(_04985_),
    .B1(_04987_),
    .C1(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__o21a_1 _11800_ (.A1(_04983_),
    .A2(_04989_),
    .B1(_04825_),
    .X(_04990_));
 sky130_fd_sc_hd__clkbuf_8 _11801_ (.A(_04844_),
    .X(_04991_));
 sky130_fd_sc_hd__a211o_1 _11802_ (.A1(_04967_),
    .A2(_04975_),
    .B1(_04990_),
    .C1(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__mux2_1 _11803_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04979_),
    .X(_04993_));
 sky130_fd_sc_hd__mux2_1 _11804_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04836_),
    .X(_04994_));
 sky130_fd_sc_hd__or2_1 _11805_ (.A(_04832_),
    .B(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__o211a_1 _11806_ (.A1(_04977_),
    .A2(_04993_),
    .B1(_04995_),
    .C1(_04829_),
    .X(_04996_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04979_),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04978_),
    .X(_04998_));
 sky130_fd_sc_hd__or2_1 _11809_ (.A(_04976_),
    .B(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__o211a_1 _11810_ (.A1(_04984_),
    .A2(_04997_),
    .B1(_04999_),
    .C1(_04988_),
    .X(_05000_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04978_),
    .X(_05001_));
 sky130_fd_sc_hd__or2_1 _11812_ (.A(_04938_),
    .B(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04978_),
    .X(_05003_));
 sky130_fd_sc_hd__o21a_1 _11814_ (.A1(_04976_),
    .A2(_05003_),
    .B1(_04828_),
    .X(_05004_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04978_),
    .X(_05005_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04836_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(_05005_),
    .A1(_05006_),
    .S(_04832_),
    .X(_05007_));
 sky130_fd_sc_hd__a221o_1 _11818_ (.A1(_05002_),
    .A2(_05004_),
    .B1(_05007_),
    .B2(_04988_),
    .C1(net85),
    .X(_05008_));
 sky130_fd_sc_hd__o31a_1 _11819_ (.A1(_04825_),
    .A2(_04996_),
    .A3(_05000_),
    .B1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__o21a_1 _11820_ (.A1(_04818_),
    .A2(_05009_),
    .B1(_04821_),
    .X(_05010_));
 sky130_fd_sc_hd__a2bb2o_1 _11821_ (.A1_N(_04821_),
    .A2_N(_04966_),
    .B1(_04992_),
    .B2(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__and2_1 _11822_ (.A(_04909_),
    .B(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__clkbuf_1 _11823_ (.A(net5968),
    .X(_05013_));
 sky130_fd_sc_hd__inv_2 _11824_ (.A(net4080),
    .Y(_05014_));
 sky130_fd_sc_hd__inv_2 _11825_ (.A(net3648),
    .Y(_05015_));
 sky130_fd_sc_hd__and2_1 _11826_ (.A(net3781),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__a21oi_1 _11827_ (.A1(_05014_),
    .A2(_05016_),
    .B1(_04909_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _11828_ (.A(net3781),
    .B(_05015_),
    .Y(_05018_));
 sky130_fd_sc_hd__nand3_1 _11829_ (.A(net4271),
    .B(net4335),
    .C(net4259),
    .Y(_05019_));
 sky130_fd_sc_hd__nor3_1 _11830_ (.A(net4271),
    .B(net4335),
    .C(net4259),
    .Y(_05020_));
 sky130_fd_sc_hd__a31o_1 _11831_ (.A1(net87),
    .A2(_04976_),
    .A3(_04851_),
    .B1(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__a21oi_1 _11832_ (.A1(_04852_),
    .A2(_05019_),
    .B1(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__and3_1 _11833_ (.A(net3781),
    .B(net3648),
    .C(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__xnor2_1 _11834_ (.A(net4080),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__or4b_1 _11835_ (.A(net87),
    .B(_04977_),
    .C(_04848_),
    .D_N(net4321),
    .X(_05025_));
 sky130_fd_sc_hd__nor2_1 _11836_ (.A(net4321),
    .B(_04848_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _11837_ (.A(net1822),
    .B(net4271),
    .Y(_05027_));
 sky130_fd_sc_hd__or4_1 _11838_ (.A(net4335),
    .B(net4259),
    .C(_04824_),
    .D(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__nand2_1 _11839_ (.A(net4335),
    .B(net4259),
    .Y(_05029_));
 sky130_fd_sc_hd__or4_1 _11840_ (.A(net1822),
    .B(net4271),
    .C(_04851_),
    .D(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__a21oi_2 _11841_ (.A1(_05028_),
    .A2(_05030_),
    .B1(net4321),
    .Y(_05031_));
 sky130_fd_sc_hd__a31o_1 _11842_ (.A1(_04828_),
    .A2(_04930_),
    .A3(_05026_),
    .B1(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__or2_1 _11843_ (.A(net4079),
    .B(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__a21bo_1 _11844_ (.A1(net4080),
    .A2(_05025_),
    .B1_N(_05033_),
    .X(_05034_));
 sky130_fd_sc_hd__nor2_2 _11845_ (.A(net3781),
    .B(_05015_),
    .Y(_05035_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(_05024_),
    .A1(_05034_),
    .S(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__nand2_1 _11847_ (.A(_05018_),
    .B(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__a21bo_1 _11848_ (.A1(_05017_),
    .A2(_05037_),
    .B1_N(net7570),
    .X(_05038_));
 sky130_fd_sc_hd__o22a_2 _11849_ (.A1(net7570),
    .A2(net7731),
    .B1(_05012_),
    .B2(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__inv_2 _11850_ (.A(_04706_),
    .Y(_05040_));
 sky130_fd_sc_hd__o22a_1 _11851_ (.A1(_04707_),
    .A2(net4155),
    .B1(_05039_),
    .B2(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__nand2_1 _11852_ (.A(net4126),
    .B(net4160),
    .Y(_05042_));
 sky130_fd_sc_hd__clkbuf_4 _11853_ (.A(net4177),
    .X(_05043_));
 sky130_fd_sc_hd__or2_1 _11854_ (.A(_05043_),
    .B(net4127),
    .X(_05044_));
 sky130_fd_sc_hd__nand2_1 _11855_ (.A(_05043_),
    .B(net4127),
    .Y(_05045_));
 sky130_fd_sc_hd__and4b_1 _11856_ (.A_N(_04658_),
    .B(net4161),
    .C(_05044_),
    .D(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__o31ai_1 _11857_ (.A1(_04664_),
    .A2(_04660_),
    .A3(net4162),
    .B1(net4139),
    .Y(_05047_));
 sky130_fd_sc_hd__o21a_1 _11858_ (.A1(net4139),
    .A2(_05041_),
    .B1(net4163),
    .X(_05048_));
 sky130_fd_sc_hd__o21a_1 _11859_ (.A1(net4115),
    .A2(net4132),
    .B1(net4145),
    .X(_05049_));
 sky130_fd_sc_hd__and3_1 _11860_ (.A(net7716),
    .B(net4138),
    .C(net4177),
    .X(_05050_));
 sky130_fd_sc_hd__a21o_1 _11861_ (.A1(net5965),
    .A2(_05050_),
    .B1(net6044),
    .X(_05051_));
 sky130_fd_sc_hd__nor2_1 _11862_ (.A(net4147),
    .B(net4066),
    .Y(_05052_));
 sky130_fd_sc_hd__o221a_1 _11863_ (.A1(_04485_),
    .A2(_04653_),
    .B1(_04656_),
    .B2(_05048_),
    .C1(net4148),
    .X(_05053_));
 sky130_fd_sc_hd__buf_6 _11864_ (.A(net45),
    .X(_05054_));
 sky130_fd_sc_hd__mux2_4 _11865_ (.A0(\reg_rgb[6] ),
    .A1(_05053_),
    .S(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_1 _11866_ (.A(_05055_),
    .X(net68));
 sky130_fd_sc_hd__or2_1 _11867_ (.A(net4147),
    .B(net4066),
    .X(_05056_));
 sky130_fd_sc_hd__nor2_1 _11868_ (.A(_04023_),
    .B(_04468_),
    .Y(_05057_));
 sky130_fd_sc_hd__and4_1 _11869_ (.A(_04461_),
    .B(_04026_),
    .C(_04601_),
    .D(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__nand2_1 _11870_ (.A(net4057),
    .B(_04665_),
    .Y(_05059_));
 sky130_fd_sc_hd__o21ai_1 _11871_ (.A1(net5911),
    .A2(_04666_),
    .B1(net5205),
    .Y(_05060_));
 sky130_fd_sc_hd__and2b_1 _11872_ (.A_N(net4115),
    .B(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__or2_1 _11873_ (.A(_04667_),
    .B(net4116),
    .X(_05062_));
 sky130_fd_sc_hd__or3_1 _11874_ (.A(net5205),
    .B(net5911),
    .C(_04666_),
    .X(_05063_));
 sky130_fd_sc_hd__nor2_1 _11875_ (.A(net3917),
    .B(_04664_),
    .Y(_05064_));
 sky130_fd_sc_hd__or2_1 _11876_ (.A(_04665_),
    .B(net3918),
    .X(_05065_));
 sky130_fd_sc_hd__o2bb2a_1 _11877_ (.A1_N(_05060_),
    .A2_N(_05063_),
    .B1(net3919),
    .B2(net4057),
    .X(_05066_));
 sky130_fd_sc_hd__nand2_1 _11878_ (.A(net5205),
    .B(net5911),
    .Y(_05067_));
 sky130_fd_sc_hd__nor2_1 _11879_ (.A(net4106),
    .B(net4058),
    .Y(_05068_));
 sky130_fd_sc_hd__o22ai_1 _11880_ (.A1(net4058),
    .A2(net5912),
    .B1(net4107),
    .B2(net5205),
    .Y(_05069_));
 sky130_fd_sc_hd__and3b_1 _11881_ (.A_N(net4117),
    .B(_05066_),
    .C(net3517),
    .X(_05070_));
 sky130_fd_sc_hd__or3_1 _11882_ (.A(_04668_),
    .B(net4121),
    .C(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__and2b_1 _11883_ (.A_N(_05071_),
    .B(net3919),
    .X(_05072_));
 sky130_fd_sc_hd__and3_1 _11884_ (.A(_04666_),
    .B(net4058),
    .C(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__nand2_1 _11885_ (.A(net4105),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__and2b_1 _11886_ (.A_N(_05066_),
    .B(_05067_),
    .X(_05075_));
 sky130_fd_sc_hd__o21ba_1 _11887_ (.A1(_04667_),
    .A2(_05075_),
    .B1_N(net4116),
    .X(_05076_));
 sky130_fd_sc_hd__xnor2_4 _11888_ (.A(net4132),
    .B(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__o21ai_1 _11889_ (.A1(_05070_),
    .A2(_05077_),
    .B1(net3517),
    .Y(_05078_));
 sky130_fd_sc_hd__a21o_4 _11890_ (.A1(_05070_),
    .A2(_05077_),
    .B1(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__nor2_4 _11891_ (.A(_05074_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__and2_1 _11892_ (.A(_04684_),
    .B(net4058),
    .X(_05081_));
 sky130_fd_sc_hd__or2_1 _11893_ (.A(net4107),
    .B(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__nor2_1 _11894_ (.A(net3919),
    .B(_05071_),
    .Y(_05083_));
 sky130_fd_sc_hd__and2_1 _11895_ (.A(net4057),
    .B(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__nand2_1 _11896_ (.A(net4108),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__a21o_1 _11897_ (.A1(_05066_),
    .A2(net3517),
    .B1(_05075_),
    .X(_05086_));
 sky130_fd_sc_hd__xnor2_1 _11898_ (.A(net4117),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_2 _11899_ (.A(_05077_),
    .B(net4118),
    .Y(_05088_));
 sky130_fd_sc_hd__or2_2 _11900_ (.A(net3517),
    .B(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__nor2_4 _11901_ (.A(_05085_),
    .B(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__a21boi_1 _11902_ (.A1(_04666_),
    .A2(net4058),
    .B1_N(_05072_),
    .Y(_05091_));
 sky130_fd_sc_hd__or2b_2 _11903_ (.A(net4108),
    .B_N(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__nor2_2 _11904_ (.A(_05079_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__or4_2 _11905_ (.A(_04465_),
    .B(net3919),
    .C(_05071_),
    .D(net4108),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_4 _11906_ (.A(_05079_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__a22o_1 _11907_ (.A1(net3443),
    .A2(_05093_),
    .B1(_05095_),
    .B2(net3457),
    .X(_05096_));
 sky130_fd_sc_hd__a221o_1 _11908_ (.A1(net3461),
    .A2(_05080_),
    .B1(_05090_),
    .B2(net3348),
    .C1(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__nand2_2 _11909_ (.A(_04465_),
    .B(_05083_),
    .Y(_05098_));
 sky130_fd_sc_hd__nor2_1 _11910_ (.A(net4105),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__and2b_1 _11911_ (.A_N(_05079_),
    .B(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__nand2_1 _11912_ (.A(_04684_),
    .B(_05073_),
    .Y(_05101_));
 sky130_fd_sc_hd__nor2_4 _11913_ (.A(_05101_),
    .B(_05089_),
    .Y(_05102_));
 sky130_fd_sc_hd__nor3_4 _11914_ (.A(_04684_),
    .B(_05079_),
    .C(_05098_),
    .Y(_05103_));
 sky130_fd_sc_hd__a22o_1 _11915_ (.A1(net3370),
    .A2(_05102_),
    .B1(_05103_),
    .B2(net2898),
    .X(_05104_));
 sky130_fd_sc_hd__or2_1 _11916_ (.A(_05067_),
    .B(_05098_),
    .X(_05105_));
 sky130_fd_sc_hd__nor2_2 _11917_ (.A(_05088_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__o22a_1 _11918_ (.A1(net4058),
    .A2(_05067_),
    .B1(net4107),
    .B2(net3516),
    .X(_05107_));
 sky130_fd_sc_hd__and3_2 _11919_ (.A(_05107_),
    .B(_05077_),
    .C(_05099_),
    .X(_05108_));
 sky130_fd_sc_hd__nor2_1 _11920_ (.A(_05079_),
    .B(_05085_),
    .Y(_05109_));
 sky130_fd_sc_hd__nor2_1 _11921_ (.A(_05079_),
    .B(_05101_),
    .Y(_05110_));
 sky130_fd_sc_hd__a22o_1 _11922_ (.A1(net3990),
    .A2(_05109_),
    .B1(_05110_),
    .B2(net3389),
    .X(_05111_));
 sky130_fd_sc_hd__a221o_1 _11923_ (.A1(net4168),
    .A2(_05106_),
    .B1(_05108_),
    .B2(net3419),
    .C1(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__nor3_4 _11924_ (.A(_04501_),
    .B(_05088_),
    .C(_05092_),
    .Y(_05113_));
 sky130_fd_sc_hd__and4_4 _11925_ (.A(_05107_),
    .B(_05077_),
    .C(net4108),
    .D(_05091_),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_1 _11926_ (.A(net4118),
    .B(_05094_),
    .Y(_05115_));
 sky130_fd_sc_hd__and3b_1 _11927_ (.A_N(_05079_),
    .B(net4108),
    .C(_05091_),
    .X(_05116_));
 sky130_fd_sc_hd__a221o_1 _11928_ (.A1(net4019),
    .A2(_05115_),
    .B1(_05116_),
    .B2(net3682),
    .C1(_04659_),
    .X(_05117_));
 sky130_fd_sc_hd__a221o_1 _11929_ (.A1(net3536),
    .A2(_05113_),
    .B1(_05114_),
    .B2(net3339),
    .C1(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__a2111o_1 _11930_ (.A1(net3431),
    .A2(_05100_),
    .B1(_05104_),
    .C1(net4169),
    .D1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__nor2_1 _11931_ (.A(_04664_),
    .B(_04660_),
    .Y(_05120_));
 sky130_fd_sc_hd__or3b_1 _11932_ (.A(\gpout0.vpos[5] ),
    .B(net4126),
    .C_N(net4160),
    .X(_05121_));
 sky130_fd_sc_hd__a221o_1 _11933_ (.A1(net3372),
    .A2(_05102_),
    .B1(_05108_),
    .B2(\rbzero.debug_overlay.playerY[-5] ),
    .C1(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__a221o_1 _11934_ (.A1(net3489),
    .A2(_05113_),
    .B1(_05090_),
    .B2(net3315),
    .C1(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__a22o_1 _11935_ (.A1(net3417),
    .A2(_05106_),
    .B1(_05114_),
    .B2(net3317),
    .X(_05124_));
 sky130_fd_sc_hd__a221o_1 _11936_ (.A1(net4188),
    .A2(_05103_),
    .B1(_05115_),
    .B2(net3469),
    .C1(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__a22o_1 _11937_ (.A1(net3473),
    .A2(_05100_),
    .B1(_05109_),
    .B2(net4052),
    .X(_05126_));
 sky130_fd_sc_hd__a221o_1 _11938_ (.A1(net3445),
    .A2(_05080_),
    .B1(_05093_),
    .B2(net3326),
    .C1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__or3_1 _11939_ (.A(_05123_),
    .B(_05125_),
    .C(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__a22o_1 _11940_ (.A1(net4436),
    .A2(_05110_),
    .B1(_05116_),
    .B2(net3552),
    .X(_05129_));
 sky130_fd_sc_hd__a211o_1 _11941_ (.A1(net3433),
    .A2(_05095_),
    .B1(_05128_),
    .C1(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__or3_1 _11942_ (.A(_05100_),
    .B(_05109_),
    .C(_05110_),
    .X(_05131_));
 sky130_fd_sc_hd__a21oi_1 _11943_ (.A1(net4108),
    .A2(_05084_),
    .B1(_05073_),
    .Y(_05132_));
 sky130_fd_sc_hd__o221a_1 _11944_ (.A1(_04501_),
    .A2(_05092_),
    .B1(_05132_),
    .B2(net3517),
    .C1(_05105_),
    .X(_05133_));
 sky130_fd_sc_hd__a31o_1 _11945_ (.A1(_05074_),
    .A2(_05094_),
    .A3(_05133_),
    .B1(net4118),
    .X(_05134_));
 sky130_fd_sc_hd__or3b_4 _11946_ (.A(_05116_),
    .B(_05131_),
    .C_N(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__a22o_1 _11947_ (.A1(net3719),
    .A2(_05103_),
    .B1(_05093_),
    .B2(\rbzero.debug_overlay.facingX[0] ),
    .X(_05136_));
 sky130_fd_sc_hd__a22o_1 _11948_ (.A1(\rbzero.debug_overlay.facingX[-6] ),
    .A2(_05102_),
    .B1(_05090_),
    .B2(\rbzero.debug_overlay.facingX[-7] ),
    .X(_05137_));
 sky130_fd_sc_hd__a211o_1 _11949_ (.A1(\rbzero.debug_overlay.facingX[-9] ),
    .A2(_05106_),
    .B1(net4161),
    .C1(\gpout0.vpos[5] ),
    .X(_05138_));
 sky130_fd_sc_hd__a22o_1 _11950_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_05108_),
    .B1(_05114_),
    .B2(\rbzero.debug_overlay.facingX[-4] ),
    .X(_05139_));
 sky130_fd_sc_hd__a211o_1 _11951_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_05095_),
    .B1(_05138_),
    .C1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__a211o_1 _11952_ (.A1(\rbzero.debug_overlay.facingX[-8] ),
    .A2(_05113_),
    .B1(_05137_),
    .C1(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__a211o_1 _11953_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(_05080_),
    .B1(_05136_),
    .C1(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__a21oi_1 _11954_ (.A1(net4446),
    .A2(_05135_),
    .B1(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__a2111o_1 _11955_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_05108_),
    .B1(_04657_),
    .C1(net4126),
    .D1(net4160),
    .X(_05144_));
 sky130_fd_sc_hd__a221o_1 _11956_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(_05106_),
    .B1(_05114_),
    .B2(\rbzero.debug_overlay.facingY[-4] ),
    .C1(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__a221o_1 _11957_ (.A1(net3927),
    .A2(_05093_),
    .B1(_05095_),
    .B2(\rbzero.debug_overlay.facingY[-3] ),
    .C1(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__a22o_1 _11958_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(_05080_),
    .B1(_05103_),
    .B2(\rbzero.debug_overlay.facingY[-1] ),
    .X(_05147_));
 sky130_fd_sc_hd__a22o_1 _11959_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_05102_),
    .B1(_05090_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .X(_05148_));
 sky130_fd_sc_hd__a211o_1 _11960_ (.A1(\rbzero.debug_overlay.facingY[-8] ),
    .A2(_05113_),
    .B1(_05147_),
    .C1(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__a211o_1 _11961_ (.A1(net4002),
    .A2(_05135_),
    .B1(_05146_),
    .C1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__clkbuf_1 _11962_ (.A(net3660),
    .X(_05151_));
 sky130_fd_sc_hd__a22o_1 _11963_ (.A1(net3565),
    .A2(_05106_),
    .B1(_05114_),
    .B2(net3509),
    .X(_05152_));
 sky130_fd_sc_hd__a211o_1 _11964_ (.A1(net3661),
    .A2(_05108_),
    .B1(_05152_),
    .C1(net4160),
    .X(_05153_));
 sky130_fd_sc_hd__a221o_1 _11965_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_05093_),
    .B1(_05095_),
    .B2(\rbzero.debug_overlay.vplaneX[-3] ),
    .C1(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__clkbuf_4 _11966_ (.A(net4713),
    .X(_05155_));
 sky130_fd_sc_hd__a22o_1 _11967_ (.A1(net3493),
    .A2(_05080_),
    .B1(_05103_),
    .B2(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_05156_));
 sky130_fd_sc_hd__a22o_1 _11968_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(_05102_),
    .B1(_05090_),
    .B2(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_05157_));
 sky130_fd_sc_hd__a211o_1 _11969_ (.A1(_05155_),
    .A2(_05113_),
    .B1(_05156_),
    .C1(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__a211o_1 _11970_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_05135_),
    .B1(_05154_),
    .C1(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a21bo_1 _11971_ (.A1(net3618),
    .A2(_05108_),
    .B1_N(net4160),
    .X(_05160_));
 sky130_fd_sc_hd__a221o_1 _11972_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_05106_),
    .B1(_05114_),
    .B2(net3575),
    .C1(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__a221o_1 _11973_ (.A1(\rbzero.debug_overlay.vplaneY[0] ),
    .A2(_05093_),
    .B1(_05095_),
    .B2(\rbzero.debug_overlay.vplaneY[-3] ),
    .C1(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__a22o_1 _11974_ (.A1(net3677),
    .A2(_05080_),
    .B1(_05103_),
    .B2(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_05163_));
 sky130_fd_sc_hd__clkbuf_4 _11975_ (.A(net4598),
    .X(_05164_));
 sky130_fd_sc_hd__a22o_1 _11976_ (.A1(_05164_),
    .A2(_05113_),
    .B1(_05102_),
    .B2(net3538),
    .X(_05165_));
 sky130_fd_sc_hd__a211o_1 _11977_ (.A1(\rbzero.debug_overlay.vplaneY[-7] ),
    .A2(_05090_),
    .B1(_05163_),
    .C1(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__a211o_1 _11978_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(_05135_),
    .B1(_05162_),
    .C1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__and3_1 _11979_ (.A(_04670_),
    .B(net4127),
    .C(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__a22o_1 _11980_ (.A1(_04670_),
    .A2(_04658_),
    .B1(_05159_),
    .B2(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__o2bb2a_1 _11981_ (.A1_N(_05150_),
    .A2_N(_05169_),
    .B1(_04670_),
    .B2(net4161),
    .X(_05170_));
 sky130_fd_sc_hd__o21ai_1 _11982_ (.A1(_05143_),
    .A2(_05170_),
    .B1(_05121_),
    .Y(_05171_));
 sky130_fd_sc_hd__a21bo_1 _11983_ (.A1(_05130_),
    .A2(_05171_),
    .B1_N(_04659_),
    .X(_05172_));
 sky130_fd_sc_hd__o211a_1 _11984_ (.A1(_05097_),
    .A2(net4170),
    .B1(_05120_),
    .C1(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__inv_2 _11985_ (.A(net4139),
    .Y(_05174_));
 sky130_fd_sc_hd__a211o_1 _11986_ (.A1(_04664_),
    .A2(_05058_),
    .B1(net4171),
    .C1(net4140),
    .X(_05175_));
 sky130_fd_sc_hd__nand2_1 _11987_ (.A(net4154),
    .B(_04747_),
    .Y(_05176_));
 sky130_fd_sc_hd__a2bb2o_1 _11988_ (.A1_N(net4126),
    .A2_N(net4057),
    .B1(_04462_),
    .B2(net4160),
    .X(_05177_));
 sky130_fd_sc_hd__a21o_1 _11989_ (.A1(net4127),
    .A2(_04600_),
    .B1(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__xor2_1 _11990_ (.A(net4176),
    .B(_04460_),
    .X(_05179_));
 sky130_fd_sc_hd__o21ai_1 _11991_ (.A1(net4160),
    .A2(_04462_),
    .B1(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__o32a_1 _11992_ (.A1(_04467_),
    .A2(_05178_),
    .A3(_05180_),
    .B1(_04659_),
    .B2(net7716),
    .X(_05181_));
 sky130_fd_sc_hd__nor2_1 _11993_ (.A(net4138),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__inv_2 _11994_ (.A(net4161),
    .Y(_05183_));
 sky130_fd_sc_hd__and3_1 _11995_ (.A(_04022_),
    .B(_04467_),
    .C(_04460_),
    .X(_05184_));
 sky130_fd_sc_hd__and3_1 _11996_ (.A(net5947),
    .B(_04600_),
    .C(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__nor3_1 _11997_ (.A(net4095),
    .B(_04462_),
    .C(_05179_),
    .Y(_05186_));
 sky130_fd_sc_hd__a211o_1 _11998_ (.A1(_05183_),
    .A2(_05050_),
    .B1(net5948),
    .C1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__o2111a_1 _11999_ (.A1(_04658_),
    .A2(_05183_),
    .B1(net4177),
    .C1(_04460_),
    .D1(_04600_),
    .X(_05188_));
 sky130_fd_sc_hd__or4b_2 _12000_ (.A(_05182_),
    .B(_05187_),
    .C(_05188_),
    .D_N(_04702_),
    .X(_05189_));
 sky130_fd_sc_hd__or4_1 _12001_ (.A(net4091),
    .B(_04682_),
    .C(net4095),
    .D(_04022_),
    .X(_05190_));
 sky130_fd_sc_hd__nand2_1 _12002_ (.A(net4127),
    .B(_04468_),
    .Y(_05191_));
 sky130_fd_sc_hd__or4b_1 _12003_ (.A(net4177),
    .B(_05191_),
    .C(_04460_),
    .D_N(_04601_),
    .X(_05192_));
 sky130_fd_sc_hd__o2bb2a_1 _12004_ (.A1_N(net4095),
    .A2_N(_04600_),
    .B1(_04467_),
    .B2(net4127),
    .X(_05193_));
 sky130_fd_sc_hd__o221a_1 _12005_ (.A1(_04657_),
    .A2(_04464_),
    .B1(_04600_),
    .B2(net4095),
    .C1(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__o22a_1 _12006_ (.A1(net4177),
    .A2(_04462_),
    .B1(_04684_),
    .B2(_04682_),
    .X(_05195_));
 sky130_fd_sc_hd__o211a_1 _12007_ (.A1(net4138),
    .A2(_04460_),
    .B1(_05191_),
    .C1(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__nand2_1 _12008_ (.A(_05194_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__o21ai_1 _12009_ (.A1(_05190_),
    .A2(_05192_),
    .B1(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__and3b_1 _12010_ (.A_N(_04736_),
    .B(_05189_),
    .C(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__o21ba_1 _12011_ (.A1(_05176_),
    .A2(_05199_),
    .B1_N(_04751_),
    .X(_05200_));
 sky130_fd_sc_hd__mux2_1 _12012_ (.A0(net3569),
    .A1(net4960),
    .S(_04845_),
    .X(_05201_));
 sky130_fd_sc_hd__inv_2 _12013_ (.A(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__clkbuf_8 _12014_ (.A(net42),
    .X(_05203_));
 sky130_fd_sc_hd__buf_4 _12015_ (.A(_04977_),
    .X(_05204_));
 sky130_fd_sc_hd__mux2_1 _12016_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_04838_),
    .X(_05205_));
 sky130_fd_sc_hd__buf_4 _12017_ (.A(_04832_),
    .X(_05206_));
 sky130_fd_sc_hd__mux2_1 _12018_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04968_),
    .X(_05207_));
 sky130_fd_sc_hd__or2_1 _12019_ (.A(_05206_),
    .B(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__o211a_1 _12020_ (.A1(_05204_),
    .A2(_05205_),
    .B1(_05208_),
    .C1(_04955_),
    .X(_05209_));
 sky130_fd_sc_hd__mux2_1 _12021_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[0] ),
    .S(_04838_),
    .X(_05210_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_04979_),
    .X(_05211_));
 sky130_fd_sc_hd__or2_1 _12023_ (.A(_05206_),
    .B(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__buf_4 _12024_ (.A(_04829_),
    .X(_05213_));
 sky130_fd_sc_hd__o211a_1 _12025_ (.A1(_05204_),
    .A2(_05210_),
    .B1(_05212_),
    .C1(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__mux2_1 _12026_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_04968_),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_1 _12027_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04968_),
    .X(_05216_));
 sky130_fd_sc_hd__mux2_1 _12028_ (.A0(_05215_),
    .A1(_05216_),
    .S(_05206_),
    .X(_05217_));
 sky130_fd_sc_hd__mux2_1 _12029_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_04979_),
    .X(_05218_));
 sky130_fd_sc_hd__or2_1 _12030_ (.A(_04984_),
    .B(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__buf_4 _12031_ (.A(_04978_),
    .X(_05220_));
 sky130_fd_sc_hd__mux2_1 _12032_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__o21a_1 _12033_ (.A1(_04977_),
    .A2(_05221_),
    .B1(_04988_),
    .X(_05222_));
 sky130_fd_sc_hd__a221o_1 _12034_ (.A1(_05213_),
    .A2(_05217_),
    .B1(_05219_),
    .B2(_05222_),
    .C1(_04825_),
    .X(_05223_));
 sky130_fd_sc_hd__o311a_1 _12035_ (.A1(_04967_),
    .A2(_05209_),
    .A3(_05214_),
    .B1(_04818_),
    .C1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__mux2_1 _12036_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_04838_),
    .X(_05225_));
 sky130_fd_sc_hd__mux2_1 _12037_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_04979_),
    .X(_05226_));
 sky130_fd_sc_hd__or2_1 _12038_ (.A(_05206_),
    .B(_05226_),
    .X(_05227_));
 sky130_fd_sc_hd__o211a_1 _12039_ (.A1(_05204_),
    .A2(_05225_),
    .B1(_05227_),
    .C1(_04955_),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _12040_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_04838_),
    .X(_05229_));
 sky130_fd_sc_hd__mux2_1 _12041_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_04979_),
    .X(_05230_));
 sky130_fd_sc_hd__or2_1 _12042_ (.A(_05206_),
    .B(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__o211a_1 _12043_ (.A1(_05204_),
    .A2(_05229_),
    .B1(_05231_),
    .C1(_05213_),
    .X(_05232_));
 sky130_fd_sc_hd__buf_4 _12044_ (.A(_04988_),
    .X(_05233_));
 sky130_fd_sc_hd__mux2_1 _12045_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_05220_),
    .X(_05234_));
 sky130_fd_sc_hd__mux2_1 _12046_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_05220_),
    .X(_05235_));
 sky130_fd_sc_hd__mux2_1 _12047_ (.A0(_05234_),
    .A1(_05235_),
    .S(_05206_),
    .X(_05236_));
 sky130_fd_sc_hd__clkbuf_8 _12048_ (.A(_04916_),
    .X(_05237_));
 sky130_fd_sc_hd__mux2_1 _12049_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__buf_4 _12050_ (.A(_04835_),
    .X(_05239_));
 sky130_fd_sc_hd__mux2_1 _12051_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__or2_1 _12052_ (.A(_04938_),
    .B(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__o211a_1 _12053_ (.A1(_04911_),
    .A2(_05238_),
    .B1(_05241_),
    .C1(_04919_),
    .X(_05242_));
 sky130_fd_sc_hd__a211o_1 _12054_ (.A1(_05233_),
    .A2(_05236_),
    .B1(_05242_),
    .C1(_04825_),
    .X(_05243_));
 sky130_fd_sc_hd__o311a_1 _12055_ (.A1(_04967_),
    .A2(_05228_),
    .A3(_05232_),
    .B1(_04991_),
    .C1(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__mux2_1 _12056_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04838_),
    .X(_05245_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_05220_),
    .X(_05246_));
 sky130_fd_sc_hd__or2_1 _12058_ (.A(_04977_),
    .B(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__o211a_1 _12059_ (.A1(_04949_),
    .A2(_05245_),
    .B1(_05247_),
    .C1(_05233_),
    .X(_05248_));
 sky130_fd_sc_hd__clkbuf_8 _12060_ (.A(_04923_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_8 _12061_ (.A(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__mux2_1 _12062_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__mux2_1 _12063_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_05237_),
    .X(_05252_));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(_04984_),
    .B(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__o211a_1 _12065_ (.A1(_05204_),
    .A2(_05251_),
    .B1(_05253_),
    .C1(_05213_),
    .X(_05254_));
 sky130_fd_sc_hd__mux2_1 _12066_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_05249_),
    .X(_05255_));
 sky130_fd_sc_hd__mux2_1 _12067_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_05249_),
    .X(_05256_));
 sky130_fd_sc_hd__mux2_1 _12068_ (.A0(_05255_),
    .A1(_05256_),
    .S(_04984_),
    .X(_05257_));
 sky130_fd_sc_hd__buf_4 _12069_ (.A(_04933_),
    .X(_05258_));
 sky130_fd_sc_hd__mux2_1 _12070_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__mux2_1 _12071_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_04923_),
    .X(_05260_));
 sky130_fd_sc_hd__or2_1 _12072_ (.A(_04930_),
    .B(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__o211a_1 _12073_ (.A1(_04943_),
    .A2(_05259_),
    .B1(_05261_),
    .C1(_04947_),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_8 _12074_ (.A(_04824_),
    .X(_05263_));
 sky130_fd_sc_hd__a211o_1 _12075_ (.A1(_05233_),
    .A2(_05257_),
    .B1(_05262_),
    .C1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__o311a_1 _12076_ (.A1(_04967_),
    .A2(_05248_),
    .A3(_05254_),
    .B1(_04818_),
    .C1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__mux2_1 _12077_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_04979_),
    .X(_05266_));
 sky130_fd_sc_hd__mux2_1 _12078_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_04979_),
    .X(_05267_));
 sky130_fd_sc_hd__mux2_1 _12079_ (.A0(_05266_),
    .A1(_05267_),
    .S(_05206_),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_1 _12080_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_05237_),
    .X(_05269_));
 sky130_fd_sc_hd__or2_1 _12081_ (.A(_04984_),
    .B(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__mux2_1 _12082_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_04913_),
    .X(_05271_));
 sky130_fd_sc_hd__o21a_1 _12083_ (.A1(_04911_),
    .A2(_05271_),
    .B1(_04988_),
    .X(_05272_));
 sky130_fd_sc_hd__a221o_1 _12084_ (.A1(_05213_),
    .A2(_05268_),
    .B1(_05270_),
    .B2(_05272_),
    .C1(_04942_),
    .X(_05273_));
 sky130_fd_sc_hd__mux2_1 _12085_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_05220_),
    .X(_05274_));
 sky130_fd_sc_hd__or2_1 _12086_ (.A(_04977_),
    .B(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__clkbuf_8 _12087_ (.A(_04930_),
    .X(_05276_));
 sky130_fd_sc_hd__mux2_1 _12088_ (.A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_04913_),
    .X(_05277_));
 sky130_fd_sc_hd__o21a_1 _12089_ (.A1(_05276_),
    .A2(_05277_),
    .B1(_04988_),
    .X(_05278_));
 sky130_fd_sc_hd__mux2_1 _12090_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_05220_),
    .X(_05279_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_05220_),
    .X(_05280_));
 sky130_fd_sc_hd__mux2_1 _12092_ (.A0(_05279_),
    .A1(_05280_),
    .S(_04977_),
    .X(_05281_));
 sky130_fd_sc_hd__a221o_1 _12093_ (.A1(_05275_),
    .A2(_05278_),
    .B1(_05281_),
    .B2(_05213_),
    .C1(_04825_),
    .X(_05282_));
 sky130_fd_sc_hd__a31o_1 _12094_ (.A1(_04991_),
    .A2(_05273_),
    .A3(_05282_),
    .B1(_04821_),
    .X(_05283_));
 sky130_fd_sc_hd__o32a_1 _12095_ (.A1(_04849_),
    .A2(_05224_),
    .A3(_05244_),
    .B1(_05265_),
    .B2(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__nand2_1 _12096_ (.A(net4080),
    .B(_05032_),
    .Y(_05285_));
 sky130_fd_sc_hd__a221o_1 _12097_ (.A1(_05014_),
    .A2(_05023_),
    .B1(_05285_),
    .B2(_05035_),
    .C1(_05016_),
    .X(_05286_));
 sky130_fd_sc_hd__and2_1 _12098_ (.A(net1822),
    .B(_04991_),
    .X(_05287_));
 sky130_fd_sc_hd__nor2_1 _12099_ (.A(net1822),
    .B(_04991_),
    .Y(_05288_));
 sky130_fd_sc_hd__o31a_1 _12100_ (.A1(_05018_),
    .A2(_05287_),
    .A3(_05288_),
    .B1(_05203_),
    .X(_05289_));
 sky130_fd_sc_hd__a2bb2o_1 _12101_ (.A1_N(_05203_),
    .A2_N(_05284_),
    .B1(_05286_),
    .B2(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__mux2_1 _12102_ (.A0(_05202_),
    .A1(_05290_),
    .S(net7570),
    .X(_05291_));
 sky130_fd_sc_hd__a2bb2o_1 _12103_ (.A1_N(_04707_),
    .A2_N(_05200_),
    .B1(_05291_),
    .B2(_04706_),
    .X(_05292_));
 sky130_fd_sc_hd__nand2_1 _12104_ (.A(net4140),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__a21oi_1 _12105_ (.A1(net4172),
    .A2(_05293_),
    .B1(_04656_),
    .Y(_05294_));
 sky130_fd_sc_hd__a211o_1 _12106_ (.A1(net3774),
    .A2(net2),
    .B1(net4067),
    .C1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__inv_2 _12107_ (.A(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__mux2_4 _12108_ (.A0(\reg_rgb[7] ),
    .A1(_05296_),
    .S(_05054_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_1 _12109_ (.A(_05297_),
    .X(net69));
 sky130_fd_sc_hd__mux2_1 _12110_ (.A0(net4964),
    .A1(net7722),
    .S(_04845_),
    .X(_05298_));
 sky130_fd_sc_hd__mux2_1 _12111_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_04951_),
    .X(_05299_));
 sky130_fd_sc_hd__or2_1 _12112_ (.A(_04949_),
    .B(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_1 _12113_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04951_),
    .X(_05301_));
 sky130_fd_sc_hd__o21a_1 _12114_ (.A1(_04943_),
    .A2(_05301_),
    .B1(_04947_),
    .X(_05302_));
 sky130_fd_sc_hd__mux2_1 _12115_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_05258_),
    .X(_05303_));
 sky130_fd_sc_hd__mux2_1 _12116_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_05258_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_1 _12117_ (.A0(_05303_),
    .A1(_05304_),
    .S(_05276_),
    .X(_05305_));
 sky130_fd_sc_hd__buf_4 _12118_ (.A(_04955_),
    .X(_05306_));
 sky130_fd_sc_hd__a221o_1 _12119_ (.A1(_05300_),
    .A2(_05302_),
    .B1(_05305_),
    .B2(_05306_),
    .C1(_05263_),
    .X(_05307_));
 sky130_fd_sc_hd__mux2_1 _12120_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04951_),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _12121_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04951_),
    .X(_05309_));
 sky130_fd_sc_hd__mux2_1 _12122_ (.A0(_05308_),
    .A1(_05309_),
    .S(_04911_),
    .X(_05310_));
 sky130_fd_sc_hd__mux2_1 _12123_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_04838_),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_04837_),
    .X(_05312_));
 sky130_fd_sc_hd__or2_1 _12125_ (.A(_04921_),
    .B(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__o211a_1 _12126_ (.A1(_05204_),
    .A2(_05311_),
    .B1(_05313_),
    .C1(_05213_),
    .X(_05314_));
 sky130_fd_sc_hd__a211o_1 _12127_ (.A1(_05306_),
    .A2(_05310_),
    .B1(_05314_),
    .C1(_04967_),
    .X(_05315_));
 sky130_fd_sc_hd__mux2_1 _12128_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_04950_),
    .X(_05316_));
 sky130_fd_sc_hd__or2_1 _12129_ (.A(_04921_),
    .B(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__mux2_1 _12130_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04950_),
    .X(_05318_));
 sky130_fd_sc_hd__o21a_1 _12131_ (.A1(_04847_),
    .A2(_05318_),
    .B1(_04829_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _12132_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04933_),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04933_),
    .X(_05321_));
 sky130_fd_sc_hd__mux2_1 _12134_ (.A0(_05320_),
    .A1(_05321_),
    .S(_04915_),
    .X(_05322_));
 sky130_fd_sc_hd__a221o_1 _12135_ (.A1(_05317_),
    .A2(_05319_),
    .B1(_05322_),
    .B2(_04928_),
    .C1(_04942_),
    .X(_05323_));
 sky130_fd_sc_hd__mux2_1 _12136_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04950_),
    .X(_05324_));
 sky130_fd_sc_hd__mux2_1 _12137_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_04950_),
    .X(_05325_));
 sky130_fd_sc_hd__mux2_1 _12138_ (.A0(_05324_),
    .A1(_05325_),
    .S(_04910_),
    .X(_05326_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_04837_),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_1 _12140_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_04836_),
    .X(_05328_));
 sky130_fd_sc_hd__or2_1 _12141_ (.A(_04832_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__o211a_1 _12142_ (.A1(_04847_),
    .A2(_05327_),
    .B1(_05329_),
    .C1(_04829_),
    .X(_05330_));
 sky130_fd_sc_hd__a211o_1 _12143_ (.A1(_04955_),
    .A2(_05326_),
    .B1(_05330_),
    .C1(_04824_),
    .X(_05331_));
 sky130_fd_sc_hd__a31o_1 _12144_ (.A1(_04991_),
    .A2(_05323_),
    .A3(_05331_),
    .B1(_04849_),
    .X(_05332_));
 sky130_fd_sc_hd__a31o_1 _12145_ (.A1(_04818_),
    .A2(_05307_),
    .A3(_05315_),
    .B1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__mux2_1 _12146_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_05220_),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _12147_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04978_),
    .X(_05335_));
 sky130_fd_sc_hd__or2_1 _12148_ (.A(_04938_),
    .B(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__o211a_1 _12149_ (.A1(_04911_),
    .A2(_05334_),
    .B1(_05336_),
    .C1(_04919_),
    .X(_05337_));
 sky130_fd_sc_hd__mux2_1 _12150_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04913_),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _12151_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_05239_),
    .X(_05339_));
 sky130_fd_sc_hd__or2_1 _12152_ (.A(_04976_),
    .B(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__o211a_1 _12153_ (.A1(_05276_),
    .A2(_05338_),
    .B1(_05340_),
    .C1(_04928_),
    .X(_05341_));
 sky130_fd_sc_hd__mux2_1 _12154_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04916_),
    .X(_05342_));
 sky130_fd_sc_hd__or2_1 _12155_ (.A(_04915_),
    .B(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__mux2_1 _12156_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04912_),
    .X(_05344_));
 sky130_fd_sc_hd__o21a_1 _12157_ (.A1(_04910_),
    .A2(_05344_),
    .B1(_04828_),
    .X(_05345_));
 sky130_fd_sc_hd__mux2_1 _12158_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_05239_),
    .X(_05346_));
 sky130_fd_sc_hd__mux2_1 _12159_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_05239_),
    .X(_05347_));
 sky130_fd_sc_hd__mux2_1 _12160_ (.A0(_05346_),
    .A1(_05347_),
    .S(_04938_),
    .X(_05348_));
 sky130_fd_sc_hd__a221o_1 _12161_ (.A1(_05343_),
    .A2(_05345_),
    .B1(_05348_),
    .B2(_04988_),
    .C1(_04824_),
    .X(_05349_));
 sky130_fd_sc_hd__o311a_1 _12162_ (.A1(_04942_),
    .A2(_05337_),
    .A3(_05341_),
    .B1(_05349_),
    .C1(_04817_),
    .X(_05350_));
 sky130_fd_sc_hd__mux2_1 _12163_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_05237_),
    .X(_05351_));
 sky130_fd_sc_hd__mux2_1 _12164_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_05239_),
    .X(_05352_));
 sky130_fd_sc_hd__or2_1 _12165_ (.A(_04915_),
    .B(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__o211a_1 _12166_ (.A1(_04911_),
    .A2(_05351_),
    .B1(_05353_),
    .C1(_04919_),
    .X(_05354_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_05249_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _12168_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04916_),
    .X(_05356_));
 sky130_fd_sc_hd__or2_1 _12169_ (.A(_04910_),
    .B(_05356_),
    .X(_05357_));
 sky130_fd_sc_hd__o211a_1 _12170_ (.A1(_05276_),
    .A2(_05355_),
    .B1(_05357_),
    .C1(_04928_),
    .X(_05358_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_04916_),
    .X(_05359_));
 sky130_fd_sc_hd__or2_1 _12172_ (.A(_04915_),
    .B(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04923_),
    .X(_05361_));
 sky130_fd_sc_hd__o21a_1 _12174_ (.A1(_04910_),
    .A2(_05361_),
    .B1(_04828_),
    .X(_05362_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_05239_),
    .X(_05363_));
 sky130_fd_sc_hd__mux2_1 _12176_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_05239_),
    .X(_05364_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(_05363_),
    .A1(_05364_),
    .S(_04938_),
    .X(_05365_));
 sky130_fd_sc_hd__a221o_1 _12178_ (.A1(_05360_),
    .A2(_05362_),
    .B1(_05365_),
    .B2(_04988_),
    .C1(net85),
    .X(_05366_));
 sky130_fd_sc_hd__o311a_1 _12179_ (.A1(_04825_),
    .A2(_05354_),
    .A3(_05358_),
    .B1(_05366_),
    .C1(_04844_),
    .X(_05367_));
 sky130_fd_sc_hd__or3_2 _12180_ (.A(_04821_),
    .B(_05350_),
    .C(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__buf_4 _12181_ (.A(_05258_),
    .X(_05369_));
 sky130_fd_sc_hd__o31a_1 _12182_ (.A1(_05213_),
    .A2(_04949_),
    .A3(_05369_),
    .B1(_05025_),
    .X(_05370_));
 sky130_fd_sc_hd__o21ai_1 _12183_ (.A1(_05031_),
    .A2(_05370_),
    .B1(net4080),
    .Y(_05371_));
 sky130_fd_sc_hd__a21o_1 _12184_ (.A1(net4080),
    .A2(_05021_),
    .B1(_05015_),
    .X(_05372_));
 sky130_fd_sc_hd__a32o_1 _12185_ (.A1(_05033_),
    .A2(_05035_),
    .A3(_05371_),
    .B1(_05372_),
    .B2(net3781),
    .X(_05373_));
 sky130_fd_sc_hd__a32o_1 _12186_ (.A1(_04909_),
    .A2(_05333_),
    .A3(_05368_),
    .B1(_05373_),
    .B2(_05017_),
    .X(_05374_));
 sky130_fd_sc_hd__mux2_2 _12187_ (.A0(net7723),
    .A1(_05374_),
    .S(net7570),
    .X(_05375_));
 sky130_fd_sc_hd__and2_1 _12188_ (.A(_05040_),
    .B(_04691_),
    .X(_05376_));
 sky130_fd_sc_hd__a211o_1 _12189_ (.A1(_04706_),
    .A2(_05375_),
    .B1(_05376_),
    .C1(net4139),
    .X(_05377_));
 sky130_fd_sc_hd__a21o_1 _12190_ (.A1(net4163),
    .A2(_05377_),
    .B1(_04656_),
    .X(_05378_));
 sky130_fd_sc_hd__o211a_1 _12191_ (.A1(net3976),
    .A2(_04653_),
    .B1(net4148),
    .C1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_2 _12192_ (.A0(\reg_rgb[14] ),
    .A1(_05379_),
    .S(_05054_),
    .X(_05380_));
 sky130_fd_sc_hd__buf_1 _12193_ (.A(_05380_),
    .X(net64));
 sky130_fd_sc_hd__mux2_1 _12194_ (.A0(net7733),
    .A1(net4952),
    .S(_04845_),
    .X(_05381_));
 sky130_fd_sc_hd__mux2_1 _12195_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_05249_),
    .X(_05382_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_04912_),
    .X(_05383_));
 sky130_fd_sc_hd__or2_1 _12197_ (.A(_04910_),
    .B(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__o211a_1 _12198_ (.A1(_05276_),
    .A2(_05382_),
    .B1(_05384_),
    .C1(_04928_),
    .X(_05385_));
 sky130_fd_sc_hd__mux2_1 _12199_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_04924_),
    .X(_05386_));
 sky130_fd_sc_hd__mux2_1 _12200_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_04923_),
    .X(_05387_));
 sky130_fd_sc_hd__or2_1 _12201_ (.A(_04930_),
    .B(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__o211a_1 _12202_ (.A1(_04943_),
    .A2(_05386_),
    .B1(_05388_),
    .C1(_04947_),
    .X(_05389_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_04916_),
    .X(_05390_));
 sky130_fd_sc_hd__mux2_1 _12204_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[0] ),
    .S(_04916_),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_1 _12205_ (.A0(_05390_),
    .A1(_05391_),
    .S(_04938_),
    .X(_05392_));
 sky130_fd_sc_hd__mux2_1 _12206_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_04923_),
    .X(_05393_));
 sky130_fd_sc_hd__or2_1 _12207_ (.A(_04930_),
    .B(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__mux2_1 _12208_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_04950_),
    .X(_05395_));
 sky130_fd_sc_hd__o21a_1 _12209_ (.A1(_04847_),
    .A2(_05395_),
    .B1(net86),
    .X(_05396_));
 sky130_fd_sc_hd__a221o_1 _12210_ (.A1(_04947_),
    .A2(_05392_),
    .B1(_05394_),
    .B2(_05396_),
    .C1(net84),
    .X(_05397_));
 sky130_fd_sc_hd__o311a_1 _12211_ (.A1(_05263_),
    .A2(_05385_),
    .A3(_05389_),
    .B1(_05397_),
    .C1(_04817_),
    .X(_05398_));
 sky130_fd_sc_hd__mux2_1 _12212_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04924_),
    .X(_05399_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_04923_),
    .X(_05400_));
 sky130_fd_sc_hd__or2_1 _12214_ (.A(_04930_),
    .B(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__o211a_1 _12215_ (.A1(_04943_),
    .A2(_05399_),
    .B1(_05401_),
    .C1(_04928_),
    .X(_05402_));
 sky130_fd_sc_hd__mux2_1 _12216_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_04951_),
    .X(_05403_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_04933_),
    .X(_05404_));
 sky130_fd_sc_hd__or2_1 _12218_ (.A(_04921_),
    .B(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__o211a_1 _12219_ (.A1(_04943_),
    .A2(_05403_),
    .B1(_05405_),
    .C1(_04947_),
    .X(_05406_));
 sky130_fd_sc_hd__mux2_1 _12220_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_04950_),
    .X(_05407_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04950_),
    .X(_05408_));
 sky130_fd_sc_hd__mux2_1 _12222_ (.A0(_05407_),
    .A1(_05408_),
    .S(_04930_),
    .X(_05409_));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_04837_),
    .X(_05410_));
 sky130_fd_sc_hd__mux2_1 _12224_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04836_),
    .X(_05411_));
 sky130_fd_sc_hd__or2_1 _12225_ (.A(net88),
    .B(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__o211a_1 _12226_ (.A1(_04921_),
    .A2(_05410_),
    .B1(_05412_),
    .C1(_04829_),
    .X(_05413_));
 sky130_fd_sc_hd__a211o_1 _12227_ (.A1(_04955_),
    .A2(_05409_),
    .B1(_05413_),
    .C1(_04824_),
    .X(_05414_));
 sky130_fd_sc_hd__o311a_1 _12228_ (.A1(_04942_),
    .A2(_05402_),
    .A3(_05406_),
    .B1(_04844_),
    .C1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__mux2_1 _12229_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_04838_),
    .X(_05416_));
 sky130_fd_sc_hd__mux2_1 _12230_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_04837_),
    .X(_05417_));
 sky130_fd_sc_hd__or2_1 _12231_ (.A(_04847_),
    .B(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__o211a_1 _12232_ (.A1(_04949_),
    .A2(_05416_),
    .B1(_05418_),
    .C1(_05213_),
    .X(_05419_));
 sky130_fd_sc_hd__mux2_1 _12233_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_04838_),
    .X(_05420_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_04837_),
    .X(_05421_));
 sky130_fd_sc_hd__or2_1 _12235_ (.A(_04921_),
    .B(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__o211a_1 _12236_ (.A1(_05204_),
    .A2(_05420_),
    .B1(_05422_),
    .C1(_04955_),
    .X(_05423_));
 sky130_fd_sc_hd__mux2_1 _12237_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_04968_),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _12238_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_04968_),
    .X(_05425_));
 sky130_fd_sc_hd__mux2_1 _12239_ (.A0(_05424_),
    .A1(_05425_),
    .S(_04847_),
    .X(_05426_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_04968_),
    .X(_05427_));
 sky130_fd_sc_hd__mux2_1 _12241_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_04836_),
    .X(_05428_));
 sky130_fd_sc_hd__or2_1 _12242_ (.A(_04832_),
    .B(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__o211a_1 _12243_ (.A1(_04977_),
    .A2(_05427_),
    .B1(_05429_),
    .C1(_04988_),
    .X(_05430_));
 sky130_fd_sc_hd__a211o_1 _12244_ (.A1(_05213_),
    .A2(_05426_),
    .B1(_05430_),
    .C1(_04825_),
    .X(_05431_));
 sky130_fd_sc_hd__o311a_1 _12245_ (.A1(_04967_),
    .A2(_05419_),
    .A3(_05423_),
    .B1(_04818_),
    .C1(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04950_),
    .X(_05433_));
 sky130_fd_sc_hd__mux2_1 _12247_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04933_),
    .X(_05434_));
 sky130_fd_sc_hd__mux2_1 _12248_ (.A0(_05433_),
    .A1(_05434_),
    .S(_04915_),
    .X(_05435_));
 sky130_fd_sc_hd__mux2_1 _12249_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_04837_),
    .X(_05436_));
 sky130_fd_sc_hd__or2_1 _12250_ (.A(_04921_),
    .B(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__mux2_1 _12251_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04968_),
    .X(_05438_));
 sky130_fd_sc_hd__o21a_1 _12252_ (.A1(_04977_),
    .A2(_05438_),
    .B1(net87),
    .X(_05439_));
 sky130_fd_sc_hd__a221o_1 _12253_ (.A1(_04947_),
    .A2(_05435_),
    .B1(_05437_),
    .B2(_05439_),
    .C1(_04942_),
    .X(_05440_));
 sky130_fd_sc_hd__mux2_1 _12254_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04933_),
    .X(_05441_));
 sky130_fd_sc_hd__mux2_1 _12255_ (.A0(\rbzero.tex_g1[63] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_04933_),
    .X(_05442_));
 sky130_fd_sc_hd__mux2_1 _12256_ (.A0(_05441_),
    .A1(_05442_),
    .S(_04910_),
    .X(_05443_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_04837_),
    .X(_05444_));
 sky130_fd_sc_hd__or2_1 _12258_ (.A(_04847_),
    .B(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_04968_),
    .X(_05446_));
 sky130_fd_sc_hd__o21a_1 _12260_ (.A1(_05206_),
    .A2(_05446_),
    .B1(_04829_),
    .X(_05447_));
 sky130_fd_sc_hd__a221o_1 _12261_ (.A1(_04955_),
    .A2(_05443_),
    .B1(_05445_),
    .B2(_05447_),
    .C1(_04824_),
    .X(_05448_));
 sky130_fd_sc_hd__a31o_1 _12262_ (.A1(_04991_),
    .A2(_05440_),
    .A3(_05448_),
    .B1(_04821_),
    .X(_05449_));
 sky130_fd_sc_hd__o32a_1 _12263_ (.A1(_04849_),
    .A2(_05398_),
    .A3(_05415_),
    .B1(_05432_),
    .B2(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__a21oi_1 _12264_ (.A1(net4335),
    .A2(_05306_),
    .B1(_05018_),
    .Y(_05451_));
 sky130_fd_sc_hd__o21ai_1 _12265_ (.A1(net4335),
    .A2(_05306_),
    .B1(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__o311a_1 _12266_ (.A1(net3781),
    .A2(_05015_),
    .A3(_05285_),
    .B1(_05452_),
    .C1(net42),
    .X(_05453_));
 sky130_fd_sc_hd__o21ba_1 _12267_ (.A1(_05203_),
    .A2(_05450_),
    .B1_N(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__mux2_1 _12268_ (.A0(net7734),
    .A1(_05454_),
    .S(net7570),
    .X(_05455_));
 sky130_fd_sc_hd__nor2_1 _12269_ (.A(_04736_),
    .B(_05176_),
    .Y(_05456_));
 sky130_fd_sc_hd__nor2_1 _12270_ (.A(_04751_),
    .B(_05198_),
    .Y(_05457_));
 sky130_fd_sc_hd__a31o_1 _12271_ (.A1(_05189_),
    .A2(_05456_),
    .A3(_05457_),
    .B1(_04707_),
    .X(_05458_));
 sky130_fd_sc_hd__o21ai_1 _12272_ (.A1(_05040_),
    .A2(_05455_),
    .B1(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__nand2_1 _12273_ (.A(net4140),
    .B(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__a21o_1 _12274_ (.A1(net4172),
    .A2(_05460_),
    .B1(_04656_),
    .X(_05461_));
 sky130_fd_sc_hd__o211a_1 _12275_ (.A1(net3871),
    .A2(_04653_),
    .B1(net4148),
    .C1(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__mux2_4 _12276_ (.A0(\reg_rgb[15] ),
    .A1(_05462_),
    .S(_05054_),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_1 _12277_ (.A(_05463_),
    .X(net65));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(net5049),
    .A1(net7719),
    .S(_04845_),
    .X(_05464_));
 sky130_fd_sc_hd__clkbuf_8 _12279_ (.A(_04947_),
    .X(_05465_));
 sky130_fd_sc_hd__mux2_1 _12280_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_05237_),
    .X(_05466_));
 sky130_fd_sc_hd__mux2_1 _12281_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_05237_),
    .X(_05467_));
 sky130_fd_sc_hd__mux2_1 _12282_ (.A0(_05466_),
    .A1(_05467_),
    .S(_05206_),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _12283_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_04913_),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04916_),
    .X(_05470_));
 sky130_fd_sc_hd__or2_1 _12285_ (.A(_04976_),
    .B(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__o211a_1 _12286_ (.A1(_05276_),
    .A2(_05469_),
    .B1(_05471_),
    .C1(_04928_),
    .X(_05472_));
 sky130_fd_sc_hd__a211o_1 _12287_ (.A1(_05465_),
    .A2(_05468_),
    .B1(_05472_),
    .C1(_04942_),
    .X(_05473_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_05237_),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_1 _12289_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_05220_),
    .X(_05475_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(_05474_),
    .A1(_05475_),
    .S(_05206_),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_1 _12291_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_04913_),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_04916_),
    .X(_05478_));
 sky130_fd_sc_hd__or2_1 _12293_ (.A(_04976_),
    .B(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__o211a_1 _12294_ (.A1(_05276_),
    .A2(_05477_),
    .B1(_05479_),
    .C1(_04919_),
    .X(_05480_));
 sky130_fd_sc_hd__a211o_1 _12295_ (.A1(_05233_),
    .A2(_05476_),
    .B1(_05480_),
    .C1(_05263_),
    .X(_05481_));
 sky130_fd_sc_hd__mux2_1 _12296_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_05220_),
    .X(_05482_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_04978_),
    .X(_05483_));
 sky130_fd_sc_hd__or2_1 _12298_ (.A(_04938_),
    .B(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__o211a_1 _12299_ (.A1(_04911_),
    .A2(_05482_),
    .B1(_05484_),
    .C1(_04919_),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _12300_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_04913_),
    .X(_05486_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_05239_),
    .X(_05487_));
 sky130_fd_sc_hd__or2_1 _12302_ (.A(_04915_),
    .B(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__o211a_1 _12303_ (.A1(_04911_),
    .A2(_05486_),
    .B1(_05488_),
    .C1(_04928_),
    .X(_05489_));
 sky130_fd_sc_hd__mux2_1 _12304_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04916_),
    .X(_05490_));
 sky130_fd_sc_hd__or2_1 _12305_ (.A(_04976_),
    .B(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__mux2_1 _12306_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_04912_),
    .X(_05492_));
 sky130_fd_sc_hd__o21a_1 _12307_ (.A1(_04930_),
    .A2(_05492_),
    .B1(net86),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _12308_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_05239_),
    .X(_05494_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_05239_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _12310_ (.A0(_05494_),
    .A1(_05495_),
    .S(_04976_),
    .X(_05496_));
 sky130_fd_sc_hd__a221o_1 _12311_ (.A1(_05491_),
    .A2(_05493_),
    .B1(_05496_),
    .B2(_04919_),
    .C1(net84),
    .X(_05497_));
 sky130_fd_sc_hd__o311a_1 _12312_ (.A1(_04825_),
    .A2(_05485_),
    .A3(_05489_),
    .B1(_05497_),
    .C1(_04844_),
    .X(_05498_));
 sky130_fd_sc_hd__a31o_1 _12313_ (.A1(_04818_),
    .A2(_05473_),
    .A3(_05481_),
    .B1(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _12314_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_04913_),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _12315_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_05237_),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(_05500_),
    .A1(_05501_),
    .S(_04984_),
    .X(_05502_));
 sky130_fd_sc_hd__mux2_1 _12317_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_05249_),
    .X(_05503_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04912_),
    .X(_05504_));
 sky130_fd_sc_hd__or2_1 _12319_ (.A(_04915_),
    .B(_05504_),
    .X(_05505_));
 sky130_fd_sc_hd__o211a_1 _12320_ (.A1(_04911_),
    .A2(_05503_),
    .B1(_05505_),
    .C1(_04919_),
    .X(_05506_));
 sky130_fd_sc_hd__a211o_1 _12321_ (.A1(_05233_),
    .A2(_05502_),
    .B1(_05506_),
    .C1(_04942_),
    .X(_05507_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_05237_),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_1 _12323_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_05237_),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(_05508_),
    .A1(_05509_),
    .S(_04984_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _12325_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_05249_),
    .X(_05511_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_04912_),
    .X(_05512_));
 sky130_fd_sc_hd__or2_1 _12327_ (.A(_04915_),
    .B(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__o211a_1 _12328_ (.A1(_04911_),
    .A2(_05511_),
    .B1(_05513_),
    .C1(_04919_),
    .X(_05514_));
 sky130_fd_sc_hd__a211o_1 _12329_ (.A1(_05233_),
    .A2(_05510_),
    .B1(_05514_),
    .C1(_05263_),
    .X(_05515_));
 sky130_fd_sc_hd__a31o_1 _12330_ (.A1(_04991_),
    .A2(_05507_),
    .A3(_05515_),
    .B1(_04821_),
    .X(_05516_));
 sky130_fd_sc_hd__buf_4 _12331_ (.A(_04943_),
    .X(_05517_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_05250_),
    .X(_05518_));
 sky130_fd_sc_hd__mux2_1 _12333_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_04913_),
    .X(_05519_));
 sky130_fd_sc_hd__or2_1 _12334_ (.A(_05276_),
    .B(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__o211a_1 _12335_ (.A1(_05517_),
    .A2(_05518_),
    .B1(_05520_),
    .C1(_05233_),
    .X(_05521_));
 sky130_fd_sc_hd__mux2_1 _12336_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_05369_),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _12337_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_05249_),
    .X(_05523_));
 sky130_fd_sc_hd__or2_1 _12338_ (.A(_05276_),
    .B(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__o211a_1 _12339_ (.A1(_05517_),
    .A2(_05522_),
    .B1(_05524_),
    .C1(_05465_),
    .X(_05525_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_05249_),
    .X(_05526_));
 sky130_fd_sc_hd__or2_1 _12341_ (.A(_04922_),
    .B(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_05258_),
    .X(_05528_));
 sky130_fd_sc_hd__o21a_1 _12343_ (.A1(_04943_),
    .A2(_05528_),
    .B1(_04947_),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_05249_),
    .X(_05530_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04913_),
    .X(_05531_));
 sky130_fd_sc_hd__mux2_1 _12346_ (.A0(_05530_),
    .A1(_05531_),
    .S(_04984_),
    .X(_05532_));
 sky130_fd_sc_hd__a221o_1 _12347_ (.A1(_05527_),
    .A2(_05529_),
    .B1(_05532_),
    .B2(_05233_),
    .C1(_04942_),
    .X(_05533_));
 sky130_fd_sc_hd__o311a_1 _12348_ (.A1(_05263_),
    .A2(_05521_),
    .A3(_05525_),
    .B1(_05533_),
    .C1(_04818_),
    .X(_05534_));
 sky130_fd_sc_hd__o22a_1 _12349_ (.A1(_04849_),
    .A2(_05499_),
    .B1(_05516_),
    .B2(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__a31o_1 _12350_ (.A1(_05306_),
    .A2(_05517_),
    .A3(_04848_),
    .B1(_05033_),
    .X(_05536_));
 sky130_fd_sc_hd__o21bai_1 _12351_ (.A1(net4080),
    .A2(_05021_),
    .B1_N(_05372_),
    .Y(_05537_));
 sky130_fd_sc_hd__a32o_1 _12352_ (.A1(_05035_),
    .A2(_05285_),
    .A3(_05536_),
    .B1(_05537_),
    .B2(net3781),
    .X(_05538_));
 sky130_fd_sc_hd__a22o_1 _12353_ (.A1(_04909_),
    .A2(_05535_),
    .B1(_05538_),
    .B2(_05017_),
    .X(_05539_));
 sky130_fd_sc_hd__mux2_1 _12354_ (.A0(net7720),
    .A1(_05539_),
    .S(net7570),
    .X(_05540_));
 sky130_fd_sc_hd__o21ai_1 _12355_ (.A1(_05189_),
    .A2(_05198_),
    .B1(_05456_),
    .Y(_05541_));
 sky130_fd_sc_hd__or3b_1 _12356_ (.A(_04706_),
    .B(_04750_),
    .C_N(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__o21ai_1 _12357_ (.A1(_05040_),
    .A2(_05540_),
    .B1(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__o21ai_1 _12358_ (.A1(_05376_),
    .A2(_05543_),
    .B1(net4140),
    .Y(_05544_));
 sky130_fd_sc_hd__nor2_1 _12359_ (.A(_04656_),
    .B(net4067),
    .Y(_05545_));
 sky130_fd_sc_hd__and3_1 _12360_ (.A(net4163),
    .B(_05544_),
    .C(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__mux2_2 _12361_ (.A0(\reg_rgb[22] ),
    .A1(_05546_),
    .S(_05054_),
    .X(_05547_));
 sky130_fd_sc_hd__clkbuf_1 _12362_ (.A(_05547_),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(net7725),
    .A1(net4956),
    .S(_04845_),
    .X(_05548_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_05250_),
    .X(_05549_));
 sky130_fd_sc_hd__mux2_1 _12365_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_05250_),
    .X(_05550_));
 sky130_fd_sc_hd__mux2_1 _12366_ (.A0(_05549_),
    .A1(_05550_),
    .S(_04949_),
    .X(_05551_));
 sky130_fd_sc_hd__mux2_1 _12367_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_05369_),
    .X(_05552_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_05258_),
    .X(_05553_));
 sky130_fd_sc_hd__or2_1 _12369_ (.A(_04922_),
    .B(_05553_),
    .X(_05554_));
 sky130_fd_sc_hd__o211a_1 _12370_ (.A1(_05517_),
    .A2(_05552_),
    .B1(_05554_),
    .C1(_05465_),
    .X(_05555_));
 sky130_fd_sc_hd__a211o_1 _12371_ (.A1(_05306_),
    .A2(_05551_),
    .B1(_05555_),
    .C1(_04967_),
    .X(_05556_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_05250_),
    .X(_05557_));
 sky130_fd_sc_hd__mux2_1 _12373_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_05250_),
    .X(_05558_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(_05557_),
    .A1(_05558_),
    .S(_04949_),
    .X(_05559_));
 sky130_fd_sc_hd__mux2_1 _12375_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_05369_),
    .X(_05560_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_04924_),
    .X(_05561_));
 sky130_fd_sc_hd__or2_1 _12377_ (.A(_04922_),
    .B(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__o211a_1 _12378_ (.A1(_05517_),
    .A2(_05560_),
    .B1(_05562_),
    .C1(_05465_),
    .X(_05563_));
 sky130_fd_sc_hd__a211o_1 _12379_ (.A1(_05306_),
    .A2(_05559_),
    .B1(_05563_),
    .C1(_05263_),
    .X(_05564_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_05369_),
    .X(_05565_));
 sky130_fd_sc_hd__mux2_1 _12381_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_04924_),
    .X(_05566_));
 sky130_fd_sc_hd__or2_1 _12382_ (.A(_04922_),
    .B(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__o211a_1 _12383_ (.A1(_05517_),
    .A2(_05565_),
    .B1(_05567_),
    .C1(_05465_),
    .X(_05568_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_05369_),
    .X(_05569_));
 sky130_fd_sc_hd__mux2_1 _12385_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_05258_),
    .X(_05570_));
 sky130_fd_sc_hd__or2_1 _12386_ (.A(_04922_),
    .B(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__o211a_1 _12387_ (.A1(_05517_),
    .A2(_05569_),
    .B1(_05571_),
    .C1(_05306_),
    .X(_05572_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04951_),
    .X(_05573_));
 sky130_fd_sc_hd__or2_1 _12389_ (.A(_04949_),
    .B(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04838_),
    .X(_05575_));
 sky130_fd_sc_hd__o21a_1 _12391_ (.A1(_05204_),
    .A2(_05575_),
    .B1(_04955_),
    .X(_05576_));
 sky130_fd_sc_hd__mux2_1 _12392_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04951_),
    .X(_05577_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04951_),
    .X(_05578_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(_05577_),
    .A1(_05578_),
    .S(_05276_),
    .X(_05579_));
 sky130_fd_sc_hd__a221o_1 _12395_ (.A1(_05574_),
    .A2(_05576_),
    .B1(_05579_),
    .B2(_05465_),
    .C1(_05263_),
    .X(_05580_));
 sky130_fd_sc_hd__o311a_1 _12396_ (.A1(_04967_),
    .A2(_05568_),
    .A3(_05572_),
    .B1(_04818_),
    .C1(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__a311o_1 _12397_ (.A1(_04991_),
    .A2(_05556_),
    .A3(_05564_),
    .B1(_04849_),
    .C1(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_05250_),
    .X(_05583_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_05250_),
    .X(_05584_));
 sky130_fd_sc_hd__mux2_1 _12400_ (.A0(_05583_),
    .A1(_05584_),
    .S(_05204_),
    .X(_05585_));
 sky130_fd_sc_hd__mux2_1 _12401_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_05369_),
    .X(_05586_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04924_),
    .X(_05587_));
 sky130_fd_sc_hd__or2_1 _12403_ (.A(_04922_),
    .B(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__o211a_1 _12404_ (.A1(_05517_),
    .A2(_05586_),
    .B1(_05588_),
    .C1(_05306_),
    .X(_05589_));
 sky130_fd_sc_hd__a211o_1 _12405_ (.A1(_05465_),
    .A2(_05585_),
    .B1(_05589_),
    .C1(_04967_),
    .X(_05590_));
 sky130_fd_sc_hd__mux2_1 _12406_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_05250_),
    .X(_05591_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_05250_),
    .X(_05592_));
 sky130_fd_sc_hd__mux2_1 _12408_ (.A0(_05591_),
    .A1(_05592_),
    .S(_05204_),
    .X(_05593_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_05369_),
    .X(_05594_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04924_),
    .X(_05595_));
 sky130_fd_sc_hd__or2_1 _12411_ (.A(_04922_),
    .B(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__o211a_1 _12412_ (.A1(_05517_),
    .A2(_05594_),
    .B1(_05596_),
    .C1(_05306_),
    .X(_05597_));
 sky130_fd_sc_hd__a211o_1 _12413_ (.A1(_05465_),
    .A2(_05593_),
    .B1(_05597_),
    .C1(_05263_),
    .X(_05598_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_05369_),
    .X(_05599_));
 sky130_fd_sc_hd__mux2_1 _12415_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04924_),
    .X(_05600_));
 sky130_fd_sc_hd__or2_1 _12416_ (.A(_04922_),
    .B(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__o211a_1 _12417_ (.A1(_05517_),
    .A2(_05599_),
    .B1(_05601_),
    .C1(_05233_),
    .X(_05602_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_05369_),
    .X(_05603_));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_05258_),
    .X(_05604_));
 sky130_fd_sc_hd__or2_1 _12420_ (.A(_04943_),
    .B(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__o211a_1 _12421_ (.A1(_04949_),
    .A2(_05603_),
    .B1(_05605_),
    .C1(_05465_),
    .X(_05606_));
 sky130_fd_sc_hd__mux2_1 _12422_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_05258_),
    .X(_05607_));
 sky130_fd_sc_hd__or2_1 _12423_ (.A(_04922_),
    .B(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04951_),
    .X(_05609_));
 sky130_fd_sc_hd__o21a_1 _12425_ (.A1(_04943_),
    .A2(_05609_),
    .B1(_04947_),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_05258_),
    .X(_05611_));
 sky130_fd_sc_hd__mux2_1 _12427_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04924_),
    .X(_05612_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(_05611_),
    .A1(_05612_),
    .S(_04984_),
    .X(_05613_));
 sky130_fd_sc_hd__a221o_1 _12429_ (.A1(_05608_),
    .A2(_05610_),
    .B1(_05613_),
    .B2(_05233_),
    .C1(_04967_),
    .X(_05614_));
 sky130_fd_sc_hd__o311a_1 _12430_ (.A1(_05263_),
    .A2(_05602_),
    .A3(_05606_),
    .B1(_05614_),
    .C1(_04991_),
    .X(_05615_));
 sky130_fd_sc_hd__a311o_1 _12431_ (.A1(_04818_),
    .A2(_05590_),
    .A3(_05598_),
    .B1(_04821_),
    .C1(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__o31a_1 _12432_ (.A1(net4080),
    .A2(_05015_),
    .A3(_05021_),
    .B1(net3781),
    .X(_05617_));
 sky130_fd_sc_hd__a21oi_1 _12433_ (.A1(_05465_),
    .A2(_04949_),
    .B1(_05031_),
    .Y(_05618_));
 sky130_fd_sc_hd__o21a_1 _12434_ (.A1(_05031_),
    .A2(_05026_),
    .B1(net4080),
    .X(_05619_));
 sky130_fd_sc_hd__o21a_1 _12435_ (.A1(_05618_),
    .A2(_05619_),
    .B1(_05035_),
    .X(_05620_));
 sky130_fd_sc_hd__and2_1 _12436_ (.A(net4321),
    .B(_04848_),
    .X(_05621_));
 sky130_fd_sc_hd__nor2_1 _12437_ (.A(_05026_),
    .B(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__o221a_1 _12438_ (.A1(_05617_),
    .A2(_05620_),
    .B1(_05622_),
    .B2(_05018_),
    .C1(_05203_),
    .X(_05623_));
 sky130_fd_sc_hd__a31o_1 _12439_ (.A1(_04909_),
    .A2(_05582_),
    .A3(_05616_),
    .B1(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__mux2_1 _12440_ (.A0(net7726),
    .A1(_05624_),
    .S(net7570),
    .X(_05625_));
 sky130_fd_sc_hd__or3_1 _12441_ (.A(_04706_),
    .B(_04751_),
    .C(_05541_),
    .X(_05626_));
 sky130_fd_sc_hd__a21bo_1 _12442_ (.A1(_04706_),
    .A2(_05625_),
    .B1_N(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__o211a_1 _12443_ (.A1(net4139),
    .A2(_05627_),
    .B1(_05545_),
    .C1(net4172),
    .X(_05628_));
 sky130_fd_sc_hd__mux2_2 _12444_ (.A0(\reg_rgb[23] ),
    .A1(_05628_),
    .S(_05054_),
    .X(_05629_));
 sky130_fd_sc_hd__clkbuf_1 _12445_ (.A(_05629_),
    .X(net67));
 sky130_fd_sc_hd__mux2_4 _12446_ (.A0(reg_vsync),
    .A1(_04477_),
    .S(_05054_),
    .X(_05630_));
 sky130_fd_sc_hd__clkbuf_1 _12447_ (.A(_05630_),
    .X(net74));
 sky130_fd_sc_hd__inv_2 _12448_ (.A(\rbzero.hsync ),
    .Y(_05631_));
 sky130_fd_sc_hd__mux2_2 _12449_ (.A0(reg_hsync),
    .A1(_05631_),
    .S(_05054_),
    .X(_05632_));
 sky130_fd_sc_hd__clkbuf_1 _12450_ (.A(_05632_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 _12451_ (.A(net4),
    .X(_05633_));
 sky130_fd_sc_hd__nor2_1 _12452_ (.A(_05633_),
    .B(net4156),
    .Y(_05634_));
 sky130_fd_sc_hd__inv_2 _12453_ (.A(net7),
    .Y(_05635_));
 sky130_fd_sc_hd__a211o_1 _12454_ (.A1(_05633_),
    .A2(net4068),
    .B1(net8),
    .C1(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__mux4_1 _12455_ (.A0(net4149),
    .A1(net4141),
    .A2(net4164),
    .A3(net7727),
    .S0(_05633_),
    .S1(net7),
    .X(_05637_));
 sky130_fd_sc_hd__a2bb2o_1 _12456_ (.A1_N(_05634_),
    .A2_N(_05636_),
    .B1(_05637_),
    .B2(net8),
    .X(_05638_));
 sky130_fd_sc_hd__and4b_1 _12457_ (.A_N(net9),
    .B(_05638_),
    .C(net5),
    .D(net6),
    .X(_05639_));
 sky130_fd_sc_hd__nor2_1 _12458_ (.A(net9),
    .B(net8),
    .Y(_05640_));
 sky130_fd_sc_hd__nor2_1 _12459_ (.A(net7),
    .B(net6),
    .Y(_05641_));
 sky130_fd_sc_hd__and2b_1 _12460_ (.A_N(net5),
    .B(_05633_),
    .X(_05642_));
 sky130_fd_sc_hd__and2_1 _12461_ (.A(net5),
    .B(net4),
    .X(_05643_));
 sky130_fd_sc_hd__and2b_1 _12462_ (.A_N(_05633_),
    .B(net5),
    .X(_05644_));
 sky130_fd_sc_hd__buf_1 _12463_ (.A(clknet_4_8__leaf_i_clk),
    .X(_05645_));
 sky130_fd_sc_hd__nor2_2 _12464_ (.A(net5),
    .B(_05633_),
    .Y(_05646_));
 sky130_fd_sc_hd__a221o_2 _12465_ (.A1(net6122),
    .A2(_05643_),
    .B1(_05644_),
    .B2(clknet_1_1__leaf__05645_),
    .C1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__a21o_2 _12466_ (.A1(_04102_),
    .A2(_05642_),
    .B1(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__inv_2 _12467_ (.A(net6),
    .Y(_05649_));
 sky130_fd_sc_hd__nor2_1 _12468_ (.A(net7),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__a22o_1 _12469_ (.A1(net52),
    .A2(_05646_),
    .B1(_05642_),
    .B2(net53),
    .X(_05651_));
 sky130_fd_sc_hd__a221o_1 _12470_ (.A1(net54),
    .A2(_05643_),
    .B1(_05644_),
    .B2(net55),
    .C1(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__a22o_2 _12471_ (.A1(_05641_),
    .A2(_05648_),
    .B1(_05650_),
    .B2(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__mux4_1 _12472_ (.A0(_04648_),
    .A1(_04461_),
    .A2(_04468_),
    .A3(_04023_),
    .S0(_05633_),
    .S1(net5),
    .X(_05654_));
 sky130_fd_sc_hd__mux2_1 _12473_ (.A0(net4133),
    .A1(net4089),
    .S(_05633_),
    .X(_05655_));
 sky130_fd_sc_hd__mux4_1 _12474_ (.A0(_04020_),
    .A1(_04495_),
    .A2(_04494_),
    .A3(_04500_),
    .S0(_05633_),
    .S1(net5),
    .X(_05656_));
 sky130_fd_sc_hd__mux2_1 _12475_ (.A0(_05655_),
    .A1(_05656_),
    .S(net7),
    .X(_05657_));
 sky130_fd_sc_hd__a21o_1 _12476_ (.A1(net5),
    .A2(net6),
    .B1(net7),
    .X(_05658_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(net8),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__a21o_1 _12478_ (.A1(net7),
    .A2(net6),
    .B1(net8),
    .X(_05660_));
 sky130_fd_sc_hd__o2111a_1 _12479_ (.A1(_05649_),
    .A2(_05657_),
    .B1(_05659_),
    .C1(_05660_),
    .D1(net9),
    .X(_05661_));
 sky130_fd_sc_hd__o21a_1 _12480_ (.A1(net6),
    .A2(_05654_),
    .B1(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__a221o_1 _12481_ (.A1(net50),
    .A2(_05643_),
    .B1(_05644_),
    .B2(net49),
    .C1(_05649_),
    .X(_05663_));
 sky130_fd_sc_hd__a221o_1 _12482_ (.A1(net4066),
    .A2(_05646_),
    .B1(_05642_),
    .B2(net71),
    .C1(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__a22o_1 _12483_ (.A1(_05203_),
    .A2(_05643_),
    .B1(_05644_),
    .B2(net41),
    .X(_05665_));
 sky130_fd_sc_hd__a221o_1 _12484_ (.A1(net51),
    .A2(_05646_),
    .B1(_05642_),
    .B2(net40),
    .C1(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__a21bo_1 _12485_ (.A1(_05649_),
    .A2(_05666_),
    .B1_N(net7),
    .X(_05667_));
 sky130_fd_sc_hd__a21bo_1 _12486_ (.A1(net44),
    .A2(_05644_),
    .B1_N(_05641_),
    .X(_05668_));
 sky130_fd_sc_hd__a22o_1 _12487_ (.A1(net43),
    .A2(_05646_),
    .B1(_05642_),
    .B2(net46),
    .X(_05669_));
 sky130_fd_sc_hd__a211o_1 _12488_ (.A1(net4147),
    .A2(_05643_),
    .B1(_05668_),
    .C1(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__and3b_1 _12489_ (.A_N(net8),
    .B(_05670_),
    .C(net9),
    .X(_05671_));
 sky130_fd_sc_hd__clkbuf_1 _12490_ (.A(net4110),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_4 _12491_ (.A(net4095),
    .X(_05673_));
 sky130_fd_sc_hd__clkbuf_1 _12492_ (.A(net4138),
    .X(_05674_));
 sky130_fd_sc_hd__clkbuf_1 _12493_ (.A(net7716),
    .X(_05675_));
 sky130_fd_sc_hd__mux4_1 _12494_ (.A0(net4111),
    .A1(_05673_),
    .A2(net4071),
    .A3(net4092),
    .S0(_05633_),
    .S1(net6),
    .X(_05676_));
 sky130_fd_sc_hd__buf_1 _12495_ (.A(net4102),
    .X(_05677_));
 sky130_fd_sc_hd__clkbuf_1 _12496_ (.A(net5981),
    .X(_05678_));
 sky130_fd_sc_hd__mux4_1 _12497_ (.A0(net4103),
    .A1(net4024),
    .A2(net5965),
    .A3(net6044),
    .S0(net4),
    .S1(net7),
    .X(_05679_));
 sky130_fd_sc_hd__clkbuf_2 _12498_ (.A(net4127),
    .X(_05680_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(net4128),
    .A1(_05043_),
    .S(net4),
    .X(_05681_));
 sky130_fd_sc_hd__mux2_1 _12500_ (.A0(_05679_),
    .A1(_05681_),
    .S(_05649_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _12501_ (.A0(_05676_),
    .A1(_05682_),
    .S(net5),
    .X(_05683_));
 sky130_fd_sc_hd__and4_1 _12502_ (.A(net9),
    .B(net8),
    .C(_05658_),
    .D(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__a31o_1 _12503_ (.A1(_05664_),
    .A2(_05667_),
    .A3(_05671_),
    .B1(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__a211o_2 _12504_ (.A1(_05640_),
    .A2(_05653_),
    .B1(_05662_),
    .C1(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__nand4b_1 _12505_ (.A_N(net4149),
    .B(_05641_),
    .C(_05640_),
    .D(_05646_),
    .Y(_05687_));
 sky130_fd_sc_hd__o21a_2 _12506_ (.A1(_05639_),
    .A2(_05686_),
    .B1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_2 _12507_ (.A0(\reg_gpout[0] ),
    .A1(clknet_1_1__leaf__05688_),
    .S(_05054_),
    .X(_05689_));
 sky130_fd_sc_hd__buf_1 _12508_ (.A(_05689_),
    .X(net56));
 sky130_fd_sc_hd__and2b_1 _12509_ (.A_N(net14),
    .B(net13),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_4 _12510_ (.A(net10),
    .X(_05691_));
 sky130_fd_sc_hd__or2_1 _12511_ (.A(_05691_),
    .B(net4156),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _12512_ (.A(_05691_),
    .B(net7571),
    .Y(_05693_));
 sky130_fd_sc_hd__mux4_1 _12513_ (.A0(net4149),
    .A1(net4141),
    .A2(net4164),
    .A3(net7727),
    .S0(_05691_),
    .S1(net13),
    .X(_05694_));
 sky130_fd_sc_hd__a32o_1 _12514_ (.A1(_05690_),
    .A2(_05692_),
    .A3(_05693_),
    .B1(_05694_),
    .B2(net14),
    .X(_05695_));
 sky130_fd_sc_hd__and4b_1 _12515_ (.A_N(net15),
    .B(_05695_),
    .C(net11),
    .D(net12),
    .X(_05696_));
 sky130_fd_sc_hd__nand2_1 _12516_ (.A(net11),
    .B(_05691_),
    .Y(_05697_));
 sky130_fd_sc_hd__inv_2 _12517_ (.A(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__and2b_1 _12518_ (.A_N(net11),
    .B(_05691_),
    .X(_05699_));
 sky130_fd_sc_hd__and2b_2 _12519_ (.A_N(net10),
    .B(net11),
    .X(_05700_));
 sky130_fd_sc_hd__nor2_2 _12520_ (.A(net11),
    .B(_05691_),
    .Y(_05701_));
 sky130_fd_sc_hd__a22o_1 _12521_ (.A1(net41),
    .A2(_05700_),
    .B1(_05701_),
    .B2(net51),
    .X(_05702_));
 sky130_fd_sc_hd__a221o_1 _12522_ (.A1(_05203_),
    .A2(_05698_),
    .B1(_05699_),
    .B2(net40),
    .C1(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__inv_2 _12523_ (.A(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21a_1 _12524_ (.A1(net12),
    .A2(_05704_),
    .B1(net13),
    .X(_05705_));
 sky130_fd_sc_hd__or2_1 _12525_ (.A(net13),
    .B(net12),
    .X(_05706_));
 sky130_fd_sc_hd__a221o_1 _12526_ (.A1(net43),
    .A2(_05701_),
    .B1(_05699_),
    .B2(net46),
    .C1(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__and2b_1 _12527_ (.A_N(net13),
    .B(net12),
    .X(_05708_));
 sky130_fd_sc_hd__a31o_1 _12528_ (.A1(net54),
    .A2(_05698_),
    .A3(_05708_),
    .B1(net15),
    .X(_05709_));
 sky130_fd_sc_hd__nand2_1 _12529_ (.A(_05707_),
    .B(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__inv_2 _12530_ (.A(net49),
    .Y(_05711_));
 sky130_fd_sc_hd__inv_2 _12531_ (.A(_05700_),
    .Y(_05712_));
 sky130_fd_sc_hd__nor2_1 _12532_ (.A(net14),
    .B(net15),
    .Y(_05713_));
 sky130_fd_sc_hd__a21oi_1 _12533_ (.A1(net54),
    .A2(_05713_),
    .B1(net50),
    .Y(_05714_));
 sky130_fd_sc_hd__o221a_1 _12534_ (.A1(_05711_),
    .A2(_05712_),
    .B1(_05697_),
    .B2(_05714_),
    .C1(net12),
    .X(_05715_));
 sky130_fd_sc_hd__a22o_1 _12535_ (.A1(net55),
    .A2(_05700_),
    .B1(_05701_),
    .B2(net52),
    .X(_05716_));
 sky130_fd_sc_hd__a21o_1 _12536_ (.A1(net53),
    .A2(_05699_),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__nor2_1 _12537_ (.A(net13),
    .B(net12),
    .Y(_05718_));
 sky130_fd_sc_hd__o221a_2 _12538_ (.A1(clknet_1_1__leaf__05645_),
    .A2(_05712_),
    .B1(_05697_),
    .B2(net6100),
    .C1(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__a21oi_2 _12539_ (.A1(_05708_),
    .A2(_05717_),
    .B1(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__o32a_2 _12540_ (.A1(_05705_),
    .A2(_05710_),
    .A3(_05715_),
    .B1(_05720_),
    .B2(net15),
    .X(_05721_));
 sky130_fd_sc_hd__a22o_1 _12541_ (.A1(_04021_),
    .A2(_05701_),
    .B1(_05699_),
    .B2(_04495_),
    .X(_05722_));
 sky130_fd_sc_hd__a221o_1 _12542_ (.A1(_04494_),
    .A2(_05700_),
    .B1(_05698_),
    .B2(_04500_),
    .C1(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__a22o_1 _12543_ (.A1(net4066),
    .A2(_05701_),
    .B1(_05699_),
    .B2(net71),
    .X(_05724_));
 sky130_fd_sc_hd__a22o_1 _12544_ (.A1(net44),
    .A2(_05700_),
    .B1(_05698_),
    .B2(net4147),
    .X(_05725_));
 sky130_fd_sc_hd__a22o_1 _12545_ (.A1(_05708_),
    .A2(_05724_),
    .B1(_05725_),
    .B2(_05718_),
    .X(_05726_));
 sky130_fd_sc_hd__mux4_1 _12546_ (.A0(_04648_),
    .A1(net4133),
    .A2(_04461_),
    .A3(net4089),
    .S0(net12),
    .S1(_05691_),
    .X(_05727_));
 sky130_fd_sc_hd__mux4_1 _12547_ (.A0(net4111),
    .A1(_05673_),
    .A2(net4071),
    .A3(net4092),
    .S0(_05691_),
    .S1(net12),
    .X(_05728_));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(_05727_),
    .A1(_05728_),
    .S(net13),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_4 _12549_ (.A(net5965),
    .X(_05730_));
 sky130_fd_sc_hd__buf_1 _12550_ (.A(net6044),
    .X(_05731_));
 sky130_fd_sc_hd__mux4_1 _12551_ (.A0(net4128),
    .A1(_05043_),
    .A2(_05730_),
    .A3(net3996),
    .S0(_05691_),
    .S1(net12),
    .X(_05732_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(net4102),
    .A1(net4024),
    .S(net10),
    .X(_05733_));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(_04468_),
    .A1(_04023_),
    .S(_05691_),
    .X(_05734_));
 sky130_fd_sc_hd__a22o_1 _12554_ (.A1(_05708_),
    .A2(_05733_),
    .B1(_05734_),
    .B2(_05718_),
    .X(_05735_));
 sky130_fd_sc_hd__a21o_1 _12555_ (.A1(net13),
    .A2(_05732_),
    .B1(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(_05729_),
    .A1(_05736_),
    .S(net11),
    .X(_05737_));
 sky130_fd_sc_hd__mux2_1 _12557_ (.A0(_05726_),
    .A1(_05737_),
    .S(net14),
    .X(_05738_));
 sky130_fd_sc_hd__a31o_1 _12558_ (.A1(net12),
    .A2(_05690_),
    .A3(_05723_),
    .B1(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__a2bb2o_2 _12559_ (.A1_N(net14),
    .A2_N(_05721_),
    .B1(_05739_),
    .B2(net15),
    .X(_05740_));
 sky130_fd_sc_hd__nand3_1 _12560_ (.A(_05701_),
    .B(_05718_),
    .C(_05713_),
    .Y(_05741_));
 sky130_fd_sc_hd__o22a_2 _12561_ (.A1(_05696_),
    .A2(_05740_),
    .B1(_05741_),
    .B2(net4141),
    .X(_05742_));
 sky130_fd_sc_hd__mux2_2 _12562_ (.A0(\reg_gpout[1] ),
    .A1(clknet_1_0__leaf__05742_),
    .S(_05054_),
    .X(_05743_));
 sky130_fd_sc_hd__buf_1 _12563_ (.A(_05743_),
    .X(net57));
 sky130_fd_sc_hd__nor2_1 _12564_ (.A(net17),
    .B(net16),
    .Y(_05744_));
 sky130_fd_sc_hd__nor2_1 _12565_ (.A(net19),
    .B(net18),
    .Y(_05745_));
 sky130_fd_sc_hd__nand2_1 _12566_ (.A(_05744_),
    .B(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__buf_2 _12567_ (.A(net17),
    .X(_05747_));
 sky130_fd_sc_hd__inv_2 _12568_ (.A(net21),
    .Y(_05748_));
 sky130_fd_sc_hd__clkbuf_4 _12569_ (.A(net16),
    .X(_05749_));
 sky130_fd_sc_hd__nor2_1 _12570_ (.A(_05749_),
    .B(net4156),
    .Y(_05750_));
 sky130_fd_sc_hd__inv_2 _12571_ (.A(net19),
    .Y(_05751_));
 sky130_fd_sc_hd__a211o_1 _12572_ (.A1(_05749_),
    .A2(net4068),
    .B1(net20),
    .C1(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__mux4_1 _12573_ (.A0(net4149),
    .A1(net4141),
    .A2(net4164),
    .A3(net7727),
    .S0(_05749_),
    .S1(net19),
    .X(_05753_));
 sky130_fd_sc_hd__a2bb2o_1 _12574_ (.A1_N(_05750_),
    .A2_N(_05752_),
    .B1(_05753_),
    .B2(net20),
    .X(_05754_));
 sky130_fd_sc_hd__a21o_1 _12575_ (.A1(_05747_),
    .A2(net18),
    .B1(net19),
    .X(_05755_));
 sky130_fd_sc_hd__and3_1 _12576_ (.A(net21),
    .B(net20),
    .C(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__mux4_1 _12577_ (.A0(net4111),
    .A1(_05673_),
    .A2(net4071),
    .A3(net4092),
    .S0(_05749_),
    .S1(net18),
    .X(_05757_));
 sky130_fd_sc_hd__mux4_1 _12578_ (.A0(net4103),
    .A1(net4024),
    .A2(_05730_),
    .A3(net3996),
    .S0(net16),
    .S1(net19),
    .X(_05758_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(net4128),
    .A1(_05043_),
    .S(net16),
    .X(_05759_));
 sky130_fd_sc_hd__inv_2 _12580_ (.A(net18),
    .Y(_05760_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(_05758_),
    .A1(_05759_),
    .S(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__mux2_1 _12582_ (.A0(_05757_),
    .A1(_05761_),
    .S(_05747_),
    .X(_05762_));
 sky130_fd_sc_hd__and2b_1 _12583_ (.A_N(net17),
    .B(net16),
    .X(_05763_));
 sky130_fd_sc_hd__and2b_1 _12584_ (.A_N(net16),
    .B(_05747_),
    .X(_05764_));
 sky130_fd_sc_hd__and3_1 _12585_ (.A(net50),
    .B(_05747_),
    .C(_05749_),
    .X(_05765_));
 sky130_fd_sc_hd__a211o_1 _12586_ (.A1(net49),
    .A2(_05764_),
    .B1(_05765_),
    .C1(_05760_),
    .X(_05766_));
 sky130_fd_sc_hd__a221o_1 _12587_ (.A1(net4066),
    .A2(_05744_),
    .B1(_05763_),
    .B2(net71),
    .C1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__mux4_1 _12588_ (.A0(net51),
    .A1(net41),
    .A2(net40),
    .A3(_05203_),
    .S0(_05747_),
    .S1(_05749_),
    .X(_05768_));
 sky130_fd_sc_hd__a21bo_1 _12589_ (.A1(_05760_),
    .A2(_05768_),
    .B1_N(net19),
    .X(_05769_));
 sky130_fd_sc_hd__a21bo_1 _12590_ (.A1(net46),
    .A2(_05763_),
    .B1_N(_05745_),
    .X(_05770_));
 sky130_fd_sc_hd__a221o_1 _12591_ (.A1(net43),
    .A2(_05744_),
    .B1(_05764_),
    .B2(net44),
    .C1(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__a31o_1 _12592_ (.A1(_05747_),
    .A2(_05749_),
    .A3(net4147),
    .B1(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__and4b_1 _12593_ (.A_N(net20),
    .B(_05769_),
    .C(_05772_),
    .D(net21),
    .X(_05773_));
 sky130_fd_sc_hd__a22oi_1 _12594_ (.A1(_05756_),
    .A2(_05762_),
    .B1(_05767_),
    .B2(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__mux4_1 _12595_ (.A0(_04648_),
    .A1(_04461_),
    .A2(_04468_),
    .A3(_04023_),
    .S0(_05749_),
    .S1(_05747_),
    .X(_05775_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(net4133),
    .A1(net4089),
    .S(_05749_),
    .X(_05776_));
 sky130_fd_sc_hd__mux4_1 _12597_ (.A0(_04020_),
    .A1(_04495_),
    .A2(net7678),
    .A3(_04500_),
    .S0(net16),
    .S1(_05747_),
    .X(_05777_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(_05776_),
    .A1(_05777_),
    .S(net19),
    .X(_05778_));
 sky130_fd_sc_hd__nand2_1 _12599_ (.A(net20),
    .B(_05755_),
    .Y(_05779_));
 sky130_fd_sc_hd__a21o_1 _12600_ (.A1(net19),
    .A2(net18),
    .B1(net20),
    .X(_05780_));
 sky130_fd_sc_hd__o2111a_1 _12601_ (.A1(_05760_),
    .A2(_05778_),
    .B1(_05779_),
    .C1(_05780_),
    .D1(net21),
    .X(_05781_));
 sky130_fd_sc_hd__o21ai_1 _12602_ (.A1(net18),
    .A2(_05775_),
    .B1(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__nor2_1 _12603_ (.A(net19),
    .B(_05760_),
    .Y(_05783_));
 sky130_fd_sc_hd__a22o_1 _12604_ (.A1(net52),
    .A2(_05744_),
    .B1(_05763_),
    .B2(net53),
    .X(_05784_));
 sky130_fd_sc_hd__a21o_1 _12605_ (.A1(net55),
    .A2(_05764_),
    .B1(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__a22o_2 _12606_ (.A1(net47),
    .A2(_05763_),
    .B1(_05764_),
    .B2(clknet_leaf_89_i_clk),
    .X(_05786_));
 sky130_fd_sc_hd__a22o_1 _12607_ (.A1(net6041),
    .A2(_05745_),
    .B1(_05783_),
    .B2(net54),
    .X(_05787_));
 sky130_fd_sc_hd__inv_2 _12608_ (.A(_05746_),
    .Y(_05788_));
 sky130_fd_sc_hd__a31o_1 _12609_ (.A1(_05747_),
    .A2(_05749_),
    .A3(_05787_),
    .B1(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__a221o_2 _12610_ (.A1(_05783_),
    .A2(_05785_),
    .B1(_05786_),
    .B2(_05745_),
    .C1(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__or3b_2 _12611_ (.A(net21),
    .B(net20),
    .C_N(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__nand3_2 _12612_ (.A(_05774_),
    .B(_05782_),
    .C(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__a41o_2 _12613_ (.A1(_05747_),
    .A2(net18),
    .A3(_05748_),
    .A4(_05754_),
    .B1(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__o41a_2 _12614_ (.A1(net21),
    .A2(net20),
    .A3(net4156),
    .A4(_05746_),
    .B1(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__mux2_2 _12615_ (.A0(\reg_gpout[2] ),
    .A1(clknet_1_1__leaf__05794_),
    .S(net45),
    .X(_05795_));
 sky130_fd_sc_hd__buf_1 _12616_ (.A(_05795_),
    .X(net58));
 sky130_fd_sc_hd__nor2_1 _12617_ (.A(net27),
    .B(net26),
    .Y(_05796_));
 sky130_fd_sc_hd__clkbuf_4 _12618_ (.A(net23),
    .X(_05797_));
 sky130_fd_sc_hd__nor2_1 _12619_ (.A(_05797_),
    .B(net22),
    .Y(_05798_));
 sky130_fd_sc_hd__nor2_1 _12620_ (.A(net25),
    .B(net24),
    .Y(_05799_));
 sky130_fd_sc_hd__and3_1 _12621_ (.A(_05796_),
    .B(_05798_),
    .C(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__inv_2 _12622_ (.A(net27),
    .Y(_05801_));
 sky130_fd_sc_hd__clkbuf_4 _12623_ (.A(net22),
    .X(_05802_));
 sky130_fd_sc_hd__nor2_1 _12624_ (.A(_05802_),
    .B(net4156),
    .Y(_05803_));
 sky130_fd_sc_hd__inv_2 _12625_ (.A(net25),
    .Y(_05804_));
 sky130_fd_sc_hd__a211o_1 _12626_ (.A1(_05802_),
    .A2(net7571),
    .B1(net26),
    .C1(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__mux4_1 _12627_ (.A0(net4149),
    .A1(net4141),
    .A2(net4164),
    .A3(net7727),
    .S0(_05802_),
    .S1(net25),
    .X(_05806_));
 sky130_fd_sc_hd__a2bb2o_1 _12628_ (.A1_N(_05803_),
    .A2_N(_05805_),
    .B1(_05806_),
    .B2(net26),
    .X(_05807_));
 sky130_fd_sc_hd__nand4_1 _12629_ (.A(_05797_),
    .B(net24),
    .C(_05801_),
    .D(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__a21o_1 _12630_ (.A1(_05797_),
    .A2(net24),
    .B1(net25),
    .X(_05809_));
 sky130_fd_sc_hd__and3_1 _12631_ (.A(net27),
    .B(net26),
    .C(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__mux4_1 _12632_ (.A0(net4111),
    .A1(_05673_),
    .A2(net4071),
    .A3(net4092),
    .S0(_05802_),
    .S1(net24),
    .X(_05811_));
 sky130_fd_sc_hd__mux4_1 _12633_ (.A0(net4103),
    .A1(net4024),
    .A2(_05730_),
    .A3(net3996),
    .S0(net22),
    .S1(net25),
    .X(_05812_));
 sky130_fd_sc_hd__mux2_1 _12634_ (.A0(net4128),
    .A1(_05043_),
    .S(net22),
    .X(_05813_));
 sky130_fd_sc_hd__inv_2 _12635_ (.A(net24),
    .Y(_05814_));
 sky130_fd_sc_hd__mux2_1 _12636_ (.A0(_05812_),
    .A1(_05813_),
    .S(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__mux2_1 _12637_ (.A0(_05811_),
    .A1(_05815_),
    .S(_05797_),
    .X(_05816_));
 sky130_fd_sc_hd__and2b_1 _12638_ (.A_N(net23),
    .B(net22),
    .X(_05817_));
 sky130_fd_sc_hd__and2b_1 _12639_ (.A_N(net22),
    .B(net23),
    .X(_05818_));
 sky130_fd_sc_hd__and3_1 _12640_ (.A(net50),
    .B(_05797_),
    .C(_05802_),
    .X(_05819_));
 sky130_fd_sc_hd__a211o_1 _12641_ (.A1(net49),
    .A2(_05818_),
    .B1(_05819_),
    .C1(_05814_),
    .X(_05820_));
 sky130_fd_sc_hd__a221o_1 _12642_ (.A1(net4066),
    .A2(_05798_),
    .B1(_05817_),
    .B2(net71),
    .C1(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__mux4_1 _12643_ (.A0(net51),
    .A1(net41),
    .A2(net40),
    .A3(_05203_),
    .S0(_05797_),
    .S1(_05802_),
    .X(_05822_));
 sky130_fd_sc_hd__nand2_1 _12644_ (.A(_05814_),
    .B(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__a21bo_1 _12645_ (.A1(net46),
    .A2(_05817_),
    .B1_N(_05799_),
    .X(_05824_));
 sky130_fd_sc_hd__a221o_1 _12646_ (.A1(net43),
    .A2(_05798_),
    .B1(_05818_),
    .B2(net44),
    .C1(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__a31oi_1 _12647_ (.A1(_05797_),
    .A2(_05802_),
    .A3(net4147),
    .B1(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__a2111oi_1 _12648_ (.A1(net25),
    .A2(_05823_),
    .B1(_05826_),
    .C1(_05801_),
    .D1(net26),
    .Y(_05827_));
 sky130_fd_sc_hd__a22o_1 _12649_ (.A1(_05810_),
    .A2(_05816_),
    .B1(_05821_),
    .B2(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__mux4_1 _12650_ (.A0(_04648_),
    .A1(_04461_),
    .A2(_04468_),
    .A3(_04023_),
    .S0(_05802_),
    .S1(_05797_),
    .X(_05829_));
 sky130_fd_sc_hd__or2_1 _12651_ (.A(net24),
    .B(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(net4133),
    .A1(net4089),
    .S(_05802_),
    .X(_05831_));
 sky130_fd_sc_hd__mux4_1 _12653_ (.A0(_04020_),
    .A1(_04495_),
    .A2(_04494_),
    .A3(_04500_),
    .S0(net22),
    .S1(_05797_),
    .X(_05832_));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(_05831_),
    .A1(_05832_),
    .S(net25),
    .X(_05833_));
 sky130_fd_sc_hd__nand2_1 _12655_ (.A(net26),
    .B(_05809_),
    .Y(_05834_));
 sky130_fd_sc_hd__a21o_1 _12656_ (.A1(net25),
    .A2(net24),
    .B1(net26),
    .X(_05835_));
 sky130_fd_sc_hd__o2111a_1 _12657_ (.A1(_05814_),
    .A2(_05833_),
    .B1(_05834_),
    .C1(_05835_),
    .D1(net27),
    .X(_05836_));
 sky130_fd_sc_hd__nor2_1 _12658_ (.A(net25),
    .B(_05814_),
    .Y(_05837_));
 sky130_fd_sc_hd__a22o_1 _12659_ (.A1(net52),
    .A2(_05798_),
    .B1(_05817_),
    .B2(net53),
    .X(_05838_));
 sky130_fd_sc_hd__a21o_1 _12660_ (.A1(net55),
    .A2(_05818_),
    .B1(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__a22o_2 _12661_ (.A1(net48),
    .A2(_05817_),
    .B1(_05818_),
    .B2(clknet_1_1__leaf__05645_),
    .X(_05840_));
 sky130_fd_sc_hd__a22o_1 _12662_ (.A1(net6627),
    .A2(_05799_),
    .B1(_05837_),
    .B2(net54),
    .X(_05841_));
 sky130_fd_sc_hd__and2_1 _12663_ (.A(_05798_),
    .B(_05799_),
    .X(_05842_));
 sky130_fd_sc_hd__a31o_1 _12664_ (.A1(_05797_),
    .A2(_05802_),
    .A3(_05841_),
    .B1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__a221o_2 _12665_ (.A1(_05837_),
    .A2(_05839_),
    .B1(_05840_),
    .B2(_05799_),
    .C1(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__a22o_2 _12666_ (.A1(_05830_),
    .A2(_05836_),
    .B1(_05844_),
    .B2(_05796_),
    .X(_05845_));
 sky130_fd_sc_hd__nor2_2 _12667_ (.A(_05828_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__a22oi_2 _12668_ (.A1(net7571),
    .A2(_05800_),
    .B1(_05808_),
    .B2(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__mux2_2 _12669_ (.A0(\reg_gpout[3] ),
    .A1(clknet_1_1__leaf__05847_),
    .S(net45),
    .X(_05848_));
 sky130_fd_sc_hd__buf_1 _12670_ (.A(_05848_),
    .X(net59));
 sky130_fd_sc_hd__nor2_1 _12671_ (.A(net32),
    .B(net33),
    .Y(_05849_));
 sky130_fd_sc_hd__buf_2 _12672_ (.A(net29),
    .X(_05850_));
 sky130_fd_sc_hd__clkbuf_4 _12673_ (.A(net28),
    .X(_05851_));
 sky130_fd_sc_hd__nor2_1 _12674_ (.A(_05850_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__nor2_1 _12675_ (.A(net31),
    .B(net30),
    .Y(_05853_));
 sky130_fd_sc_hd__and2_1 _12676_ (.A(_05852_),
    .B(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__nand2_1 _12677_ (.A(_05849_),
    .B(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__nor2_1 _12678_ (.A(_05851_),
    .B(net4156),
    .Y(_05856_));
 sky130_fd_sc_hd__inv_2 _12679_ (.A(net31),
    .Y(_05857_));
 sky130_fd_sc_hd__a211o_1 _12680_ (.A1(_05851_),
    .A2(net4068),
    .B1(net32),
    .C1(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__mux4_1 _12681_ (.A0(net4149),
    .A1(net4141),
    .A2(net4164),
    .A3(net7727),
    .S0(_05851_),
    .S1(net31),
    .X(_05859_));
 sky130_fd_sc_hd__a2bb2o_1 _12682_ (.A1_N(_05856_),
    .A2_N(_05858_),
    .B1(_05859_),
    .B2(net32),
    .X(_05860_));
 sky130_fd_sc_hd__and4b_1 _12683_ (.A_N(net33),
    .B(_05860_),
    .C(_05850_),
    .D(net30),
    .X(_05861_));
 sky130_fd_sc_hd__inv_2 _12684_ (.A(net30),
    .Y(_05862_));
 sky130_fd_sc_hd__nor2_1 _12685_ (.A(net31),
    .B(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__and2b_1 _12686_ (.A_N(net28),
    .B(net29),
    .X(_05864_));
 sky130_fd_sc_hd__and2b_1 _12687_ (.A_N(net29),
    .B(net28),
    .X(_05865_));
 sky130_fd_sc_hd__a22o_1 _12688_ (.A1(net52),
    .A2(_05852_),
    .B1(_05865_),
    .B2(net53),
    .X(_05866_));
 sky130_fd_sc_hd__a21o_1 _12689_ (.A1(net55),
    .A2(_05864_),
    .B1(_05866_),
    .X(_05867_));
 sky130_fd_sc_hd__a22o_2 _12690_ (.A1(net3),
    .A2(_05865_),
    .B1(_05864_),
    .B2(clknet_1_1__leaf__05645_),
    .X(_05868_));
 sky130_fd_sc_hd__a22o_1 _12691_ (.A1(net6111),
    .A2(_05853_),
    .B1(_05863_),
    .B2(net54),
    .X(_05869_));
 sky130_fd_sc_hd__a31o_1 _12692_ (.A1(_05850_),
    .A2(_05851_),
    .A3(_05869_),
    .B1(_05854_),
    .X(_05870_));
 sky130_fd_sc_hd__a221o_2 _12693_ (.A1(_05863_),
    .A2(_05867_),
    .B1(_05868_),
    .B2(_05853_),
    .C1(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__mux4_1 _12694_ (.A0(_04648_),
    .A1(_04461_),
    .A2(_04468_),
    .A3(_04023_),
    .S0(_05851_),
    .S1(_05850_),
    .X(_05872_));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(net4133),
    .A1(net4089),
    .S(_05851_),
    .X(_05873_));
 sky130_fd_sc_hd__mux4_1 _12696_ (.A0(_04020_),
    .A1(_04495_),
    .A2(net7678),
    .A3(_04500_),
    .S0(net28),
    .S1(_05850_),
    .X(_05874_));
 sky130_fd_sc_hd__mux2_1 _12697_ (.A0(_05873_),
    .A1(_05874_),
    .S(net31),
    .X(_05875_));
 sky130_fd_sc_hd__a21o_1 _12698_ (.A1(_05850_),
    .A2(net30),
    .B1(net31),
    .X(_05876_));
 sky130_fd_sc_hd__nand2_1 _12699_ (.A(net32),
    .B(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__a21o_1 _12700_ (.A1(net31),
    .A2(net30),
    .B1(net32),
    .X(_05878_));
 sky130_fd_sc_hd__o2111a_1 _12701_ (.A1(_05862_),
    .A2(_05875_),
    .B1(_05877_),
    .C1(_05878_),
    .D1(net33),
    .X(_05879_));
 sky130_fd_sc_hd__o21a_1 _12702_ (.A1(net30),
    .A2(_05872_),
    .B1(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__and3_1 _12703_ (.A(net50),
    .B(_05850_),
    .C(_05851_),
    .X(_05881_));
 sky130_fd_sc_hd__a211o_1 _12704_ (.A1(net49),
    .A2(_05864_),
    .B1(_05881_),
    .C1(_05862_),
    .X(_05882_));
 sky130_fd_sc_hd__a221o_1 _12705_ (.A1(net4066),
    .A2(_05852_),
    .B1(_05865_),
    .B2(net71),
    .C1(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__mux4_1 _12706_ (.A0(net51),
    .A1(net41),
    .A2(net40),
    .A3(_05203_),
    .S0(_05850_),
    .S1(_05851_),
    .X(_05884_));
 sky130_fd_sc_hd__a21bo_1 _12707_ (.A1(_05862_),
    .A2(_05884_),
    .B1_N(net31),
    .X(_05885_));
 sky130_fd_sc_hd__a21bo_1 _12708_ (.A1(net46),
    .A2(_05865_),
    .B1_N(_05853_),
    .X(_05886_));
 sky130_fd_sc_hd__a221o_1 _12709_ (.A1(net43),
    .A2(_05852_),
    .B1(_05864_),
    .B2(net44),
    .C1(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__a31o_1 _12710_ (.A1(_05850_),
    .A2(_05851_),
    .A3(net4147),
    .B1(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__and3b_1 _12711_ (.A_N(net32),
    .B(net33),
    .C(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__mux4_1 _12712_ (.A0(net4111),
    .A1(_05673_),
    .A2(net4071),
    .A3(net4092),
    .S0(net28),
    .S1(net30),
    .X(_05890_));
 sky130_fd_sc_hd__mux4_1 _12713_ (.A0(net4102),
    .A1(net4024),
    .A2(net5965),
    .A3(net6044),
    .S0(net28),
    .S1(net31),
    .X(_05891_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(net4128),
    .A1(_05043_),
    .S(net28),
    .X(_05892_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(_05891_),
    .A1(_05892_),
    .S(_05862_),
    .X(_05893_));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(_05890_),
    .A1(_05893_),
    .S(_05850_),
    .X(_05894_));
 sky130_fd_sc_hd__and4_1 _12717_ (.A(net32),
    .B(net33),
    .C(_05876_),
    .D(_05894_),
    .X(_05895_));
 sky130_fd_sc_hd__a31o_1 _12718_ (.A1(_05883_),
    .A2(_05885_),
    .A3(_05889_),
    .B1(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__a211o_2 _12719_ (.A1(_05849_),
    .A2(_05871_),
    .B1(_05880_),
    .C1(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__o22a_2 _12720_ (.A1(net4164),
    .A2(_05855_),
    .B1(_05861_),
    .B2(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__mux2_2 _12721_ (.A0(\reg_gpout[4] ),
    .A1(clknet_1_1__leaf__05898_),
    .S(net45),
    .X(_05899_));
 sky130_fd_sc_hd__buf_1 _12722_ (.A(_05899_),
    .X(net60));
 sky130_fd_sc_hd__or2_1 _12723_ (.A(net38),
    .B(net39),
    .X(_05900_));
 sky130_fd_sc_hd__clkbuf_4 _12724_ (.A(net34),
    .X(_05901_));
 sky130_fd_sc_hd__nor2_2 _12725_ (.A(net35),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__or4b_1 _12726_ (.A(net37),
    .B(net36),
    .C(_05900_),
    .D_N(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__inv_2 _12727_ (.A(net35),
    .Y(_05904_));
 sky130_fd_sc_hd__inv_2 _12728_ (.A(net36),
    .Y(_05905_));
 sky130_fd_sc_hd__and2b_1 _12729_ (.A_N(net38),
    .B(net37),
    .X(_05906_));
 sky130_fd_sc_hd__or2_1 _12730_ (.A(_05901_),
    .B(net4156),
    .X(_05907_));
 sky130_fd_sc_hd__nand2_1 _12731_ (.A(_05901_),
    .B(net4068),
    .Y(_05908_));
 sky130_fd_sc_hd__mux4_1 _12732_ (.A0(net4149),
    .A1(net4141),
    .A2(net4164),
    .A3(net4173),
    .S0(_05901_),
    .S1(net37),
    .X(_05909_));
 sky130_fd_sc_hd__a32o_1 _12733_ (.A1(_05906_),
    .A2(_05907_),
    .A3(_05908_),
    .B1(_05909_),
    .B2(net38),
    .X(_05910_));
 sky130_fd_sc_hd__or3b_1 _12734_ (.A(_05904_),
    .B(_05905_),
    .C_N(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__and2_2 _12735_ (.A(net35),
    .B(net34),
    .X(_05912_));
 sky130_fd_sc_hd__a21oi_2 _12736_ (.A1(net144),
    .A2(net35),
    .B1(_05901_),
    .Y(_05913_));
 sky130_fd_sc_hd__a21oi_2 _12737_ (.A1(net6058),
    .A2(_05912_),
    .B1(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__and2_1 _12738_ (.A(_05904_),
    .B(net34),
    .X(_05915_));
 sky130_fd_sc_hd__nor2_1 _12739_ (.A(_05904_),
    .B(net34),
    .Y(_05916_));
 sky130_fd_sc_hd__a22o_1 _12740_ (.A1(net52),
    .A2(_05902_),
    .B1(_05916_),
    .B2(net55),
    .X(_05917_));
 sky130_fd_sc_hd__a221o_1 _12741_ (.A1(net54),
    .A2(_05912_),
    .B1(_05915_),
    .B2(net53),
    .C1(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__or3b_1 _12742_ (.A(net37),
    .B(_05905_),
    .C_N(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__o31a_2 _12743_ (.A1(net37),
    .A2(net36),
    .A3(_05914_),
    .B1(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__mux4_1 _12744_ (.A0(_04648_),
    .A1(net4133),
    .A2(_04461_),
    .A3(net4089),
    .S0(net36),
    .S1(_05901_),
    .X(_05921_));
 sky130_fd_sc_hd__mux2_1 _12745_ (.A0(_04468_),
    .A1(_04023_),
    .S(_05901_),
    .X(_05922_));
 sky130_fd_sc_hd__mux2_1 _12746_ (.A0(net4103),
    .A1(net4024),
    .S(net34),
    .X(_05923_));
 sky130_fd_sc_hd__and3_1 _12747_ (.A(net35),
    .B(net36),
    .C(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__a31o_1 _12748_ (.A1(net35),
    .A2(_05905_),
    .A3(_05922_),
    .B1(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__a21oi_1 _12749_ (.A1(_05904_),
    .A2(_05921_),
    .B1(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__mux4_1 _12750_ (.A0(net4111),
    .A1(_05673_),
    .A2(net4071),
    .A3(net4092),
    .S0(_05901_),
    .S1(net36),
    .X(_05927_));
 sky130_fd_sc_hd__mux4_1 _12751_ (.A0(_05680_),
    .A1(_05043_),
    .A2(_05730_),
    .A3(net3996),
    .S0(_05901_),
    .S1(net36),
    .X(_05928_));
 sky130_fd_sc_hd__o21a_1 _12752_ (.A1(_05904_),
    .A2(_05928_),
    .B1(net37),
    .X(_05929_));
 sky130_fd_sc_hd__o21ai_1 _12753_ (.A1(net35),
    .A2(_05927_),
    .B1(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__o21ai_1 _12754_ (.A1(net37),
    .A2(_05926_),
    .B1(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__mux4_1 _12755_ (.A0(_04020_),
    .A1(_04495_),
    .A2(_04494_),
    .A3(_04500_),
    .S0(_05901_),
    .S1(net35),
    .X(_05932_));
 sky130_fd_sc_hd__a221o_1 _12756_ (.A1(_05203_),
    .A2(_05912_),
    .B1(_05916_),
    .B2(net41),
    .C1(net36),
    .X(_05933_));
 sky130_fd_sc_hd__o211a_1 _12757_ (.A1(_05905_),
    .A2(_05932_),
    .B1(_05933_),
    .C1(_05906_),
    .X(_05934_));
 sky130_fd_sc_hd__a211o_1 _12758_ (.A1(net43),
    .A2(_05902_),
    .B1(net36),
    .C1(net37),
    .X(_05935_));
 sky130_fd_sc_hd__a22o_1 _12759_ (.A1(net44),
    .A2(_05916_),
    .B1(_05915_),
    .B2(net46),
    .X(_05936_));
 sky130_fd_sc_hd__a211o_1 _12760_ (.A1(net4147),
    .A2(_05912_),
    .B1(_05935_),
    .C1(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__a221o_1 _12761_ (.A1(net50),
    .A2(_05912_),
    .B1(_05916_),
    .B2(net49),
    .C1(_05905_),
    .X(_05938_));
 sky130_fd_sc_hd__a221o_1 _12762_ (.A1(net4066),
    .A2(_05902_),
    .B1(_05915_),
    .B2(net71),
    .C1(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__a22o_1 _12763_ (.A1(net51),
    .A2(_05902_),
    .B1(_05915_),
    .B2(net40),
    .X(_05940_));
 sky130_fd_sc_hd__a21bo_1 _12764_ (.A1(_05905_),
    .A2(_05940_),
    .B1_N(net37),
    .X(_05941_));
 sky130_fd_sc_hd__and4b_1 _12765_ (.A_N(net38),
    .B(_05937_),
    .C(_05939_),
    .D(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__a211o_1 _12766_ (.A1(net38),
    .A2(_05931_),
    .B1(_05934_),
    .C1(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__nand2_1 _12767_ (.A(net39),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__o221a_2 _12768_ (.A1(net39),
    .A2(_05911_),
    .B1(_05920_),
    .B2(_05900_),
    .C1(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__o21ba_2 _12769_ (.A1(net7727),
    .A2(_05903_),
    .B1_N(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__mux2_2 _12770_ (.A0(\reg_gpout[5] ),
    .A1(clknet_1_1__leaf__05946_),
    .S(net45),
    .X(_05947_));
 sky130_fd_sc_hd__buf_1 _12771_ (.A(_05947_),
    .X(net61));
 sky130_fd_sc_hd__nand2_2 _12772_ (.A(net4416),
    .B(net3761),
    .Y(_05948_));
 sky130_fd_sc_hd__nor2_2 _12773_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_05949_));
 sky130_fd_sc_hd__and2_2 _12774_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_05950_));
 sky130_fd_sc_hd__nor2_1 _12775_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_05951_));
 sky130_fd_sc_hd__nor2_4 _12776_ (.A(_05950_),
    .B(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__xor2_4 _12777_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_05953_));
 sky130_fd_sc_hd__and2_1 _12778_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_05954_));
 sky130_fd_sc_hd__a31o_4 _12779_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_05953_),
    .B1(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__a221oi_4 _12780_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_05952_),
    .B2(_05955_),
    .C1(_05950_),
    .Y(_05956_));
 sky130_fd_sc_hd__nand2_1 _12781_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_05957_));
 sky130_fd_sc_hd__or2_1 _12782_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_05958_));
 sky130_fd_sc_hd__and2_1 _12783_ (.A(_05957_),
    .B(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__inv_2 _12784_ (.A(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__nand2_1 _12785_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_05961_));
 sky130_fd_sc_hd__or2_1 _12786_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_05962_));
 sky130_fd_sc_hd__xor2_1 _12787_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_05963_));
 sky130_fd_sc_hd__nand3_1 _12788_ (.A(_05961_),
    .B(_05962_),
    .C(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__nor2_1 _12789_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_05965_));
 sky130_fd_sc_hd__nand2_1 _12790_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_05966_));
 sky130_fd_sc_hd__or2b_2 _12791_ (.A(_05965_),
    .B_N(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__or2_1 _12792_ (.A(_05964_),
    .B(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__or4_4 _12793_ (.A(_05949_),
    .B(_05956_),
    .C(_05960_),
    .D(_05968_),
    .X(_05969_));
 sky130_fd_sc_hd__a21o_1 _12794_ (.A1(_05957_),
    .A2(_05966_),
    .B1(_05965_),
    .X(_05970_));
 sky130_fd_sc_hd__nand2_1 _12795_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_05971_));
 sky130_fd_sc_hd__or2b_1 _12796_ (.A(_05971_),
    .B_N(_05962_),
    .X(_05972_));
 sky130_fd_sc_hd__o211a_1 _12797_ (.A1(_05964_),
    .A2(_05970_),
    .B1(_05972_),
    .C1(_05961_),
    .X(_05973_));
 sky130_fd_sc_hd__or2_1 _12798_ (.A(net4416),
    .B(net3761),
    .X(_05974_));
 sky130_fd_sc_hd__nand2_1 _12799_ (.A(_05948_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__a21o_4 _12800_ (.A1(_05969_),
    .A2(_05973_),
    .B1(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__nand2_2 _12801_ (.A(net7744),
    .B(net6046),
    .Y(_05977_));
 sky130_fd_sc_hd__nor2_2 _12802_ (.A(net7744),
    .B(net6046),
    .Y(_05978_));
 sky130_fd_sc_hd__nor2_1 _12803_ (.A(net7746),
    .B(net4838),
    .Y(_05979_));
 sky130_fd_sc_hd__a311o_4 _12804_ (.A1(_05948_),
    .A2(_05976_),
    .A3(_05977_),
    .B1(_05978_),
    .C1(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__nor2_1 _12805_ (.A(net7746),
    .B(net5955),
    .Y(_05981_));
 sky130_fd_sc_hd__nand2_1 _12806_ (.A(net7746),
    .B(net4838),
    .Y(_05982_));
 sky130_fd_sc_hd__and2b_1 _12807_ (.A_N(_05981_),
    .B(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__and2_1 _12808_ (.A(net7746),
    .B(net5955),
    .X(_05984_));
 sky130_fd_sc_hd__a21oi_2 _12809_ (.A1(_05980_),
    .A2(_05983_),
    .B1(_05984_),
    .Y(_05985_));
 sky130_fd_sc_hd__or2_1 _12810_ (.A(_05984_),
    .B(_05981_),
    .X(_05986_));
 sky130_fd_sc_hd__a21bo_1 _12811_ (.A1(_05980_),
    .A2(_05982_),
    .B1_N(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__nand3b_1 _12812_ (.A_N(_05986_),
    .B(_05982_),
    .C(_05980_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand2_1 _12813_ (.A(_05987_),
    .B(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__and2b_1 _12814_ (.A_N(_05979_),
    .B(_05982_),
    .X(_05990_));
 sky130_fd_sc_hd__inv_2 _12815_ (.A(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__a311oi_4 _12816_ (.A1(_05948_),
    .A2(_05976_),
    .A3(_05977_),
    .B1(_05991_),
    .C1(_05978_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand3b_1 _12817_ (.A_N(_05978_),
    .B(net3761),
    .C(net4416),
    .Y(_05993_));
 sky130_fd_sc_hd__o2111a_1 _12818_ (.A1(_05978_),
    .A2(_05976_),
    .B1(_05977_),
    .C1(_05993_),
    .D1(_05991_),
    .X(_05994_));
 sky130_fd_sc_hd__nor2_1 _12819_ (.A(_05992_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__o41a_1 _12820_ (.A1(_05949_),
    .A2(_05956_),
    .A3(_05960_),
    .A4(_05967_),
    .B1(_05970_),
    .X(_05996_));
 sky130_fd_sc_hd__xnor2_1 _12821_ (.A(_05963_),
    .B(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__nand3_1 _12822_ (.A(_05975_),
    .B(_05969_),
    .C(_05973_),
    .Y(_05998_));
 sky130_fd_sc_hd__and2_1 _12823_ (.A(_05976_),
    .B(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__or3_4 _12824_ (.A(_05949_),
    .B(_05956_),
    .C(_05960_),
    .X(_06000_));
 sky130_fd_sc_hd__o21ai_1 _12825_ (.A1(_05949_),
    .A2(_05956_),
    .B1(_05960_),
    .Y(_06001_));
 sky130_fd_sc_hd__and2_1 _12826_ (.A(_06000_),
    .B(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__nand2_1 _12827_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_06003_));
 sky130_fd_sc_hd__or2b_1 _12828_ (.A(_05949_),
    .B_N(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__a21o_1 _12829_ (.A1(_05952_),
    .A2(_05955_),
    .B1(_05950_),
    .X(_06005_));
 sky130_fd_sc_hd__xnor2_2 _12830_ (.A(_06004_),
    .B(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__xor2_2 _12831_ (.A(_05952_),
    .B(_05955_),
    .X(_06007_));
 sky130_fd_sc_hd__nand2_1 _12832_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_06008_));
 sky130_fd_sc_hd__xnor2_2 _12833_ (.A(_06008_),
    .B(_05953_),
    .Y(_06009_));
 sky130_fd_sc_hd__xor2_1 _12834_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_06010_));
 sky130_fd_sc_hd__or4_1 _12835_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C(_06009_),
    .D(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__or2_1 _12836_ (.A(_06007_),
    .B(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__or4_1 _12837_ (.A(_05999_),
    .B(_06002_),
    .C(_06006_),
    .D(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__o31a_1 _12838_ (.A1(_05949_),
    .A2(_05956_),
    .A3(_05960_),
    .B1(_05957_),
    .X(_06014_));
 sky130_fd_sc_hd__xnor2_2 _12839_ (.A(_05967_),
    .B(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__inv_2 _12840_ (.A(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__or2b_1 _12841_ (.A(_05978_),
    .B_N(_05977_),
    .X(_06017_));
 sky130_fd_sc_hd__a21oi_1 _12842_ (.A1(_05948_),
    .A2(_05976_),
    .B1(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__and3_1 _12843_ (.A(_05948_),
    .B(_05976_),
    .C(_06017_),
    .X(_06019_));
 sky130_fd_sc_hd__or2_1 _12844_ (.A(_06018_),
    .B(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__or4b_1 _12845_ (.A(_05997_),
    .B(_06013_),
    .C(_06016_),
    .D_N(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__nand2_1 _12846_ (.A(_05961_),
    .B(_05962_),
    .Y(_06022_));
 sky130_fd_sc_hd__nor2_1 _12847_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06023_));
 sky130_fd_sc_hd__o21a_1 _12848_ (.A1(_06023_),
    .A2(_05996_),
    .B1(_05971_),
    .X(_06024_));
 sky130_fd_sc_hd__xnor2_2 _12849_ (.A(_06022_),
    .B(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__or4b_1 _12850_ (.A(_05989_),
    .B(_05995_),
    .C(_06021_),
    .D_N(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__nand2_4 _12851_ (.A(_05985_),
    .B(net7775),
    .Y(_06027_));
 sky130_fd_sc_hd__clkbuf_4 _12852_ (.A(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__xor2_1 _12853_ (.A(net5605),
    .B(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__inv_2 _12854_ (.A(net7575),
    .Y(_06030_));
 sky130_fd_sc_hd__xnor2_2 _12855_ (.A(_06030_),
    .B(_06028_),
    .Y(_06031_));
 sky130_fd_sc_hd__inv_2 _12856_ (.A(net4043),
    .Y(_06032_));
 sky130_fd_sc_hd__inv_2 _12857_ (.A(net7776),
    .Y(_06033_));
 sky130_fd_sc_hd__nor2_1 _12858_ (.A(_06032_),
    .B(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__buf_1 _12859_ (.A(net4043),
    .X(_06035_));
 sky130_fd_sc_hd__or2_1 _12860_ (.A(net4044),
    .B(_06028_),
    .X(_06036_));
 sky130_fd_sc_hd__inv_2 _12861_ (.A(net4641),
    .Y(_06037_));
 sky130_fd_sc_hd__nor2_1 _12862_ (.A(net4642),
    .B(_06033_),
    .Y(_06038_));
 sky130_fd_sc_hd__buf_2 _12863_ (.A(net5937),
    .X(_06039_));
 sky130_fd_sc_hd__nor2_1 _12864_ (.A(_06039_),
    .B(_06028_),
    .Y(_06040_));
 sky130_fd_sc_hd__nor2_1 _12865_ (.A(_06038_),
    .B(_06040_),
    .Y(_06041_));
 sky130_fd_sc_hd__and2_1 _12866_ (.A(net3893),
    .B(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__inv_2 _12867_ (.A(net3848),
    .Y(_06043_));
 sky130_fd_sc_hd__xnor2_1 _12868_ (.A(_06043_),
    .B(_06028_),
    .Y(_06044_));
 sky130_fd_sc_hd__o21a_1 _12869_ (.A1(_06038_),
    .A2(_06042_),
    .B1(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__a21o_1 _12870_ (.A1(net3848),
    .A2(_06028_),
    .B1(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__and2_1 _12871_ (.A(_06036_),
    .B(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__inv_2 _12872_ (.A(net3807),
    .Y(_06048_));
 sky130_fd_sc_hd__xnor2_1 _12873_ (.A(_06048_),
    .B(_06028_),
    .Y(_06049_));
 sky130_fd_sc_hd__o21a_1 _12874_ (.A1(_06034_),
    .A2(_06047_),
    .B1(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__o21a_1 _12875_ (.A1(net3807),
    .A2(net3447),
    .B1(_06028_),
    .X(_06051_));
 sky130_fd_sc_hd__a21o_1 _12876_ (.A1(_06031_),
    .A2(_06050_),
    .B1(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__or2_1 _12877_ (.A(_06029_),
    .B(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__nand2_1 _12878_ (.A(_06029_),
    .B(_06052_),
    .Y(_06054_));
 sky130_fd_sc_hd__or3b_1 _12879_ (.A(net3975),
    .B(_04476_),
    .C_N(net3871),
    .X(_06055_));
 sky130_fd_sc_hd__buf_1 _12880_ (.A(net4864),
    .X(_06056_));
 sky130_fd_sc_hd__buf_8 _12881_ (.A(net4865),
    .X(_06057_));
 sky130_fd_sc_hd__buf_4 _12882_ (.A(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__inv_2 _12883_ (.A(net3682),
    .Y(_06059_));
 sky130_fd_sc_hd__buf_2 _12884_ (.A(net4048),
    .X(_06060_));
 sky130_fd_sc_hd__inv_2 _12885_ (.A(net5974),
    .Y(_06061_));
 sky130_fd_sc_hd__inv_2 _12886_ (.A(net3964),
    .Y(_06062_));
 sky130_fd_sc_hd__a2bb2o_1 _12887_ (.A1_N(net3326),
    .A2_N(_06061_),
    .B1(_06062_),
    .B2(net3389),
    .X(_06063_));
 sky130_fd_sc_hd__inv_2 _12888_ (.A(net4048),
    .Y(_06064_));
 sky130_fd_sc_hd__a22o_1 _12889_ (.A1(_04686_),
    .A2(net3964),
    .B1(_06030_),
    .B2(net3469),
    .X(_06065_));
 sky130_fd_sc_hd__a221o_1 _12890_ (.A1(net3682),
    .A2(net4007),
    .B1(_06043_),
    .B2(net4436),
    .C1(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__inv_2 _12891_ (.A(net4748),
    .Y(_06067_));
 sky130_fd_sc_hd__inv_2 _12892_ (.A(net7712),
    .Y(_06068_));
 sky130_fd_sc_hd__a2bb2o_1 _12893_ (.A1_N(net3469),
    .A2_N(_06030_),
    .B1(_06068_),
    .B2(net3990),
    .X(_06069_));
 sky130_fd_sc_hd__a221o_1 _12894_ (.A1(net4053),
    .A2(net4641),
    .B1(_06048_),
    .B2(net3552),
    .C1(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__clkbuf_1 _12895_ (.A(net4033),
    .X(_06071_));
 sky130_fd_sc_hd__a2bb2o_1 _12896_ (.A1_N(net4436),
    .A2_N(_06043_),
    .B1(net4044),
    .B2(_04674_),
    .X(_06072_));
 sky130_fd_sc_hd__a221o_1 _12897_ (.A1(net3991),
    .A2(net4034),
    .B1(net3807),
    .B2(net3553),
    .C1(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__or3_1 _12898_ (.A(_06066_),
    .B(_06070_),
    .C(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__a211o_1 _12899_ (.A1(net3683),
    .A2(net4049),
    .B1(_06063_),
    .C1(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__nand2_1 _12900_ (.A(net3431),
    .B(net3998),
    .Y(_06076_));
 sky130_fd_sc_hd__or2_1 _12901_ (.A(net3431),
    .B(net3998),
    .X(_06077_));
 sky130_fd_sc_hd__or4_1 _12902_ (.A(net2277),
    .B(net2058),
    .C(net1006),
    .D(net894),
    .X(_06078_));
 sky130_fd_sc_hd__or4_1 _12903_ (.A(net2968),
    .B(net1161),
    .C(net832),
    .D(net1611),
    .X(_06079_));
 sky130_fd_sc_hd__a211o_1 _12904_ (.A1(_06076_),
    .A2(_06077_),
    .B1(_06078_),
    .C1(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__inv_2 _12905_ (.A(net3959),
    .Y(_06081_));
 sky130_fd_sc_hd__a22o_1 _12906_ (.A1(net3326),
    .A2(_06061_),
    .B1(_06032_),
    .B2(net3473),
    .X(_06082_));
 sky130_fd_sc_hd__a221o_1 _12907_ (.A1(net3443),
    .A2(net3960),
    .B1(net4642),
    .B2(net4748),
    .C1(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__inv_2 _12908_ (.A(net4019),
    .Y(_06084_));
 sky130_fd_sc_hd__a211o_1 _12909_ (.A1(_06084_),
    .A2(net3884),
    .B1(net2379),
    .C1(net2006),
    .X(_06085_));
 sky130_fd_sc_hd__o22a_1 _12910_ (.A1(net3443),
    .A2(net3960),
    .B1(net3884),
    .B2(_06084_),
    .X(_06086_));
 sky130_fd_sc_hd__or4b_1 _12911_ (.A(_06080_),
    .B(_06083_),
    .C(_06085_),
    .D_N(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__or4_1 _12912_ (.A(net4705),
    .B(net4718),
    .C(net4751),
    .D(net4757),
    .X(_06088_));
 sky130_fd_sc_hd__or4_1 _12913_ (.A(net4737),
    .B(net4690),
    .C(net4694),
    .D(net4584),
    .X(_06089_));
 sky130_fd_sc_hd__or4_1 _12914_ (.A(net4576),
    .B(net4550),
    .C(net4293),
    .D(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__or4_1 _12915_ (.A(net4777),
    .B(net4674),
    .C(_06088_),
    .D(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__inv_4 _12916_ (.A(net8034),
    .Y(_06092_));
 sky130_fd_sc_hd__o211a_1 _12917_ (.A1(_06075_),
    .A2(_06087_),
    .B1(net4778),
    .C1(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__xnor2_1 _12918_ (.A(net4384),
    .B(net4044),
    .Y(_06094_));
 sky130_fd_sc_hd__o221a_1 _12919_ (.A1(_04731_),
    .A2(net3893),
    .B1(_06048_),
    .B2(net4357),
    .C1(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__o221a_1 _12920_ (.A1(net2587),
    .A2(_06061_),
    .B1(net4642),
    .B2(net4366),
    .C1(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__or4_1 _12921_ (.A(_06039_),
    .B(net3848),
    .C(net4044),
    .D(net3807),
    .X(_06097_));
 sky130_fd_sc_hd__nor2_1 _12922_ (.A(net3893),
    .B(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__xor2_1 _12923_ (.A(net4393),
    .B(net3848),
    .X(_06099_));
 sky130_fd_sc_hd__a221o_1 _12924_ (.A1(net4366),
    .A2(net4642),
    .B1(_06048_),
    .B2(net4357),
    .C1(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__nor2_1 _12925_ (.A(_06098_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__and3_1 _12926_ (.A(net4779),
    .B(net4643),
    .C(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__a21oi_1 _12927_ (.A1(net3983),
    .A2(_04743_),
    .B1(_06060_),
    .Y(_06103_));
 sky130_fd_sc_hd__clkbuf_4 _12928_ (.A(net7687),
    .X(_06104_));
 sky130_fd_sc_hd__or2_1 _12929_ (.A(net4354),
    .B(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__nand2_1 _12930_ (.A(net4354),
    .B(_06104_),
    .Y(_06106_));
 sky130_fd_sc_hd__clkbuf_1 _12931_ (.A(net3964),
    .X(_06107_));
 sky130_fd_sc_hd__inv_2 _12932_ (.A(net4420),
    .Y(_06108_));
 sky130_fd_sc_hd__clkbuf_1 _12933_ (.A(net3998),
    .X(_06109_));
 sky130_fd_sc_hd__xor2_1 _12934_ (.A(net4431),
    .B(net3999),
    .X(_06110_));
 sky130_fd_sc_hd__a221o_1 _12935_ (.A1(_04738_),
    .A2(net4034),
    .B1(net3965),
    .B2(_06108_),
    .C1(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__a221o_1 _12936_ (.A1(net4369),
    .A2(_06068_),
    .B1(_06105_),
    .B2(_06106_),
    .C1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__a221o_1 _12937_ (.A1(net4420),
    .A2(_06062_),
    .B1(_06060_),
    .B2(net3983),
    .C1(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__or3b_1 _12938_ (.A(net3984),
    .B(_06113_),
    .C_N(_06093_),
    .X(_06114_));
 sky130_fd_sc_hd__or2b_2 _12939_ (.A(net4644),
    .B_N(net3985),
    .X(_06115_));
 sky130_fd_sc_hd__nor2_1 _12940_ (.A(_06056_),
    .B(net4645),
    .Y(_06116_));
 sky130_fd_sc_hd__and2b_1 _12941_ (.A_N(net5922),
    .B(net3975),
    .X(_06117_));
 sky130_fd_sc_hd__and3b_2 _12942_ (.A_N(_04485_),
    .B(_06117_),
    .C(net3773),
    .X(_06118_));
 sky130_fd_sc_hd__clkbuf_4 _12943_ (.A(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__buf_4 _12944_ (.A(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__buf_4 _12945_ (.A(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__clkbuf_4 _12946_ (.A(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__clkbuf_4 _12947_ (.A(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__buf_4 _12948_ (.A(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__xor2_1 _12949_ (.A(net3965),
    .B(net4044),
    .X(_06125_));
 sky130_fd_sc_hd__o221a_1 _12950_ (.A1(_06068_),
    .A2(_06061_),
    .B1(_06043_),
    .B2(net3960),
    .C1(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__o2bb2a_1 _12951_ (.A1_N(net3999),
    .A2_N(_06039_),
    .B1(net3848),
    .B2(_06104_),
    .X(_06127_));
 sky130_fd_sc_hd__o221a_1 _12952_ (.A1(net4034),
    .A2(net3893),
    .B1(_06039_),
    .B2(net3999),
    .C1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__and4_1 _12953_ (.A(net3960),
    .B(_06062_),
    .C(_06061_),
    .D(_06043_),
    .X(_06129_));
 sky130_fd_sc_hd__and4_1 _12954_ (.A(net3999),
    .B(_06039_),
    .C(_06035_),
    .D(_06048_),
    .X(_06130_));
 sky130_fd_sc_hd__and4_1 _12955_ (.A(_06068_),
    .B(net4007),
    .C(_06129_),
    .D(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__a21oi_1 _12956_ (.A1(_06126_),
    .A2(_06128_),
    .B1(net4008),
    .Y(_06132_));
 sky130_fd_sc_hd__and4_1 _12957_ (.A(_06039_),
    .B(net3848),
    .C(net4044),
    .D(net3807),
    .X(_06133_));
 sky130_fd_sc_hd__and3_1 _12958_ (.A(net3965),
    .B(net3999),
    .C(_06060_),
    .X(_06134_));
 sky130_fd_sc_hd__xnor2_1 _12959_ (.A(net3893),
    .B(_06039_),
    .Y(_06135_));
 sky130_fd_sc_hd__a22o_1 _12960_ (.A1(net3960),
    .A2(_06061_),
    .B1(_06135_),
    .B2(net4034),
    .X(_06136_));
 sky130_fd_sc_hd__or4_1 _12961_ (.A(_06104_),
    .B(net4034),
    .C(net3965),
    .D(_06060_),
    .X(_06137_));
 sky130_fd_sc_hd__a21o_1 _12962_ (.A1(_06062_),
    .A2(_06043_),
    .B1(net4044),
    .X(_06138_));
 sky130_fd_sc_hd__a22o_1 _12963_ (.A1(net3960),
    .A2(_06061_),
    .B1(net3848),
    .B2(net3965),
    .X(_06139_));
 sky130_fd_sc_hd__a22o_1 _12964_ (.A1(_06104_),
    .A2(net3893),
    .B1(_06039_),
    .B2(net4034),
    .X(_06140_));
 sky130_fd_sc_hd__a2111o_1 _12965_ (.A1(_06068_),
    .A2(net4642),
    .B1(_06138_),
    .C1(_06139_),
    .D1(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__a21oi_1 _12966_ (.A1(_06137_),
    .A2(_06141_),
    .B1(net3999),
    .Y(_06142_));
 sky130_fd_sc_hd__a31o_1 _12967_ (.A1(net3965),
    .A2(net3848),
    .A3(_06136_),
    .B1(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__a311o_1 _12968_ (.A1(_06104_),
    .A2(net4034),
    .A3(_06134_),
    .B1(_06143_),
    .C1(_06129_),
    .X(_06144_));
 sky130_fd_sc_hd__a211oi_1 _12969_ (.A1(net3893),
    .A2(_06133_),
    .B1(_06144_),
    .C1(_06098_),
    .Y(_06145_));
 sky130_fd_sc_hd__nand2_1 _12970_ (.A(net4009),
    .B(net5975),
    .Y(_06146_));
 sky130_fd_sc_hd__xnor2_1 _12971_ (.A(net2185),
    .B(net4049),
    .Y(_06147_));
 sky130_fd_sc_hd__o221a_1 _12972_ (.A1(_04718_),
    .A2(net4034),
    .B1(net3807),
    .B2(_04721_),
    .C1(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__xor2_1 _12973_ (.A(net4152),
    .B(_06104_),
    .X(_06149_));
 sky130_fd_sc_hd__a221oi_1 _12974_ (.A1(net1817),
    .A2(_06061_),
    .B1(_06043_),
    .B2(net4324),
    .C1(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__xnor2_1 _12975_ (.A(net4347),
    .B(net3999),
    .Y(_06151_));
 sky130_fd_sc_hd__xnor2_1 _12976_ (.A(net2038),
    .B(_06039_),
    .Y(_06152_));
 sky130_fd_sc_hd__o22a_1 _12977_ (.A1(net1817),
    .A2(_06061_),
    .B1(_06043_),
    .B2(net4324),
    .X(_06153_));
 sky130_fd_sc_hd__o221a_1 _12978_ (.A1(net4315),
    .A2(_06062_),
    .B1(_06048_),
    .B2(net1803),
    .C1(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__xnor2_1 _12979_ (.A(net4306),
    .B(net4044),
    .Y(_06155_));
 sky130_fd_sc_hd__o221a_1 _12980_ (.A1(net4309),
    .A2(_06068_),
    .B1(net3965),
    .B2(_04722_),
    .C1(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__and4_1 _12981_ (.A(_06151_),
    .B(_06152_),
    .C(_06154_),
    .D(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__and4_1 _12982_ (.A(net4779),
    .B(_06148_),
    .C(_06150_),
    .D(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__a21oi_1 _12983_ (.A1(net4779),
    .A2(_06146_),
    .B1(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__o31a_1 _12984_ (.A1(_06056_),
    .A2(net4645),
    .A3(net4780),
    .B1(_04479_),
    .X(_06160_));
 sky130_fd_sc_hd__o21a_1 _12985_ (.A1(net4646),
    .A2(_06124_),
    .B1(net4781),
    .X(_06161_));
 sky130_fd_sc_hd__inv_2 _12986_ (.A(net4498),
    .Y(_06162_));
 sky130_fd_sc_hd__and2_2 _12987_ (.A(_06162_),
    .B(net4742),
    .X(_06163_));
 sky130_fd_sc_hd__inv_2 _12988_ (.A(net4569),
    .Y(_06164_));
 sky130_fd_sc_hd__inv_2 _12989_ (.A(net3945),
    .Y(_06165_));
 sky130_fd_sc_hd__a22o_1 _12990_ (.A1(_06164_),
    .A2(net3787),
    .B1(_06165_),
    .B2(net3932),
    .X(_06166_));
 sky130_fd_sc_hd__inv_2 _12991_ (.A(net3926),
    .Y(_06167_));
 sky130_fd_sc_hd__o22a_1 _12992_ (.A1(_06162_),
    .A2(net4742),
    .B1(net4762),
    .B2(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__inv_2 _12993_ (.A(net3768),
    .Y(_06169_));
 sky130_fd_sc_hd__inv_2 _12994_ (.A(net3757),
    .Y(_06170_));
 sky130_fd_sc_hd__o22a_1 _12995_ (.A1(net4500),
    .A2(_06169_),
    .B1(net4508),
    .B2(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__inv_2 _12996_ (.A(net3932),
    .Y(_06172_));
 sky130_fd_sc_hd__nor2_1 _12997_ (.A(_06164_),
    .B(net3787),
    .Y(_06173_));
 sky130_fd_sc_hd__inv_2 _12998_ (.A(net4667),
    .Y(_06174_));
 sky130_fd_sc_hd__inv_2 _12999_ (.A(net4518),
    .Y(_06175_));
 sky130_fd_sc_hd__a2bb2o_1 _13000_ (.A1_N(net3749),
    .A2_N(_06174_),
    .B1(net4506),
    .B2(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__inv_2 _13001_ (.A(net4541),
    .Y(_06177_));
 sky130_fd_sc_hd__nor2_1 _13002_ (.A(net4565),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__inv_2 _13003_ (.A(net4547),
    .Y(_06179_));
 sky130_fd_sc_hd__nor2_1 _13004_ (.A(_06179_),
    .B(net3847),
    .Y(_06180_));
 sky130_fd_sc_hd__and2_1 _13005_ (.A(net4508),
    .B(_06170_),
    .X(_06181_));
 sky130_fd_sc_hd__and2_1 _13006_ (.A(net4762),
    .B(_06167_),
    .X(_06182_));
 sky130_fd_sc_hd__or4_1 _13007_ (.A(_06178_),
    .B(_06180_),
    .C(_06181_),
    .D(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__a22o_1 _13008_ (.A1(_06179_),
    .A2(net3847),
    .B1(net4565),
    .B2(_06177_),
    .X(_06184_));
 sky130_fd_sc_hd__and2_1 _13009_ (.A(net4500),
    .B(_06169_),
    .X(_06185_));
 sky130_fd_sc_hd__a211o_1 _13010_ (.A1(net3749),
    .A2(_06174_),
    .B1(_06184_),
    .C1(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__or2_1 _13011_ (.A(net4506),
    .B(_06175_),
    .X(_06187_));
 sky130_fd_sc_hd__or4b_1 _13012_ (.A(_06176_),
    .B(_06183_),
    .C(_06186_),
    .D_N(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__a2111oi_1 _13013_ (.A1(net3945),
    .A2(_06172_),
    .B1(_06163_),
    .C1(_06173_),
    .D1(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__and4b_1 _13014_ (.A_N(_06166_),
    .B(_06168_),
    .C(_06171_),
    .D(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__inv_2 _13015_ (.A(net4723),
    .Y(_06191_));
 sky130_fd_sc_hd__inv_2 _13016_ (.A(net3835),
    .Y(_06192_));
 sky130_fd_sc_hd__o2bb2a_1 _13017_ (.A1_N(net3820),
    .A2_N(_06191_),
    .B1(_06192_),
    .B2(net4655),
    .X(_06193_));
 sky130_fd_sc_hd__inv_2 _13018_ (.A(net3875),
    .Y(_06194_));
 sky130_fd_sc_hd__and2_1 _13019_ (.A(net4655),
    .B(_06192_),
    .X(_06195_));
 sky130_fd_sc_hd__o21ba_1 _13020_ (.A1(_06194_),
    .A2(net4575),
    .B1_N(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__o211a_1 _13021_ (.A1(_06191_),
    .A2(net3820),
    .B1(_06193_),
    .C1(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__inv_2 _13022_ (.A(net4659),
    .Y(_06198_));
 sky130_fd_sc_hd__a22o_1 _13023_ (.A1(_06194_),
    .A2(net4575),
    .B1(net3803),
    .B2(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__o21ba_1 _13024_ (.A1(net3803),
    .A2(_06198_),
    .B1_N(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__inv_2 _13025_ (.A(net4581),
    .Y(_06201_));
 sky130_fd_sc_hd__inv_2 _13026_ (.A(net4665),
    .Y(_06202_));
 sky130_fd_sc_hd__o22a_1 _13027_ (.A1(_06201_),
    .A2(net3790),
    .B1(_06202_),
    .B2(net4567),
    .X(_06203_));
 sky130_fd_sc_hd__inv_2 _13028_ (.A(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__inv_2 _13029_ (.A(net3785),
    .Y(_06205_));
 sky130_fd_sc_hd__a2bb2o_1 _13030_ (.A1_N(_06205_),
    .A2_N(net3888),
    .B1(_06202_),
    .B2(net4567),
    .X(_06206_));
 sky130_fd_sc_hd__inv_2 _13031_ (.A(net4669),
    .Y(_06207_));
 sky130_fd_sc_hd__a22o_1 _13032_ (.A1(_06207_),
    .A2(net4526),
    .B1(_06201_),
    .B2(net3790),
    .X(_06208_));
 sky130_fd_sc_hd__inv_2 _13033_ (.A(net3751),
    .Y(_06209_));
 sky130_fd_sc_hd__a2bb2o_1 _13034_ (.A1_N(_06207_),
    .A2_N(net4526),
    .B1(_06209_),
    .B2(net4589),
    .X(_06210_));
 sky130_fd_sc_hd__or4_1 _13035_ (.A(_06204_),
    .B(_06206_),
    .C(_06208_),
    .D(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__inv_2 _13036_ (.A(net4651),
    .Y(_06212_));
 sky130_fd_sc_hd__inv_2 _13037_ (.A(net4610),
    .Y(_06213_));
 sky130_fd_sc_hd__a22o_1 _13038_ (.A1(_06212_),
    .A2(net3669),
    .B1(_06213_),
    .B2(net3811),
    .X(_06214_));
 sky130_fd_sc_hd__nor2_1 _13039_ (.A(_06212_),
    .B(net3669),
    .Y(_06215_));
 sky130_fd_sc_hd__a211o_1 _13040_ (.A1(_06205_),
    .A2(net3888),
    .B1(_06214_),
    .C1(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__inv_2 _13041_ (.A(net4657),
    .Y(_06217_));
 sky130_fd_sc_hd__o22a_1 _13042_ (.A1(_06213_),
    .A2(net3811),
    .B1(_06217_),
    .B2(net3766),
    .X(_06218_));
 sky130_fd_sc_hd__o2bb2a_1 _13043_ (.A1_N(_06217_),
    .A2_N(net3766),
    .B1(_06209_),
    .B2(net4589),
    .X(_06219_));
 sky130_fd_sc_hd__and4bb_1 _13044_ (.A_N(_06211_),
    .B_N(_06216_),
    .C(_06218_),
    .D(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__nor2_1 _13045_ (.A(_06173_),
    .B(_06178_),
    .Y(_06221_));
 sky130_fd_sc_hd__o2bb2a_1 _13046_ (.A1_N(_06187_),
    .A2_N(_06176_),
    .B1(_06165_),
    .B2(net3729),
    .X(_06222_));
 sky130_fd_sc_hd__or2_1 _13047_ (.A(_06166_),
    .B(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__a21oi_1 _13048_ (.A1(_06221_),
    .A2(_06223_),
    .B1(_06184_),
    .Y(_06224_));
 sky130_fd_sc_hd__o31a_1 _13049_ (.A1(_06180_),
    .A2(_06181_),
    .A3(_06224_),
    .B1(_06171_),
    .X(_06225_));
 sky130_fd_sc_hd__nor2_1 _13050_ (.A(_06185_),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__a21oi_1 _13051_ (.A1(_06203_),
    .A2(_06206_),
    .B1(_06208_),
    .Y(_06227_));
 sky130_fd_sc_hd__o21ai_1 _13052_ (.A1(_06210_),
    .A2(_06227_),
    .B1(_06219_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21oi_1 _13053_ (.A1(_06218_),
    .A2(_06228_),
    .B1(_06214_),
    .Y(_06229_));
 sky130_fd_sc_hd__o2bb2a_1 _13054_ (.A1_N(_06220_),
    .A2_N(_06226_),
    .B1(_06229_),
    .B2(_06215_),
    .X(_06230_));
 sky130_fd_sc_hd__nand3b_1 _13055_ (.A_N(_06230_),
    .B(_06200_),
    .C(_06197_),
    .Y(_06231_));
 sky130_fd_sc_hd__nand2_1 _13056_ (.A(_06197_),
    .B(_06199_),
    .Y(_06232_));
 sky130_fd_sc_hd__o211a_1 _13057_ (.A1(_06193_),
    .A2(_06195_),
    .B1(_06231_),
    .C1(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__o21a_1 _13058_ (.A1(_06182_),
    .A2(_06233_),
    .B1(_06168_),
    .X(_06234_));
 sky130_fd_sc_hd__a41o_1 _13059_ (.A1(_06190_),
    .A2(_06197_),
    .A3(_06200_),
    .A4(_06220_),
    .B1(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__and2_1 _13060_ (.A(net4646),
    .B(net4780),
    .X(_06236_));
 sky130_fd_sc_hd__buf_2 _13061_ (.A(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__or3b_1 _13062_ (.A(_06163_),
    .B(_06235_),
    .C_N(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__buf_2 _13063_ (.A(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__nand2_2 _13064_ (.A(net4647),
    .B(_06239_),
    .Y(_06240_));
 sky130_fd_sc_hd__nor2_2 _13065_ (.A(_06058_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__clkbuf_4 _13066_ (.A(_06240_),
    .X(_06242_));
 sky130_fd_sc_hd__a32o_1 _13067_ (.A1(_06053_),
    .A2(_06054_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(net5605),
    .X(_00386_));
 sky130_fd_sc_hd__xor2_1 _13068_ (.A(net5531),
    .B(_06028_),
    .X(_06243_));
 sky130_fd_sc_hd__buf_2 _13069_ (.A(_06028_),
    .X(_06244_));
 sky130_fd_sc_hd__a21bo_1 _13070_ (.A1(net2277),
    .A2(_06244_),
    .B1_N(_06054_),
    .X(_06245_));
 sky130_fd_sc_hd__xor2_1 _13071_ (.A(_06243_),
    .B(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__a22o_1 _13072_ (.A1(net5531),
    .A2(_06242_),
    .B1(_06241_),
    .B2(_06246_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _13073_ (.A(net5428),
    .B(_06244_),
    .X(_06247_));
 sky130_fd_sc_hd__nor2_1 _13074_ (.A(net5428),
    .B(_06244_),
    .Y(_06248_));
 sky130_fd_sc_hd__nor2_1 _13075_ (.A(_06247_),
    .B(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__and4_1 _13076_ (.A(_06029_),
    .B(_06031_),
    .C(_06050_),
    .D(_06243_),
    .X(_06250_));
 sky130_fd_sc_hd__o21a_1 _13077_ (.A1(net5531),
    .A2(net5605),
    .B1(_06244_),
    .X(_06251_));
 sky130_fd_sc_hd__or3_1 _13078_ (.A(_06051_),
    .B(_06250_),
    .C(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__xor2_1 _13079_ (.A(_06249_),
    .B(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__a22o_1 _13080_ (.A1(net5428),
    .A2(_06242_),
    .B1(_06241_),
    .B2(_06253_),
    .X(_00388_));
 sky130_fd_sc_hd__xnor2_1 _13081_ (.A(net5618),
    .B(_06244_),
    .Y(_06254_));
 sky130_fd_sc_hd__a21oi_1 _13082_ (.A1(_06249_),
    .A2(_06252_),
    .B1(_06247_),
    .Y(_06255_));
 sky130_fd_sc_hd__nand2_1 _13083_ (.A(_06254_),
    .B(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__or2_1 _13084_ (.A(_06254_),
    .B(_06255_),
    .X(_06257_));
 sky130_fd_sc_hd__a32o_1 _13085_ (.A1(_06241_),
    .A2(_06256_),
    .A3(_06257_),
    .B1(_06242_),
    .B2(net5618),
    .X(_00389_));
 sky130_fd_sc_hd__o21ba_1 _13086_ (.A1(net2058),
    .A2(_06244_),
    .B1_N(_06255_),
    .X(_06258_));
 sky130_fd_sc_hd__a21oi_1 _13087_ (.A1(net2058),
    .A2(_06244_),
    .B1(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__xnor2_1 _13088_ (.A(net5408),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__nand2_1 _13089_ (.A(_06244_),
    .B(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__or2_1 _13090_ (.A(_06244_),
    .B(_06260_),
    .X(_06262_));
 sky130_fd_sc_hd__a32o_1 _13091_ (.A1(_06241_),
    .A2(_06261_),
    .A3(_06262_),
    .B1(_06242_),
    .B2(net5408),
    .X(_00390_));
 sky130_fd_sc_hd__a211oi_4 _13092_ (.A1(_05980_),
    .A2(_05983_),
    .B1(net8051),
    .C1(_05984_),
    .Y(_06263_));
 sky130_fd_sc_hd__nor2_2 _13093_ (.A(net8217),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__clkbuf_4 _13094_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06265_));
 sky130_fd_sc_hd__buf_2 _13095_ (.A(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__or2_1 _13096_ (.A(net8265),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__or2_1 _13097_ (.A(net4446),
    .B(net4828),
    .X(_06268_));
 sky130_fd_sc_hd__or2_2 _13098_ (.A(net4513),
    .B(net6015),
    .X(_06269_));
 sky130_fd_sc_hd__nor2_1 _13099_ (.A(net4462),
    .B(net3604),
    .Y(_06270_));
 sky130_fd_sc_hd__xor2_2 _13100_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_06271_));
 sky130_fd_sc_hd__and2_1 _13101_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_06272_));
 sky130_fd_sc_hd__a31oi_2 _13102_ (.A1(\rbzero.debug_overlay.facingX[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A3(_06271_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nor2_1 _13103_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06274_));
 sky130_fd_sc_hd__nand2_1 _13104_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06275_));
 sky130_fd_sc_hd__o21a_2 _13105_ (.A1(_06273_),
    .A2(_06274_),
    .B1(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__nand2_1 _13106_ (.A(net4462),
    .B(net3604),
    .Y(_06277_));
 sky130_fd_sc_hd__o21ai_4 _13107_ (.A1(_06270_),
    .A2(_06276_),
    .B1(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__and2_1 _13108_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06279_));
 sky130_fd_sc_hd__nor2_1 _13109_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_06280_));
 sky130_fd_sc_hd__nor2_2 _13110_ (.A(_06279_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_1 _13111_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_06282_));
 sky130_fd_sc_hd__or2_1 _13112_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06283_));
 sky130_fd_sc_hd__and3_1 _13113_ (.A(_06281_),
    .B(_06282_),
    .C(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__nand2_1 _13114_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_06285_));
 sky130_fd_sc_hd__inv_2 _13115_ (.A(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__nor2_1 _13116_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_06287_));
 sky130_fd_sc_hd__nor2_1 _13117_ (.A(_06286_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__and2_1 _13118_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_06289_));
 sky130_fd_sc_hd__nor2_1 _13119_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_06290_));
 sky130_fd_sc_hd__nor2_2 _13120_ (.A(_06289_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__and3_1 _13121_ (.A(_06284_),
    .B(_06288_),
    .C(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__o21ba_1 _13122_ (.A1(_06286_),
    .A2(_06289_),
    .B1_N(_06287_),
    .X(_06293_));
 sky130_fd_sc_hd__and2_1 _13123_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06294_));
 sky130_fd_sc_hd__a221o_1 _13124_ (.A1(_06279_),
    .A2(_06283_),
    .B1(_06284_),
    .B2(_06293_),
    .C1(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__a21o_1 _13125_ (.A1(_06278_),
    .A2(_06292_),
    .B1(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__and2_1 _13126_ (.A(net3719),
    .B(net3614),
    .X(_06297_));
 sky130_fd_sc_hd__nor2_1 _13127_ (.A(net3719),
    .B(net3614),
    .Y(_06298_));
 sky130_fd_sc_hd__nor2_1 _13128_ (.A(_06297_),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__a221o_1 _13129_ (.A1(net4513),
    .A2(net6015),
    .B1(_06296_),
    .B2(_06299_),
    .C1(_06297_),
    .X(_06300_));
 sky130_fd_sc_hd__and2_1 _13130_ (.A(net4446),
    .B(net4828),
    .X(_06301_));
 sky130_fd_sc_hd__nor2_1 _13131_ (.A(net4446),
    .B(net5952),
    .Y(_06302_));
 sky130_fd_sc_hd__a311o_2 _13132_ (.A1(_06268_),
    .A2(_06269_),
    .A3(_06300_),
    .B1(_06301_),
    .C1(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__nand2_2 _13133_ (.A(net4446),
    .B(net5952),
    .Y(_06304_));
 sky130_fd_sc_hd__inv_2 _13134_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06305_));
 sky130_fd_sc_hd__clkbuf_4 _13135_ (.A(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__a21oi_4 _13136_ (.A1(_06303_),
    .A2(_06304_),
    .B1(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__a21oi_2 _13137_ (.A1(_06264_),
    .A2(_06267_),
    .B1(_06307_),
    .Y(_06308_));
 sky130_fd_sc_hd__or2_1 _13138_ (.A(net8267),
    .B(_06266_),
    .X(_06309_));
 sky130_fd_sc_hd__a21oi_4 _13139_ (.A1(_06264_),
    .A2(_06309_),
    .B1(_06307_),
    .Y(_06310_));
 sky130_fd_sc_hd__nand2_2 _13140_ (.A(_06282_),
    .B(_06283_),
    .Y(_06311_));
 sky130_fd_sc_hd__a31o_1 _13141_ (.A1(_06288_),
    .A2(_06278_),
    .A3(_06291_),
    .B1(_06293_),
    .X(_06312_));
 sky130_fd_sc_hd__a21o_1 _13142_ (.A1(_06281_),
    .A2(_06312_),
    .B1(_06279_),
    .X(_06313_));
 sky130_fd_sc_hd__xnor2_4 _13143_ (.A(_06311_),
    .B(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__nor2_1 _13144_ (.A(net8263),
    .B(_06265_),
    .Y(_06315_));
 sky130_fd_sc_hd__a211oi_1 _13145_ (.A1(_06265_),
    .A2(_06025_),
    .B1(_06315_),
    .C1(_04491_),
    .Y(_06316_));
 sky130_fd_sc_hd__xor2_2 _13146_ (.A(_06281_),
    .B(_06312_),
    .X(_06317_));
 sky130_fd_sc_hd__mux2_1 _13147_ (.A0(net4293),
    .A1(_05997_),
    .S(_06265_),
    .X(_06318_));
 sky130_fd_sc_hd__mux2_4 _13148_ (.A0(_06317_),
    .A1(_06318_),
    .S(_06306_),
    .X(_06319_));
 sky130_fd_sc_hd__a21oi_1 _13149_ (.A1(_06278_),
    .A2(_06291_),
    .B1(_06289_),
    .Y(_06320_));
 sky130_fd_sc_hd__xnor2_2 _13150_ (.A(_06288_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__nor2_1 _13151_ (.A(net4280),
    .B(_06265_),
    .Y(_06322_));
 sky130_fd_sc_hd__a211oi_2 _13152_ (.A1(_06265_),
    .A2(_06015_),
    .B1(_06322_),
    .C1(_04491_),
    .Y(_06323_));
 sky130_fd_sc_hd__xor2_2 _13153_ (.A(_06278_),
    .B(_06291_),
    .X(_06324_));
 sky130_fd_sc_hd__and2_1 _13154_ (.A(net4236),
    .B(net8051),
    .X(_06325_));
 sky130_fd_sc_hd__a31o_1 _13155_ (.A1(_06265_),
    .A2(_06000_),
    .A3(_06001_),
    .B1(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__mux2_4 _13156_ (.A0(_06324_),
    .A1(_06326_),
    .S(_06306_),
    .X(_06327_));
 sky130_fd_sc_hd__or2_1 _13157_ (.A(net4268),
    .B(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06328_));
 sky130_fd_sc_hd__o21ai_2 _13158_ (.A1(net8051),
    .A2(_06006_),
    .B1(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__and2b_1 _13159_ (.A_N(_06270_),
    .B(_06277_),
    .X(_06330_));
 sky130_fd_sc_hd__xnor2_2 _13160_ (.A(_06276_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__nand2_1 _13161_ (.A(_04491_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__and2b_1 _13162_ (.A_N(_06274_),
    .B(_06275_),
    .X(_06333_));
 sky130_fd_sc_hd__xnor2_1 _13163_ (.A(_06273_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__or2_1 _13164_ (.A(_06305_),
    .B(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__and2_1 _13165_ (.A(net4277),
    .B(net8051),
    .X(_06336_));
 sky130_fd_sc_hd__a211o_1 _13166_ (.A1(_06265_),
    .A2(_06007_),
    .B1(_06336_),
    .C1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06337_));
 sky130_fd_sc_hd__mux2_2 _13167_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_06009_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06338_));
 sky130_fd_sc_hd__nand2_1 _13168_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_06339_));
 sky130_fd_sc_hd__xnor2_1 _13169_ (.A(_06339_),
    .B(_06271_),
    .Y(_06340_));
 sky130_fd_sc_hd__and2_1 _13170_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .B(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__mux2_4 _13171_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06342_));
 sky130_fd_sc_hd__mux2_4 _13172_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_06342_),
    .S(_06305_),
    .X(_06343_));
 sky130_fd_sc_hd__mux2_4 _13173_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06344_));
 sky130_fd_sc_hd__mux2_4 _13174_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_06344_),
    .S(_06305_),
    .X(_06345_));
 sky130_fd_sc_hd__or2_4 _13175_ (.A(_06343_),
    .B(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_06010_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06347_));
 sky130_fd_sc_hd__or2_1 _13177_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_06348_));
 sky130_fd_sc_hd__and2_1 _13178_ (.A(_06339_),
    .B(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__mux2_4 _13179_ (.A0(_06347_),
    .A1(_06349_),
    .S(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06350_));
 sky130_fd_sc_hd__a2111o_1 _13180_ (.A1(_06305_),
    .A2(_06338_),
    .B1(_06341_),
    .C1(_06346_),
    .D1(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__a21oi_2 _13181_ (.A1(_06335_),
    .A2(_06337_),
    .B1(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__o211ai_2 _13182_ (.A1(_04491_),
    .A2(_06329_),
    .B1(_06332_),
    .C1(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__a2111o_1 _13183_ (.A1(_04491_),
    .A2(_06321_),
    .B1(_06323_),
    .C1(_06327_),
    .D1(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__a2111o_1 _13184_ (.A1(_04491_),
    .A2(_06314_),
    .B1(_06316_),
    .C1(_06319_),
    .D1(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__o21ai_1 _13185_ (.A1(_06018_),
    .A2(_06019_),
    .B1(_06266_),
    .Y(_06356_));
 sky130_fd_sc_hd__o21a_1 _13186_ (.A1(net8269),
    .A2(_06265_),
    .B1(_06306_),
    .X(_06357_));
 sky130_fd_sc_hd__nand2_1 _13187_ (.A(net4513),
    .B(net6015),
    .Y(_06358_));
 sky130_fd_sc_hd__nand2_1 _13188_ (.A(_06269_),
    .B(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__a21o_1 _13189_ (.A1(_06296_),
    .A2(_06299_),
    .B1(_06297_),
    .X(_06360_));
 sky130_fd_sc_hd__xnor2_2 _13190_ (.A(_06359_),
    .B(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__a21o_1 _13191_ (.A1(_05976_),
    .A2(_05998_),
    .B1(net8051),
    .X(_06362_));
 sky130_fd_sc_hd__o21a_1 _13192_ (.A1(net8021),
    .A2(_06265_),
    .B1(_06306_),
    .X(_06363_));
 sky130_fd_sc_hd__xor2_2 _13193_ (.A(_06296_),
    .B(_06299_),
    .X(_06364_));
 sky130_fd_sc_hd__a22o_2 _13194_ (.A1(_06362_),
    .A2(_06363_),
    .B1(_06364_),
    .B2(_04491_),
    .X(_06365_));
 sky130_fd_sc_hd__a221o_1 _13195_ (.A1(_06356_),
    .A2(_06357_),
    .B1(_06361_),
    .B2(net8217),
    .C1(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__nor2_2 _13196_ (.A(_06355_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__a31o_2 _13197_ (.A1(_06268_),
    .A2(_06269_),
    .A3(_06300_),
    .B1(_06301_),
    .X(_06368_));
 sky130_fd_sc_hd__and2b_1 _13198_ (.A_N(_06302_),
    .B(_06304_),
    .X(_06369_));
 sky130_fd_sc_hd__xnor2_4 _13199_ (.A(_06368_),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_1 _13200_ (.A(net4446),
    .B(net4828),
    .Y(_06371_));
 sky130_fd_sc_hd__nor2_1 _13201_ (.A(_06371_),
    .B(_06301_),
    .Y(_06372_));
 sky130_fd_sc_hd__inv_2 _13202_ (.A(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__nand3_1 _13203_ (.A(_06269_),
    .B(_06300_),
    .C(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__a21o_1 _13204_ (.A1(_06269_),
    .A2(_06300_),
    .B1(_06373_),
    .X(_06375_));
 sky130_fd_sc_hd__a21oi_1 _13205_ (.A1(net4917),
    .A2(net8051),
    .B1(_04491_),
    .Y(_06376_));
 sky130_fd_sc_hd__o31a_1 _13206_ (.A1(net8051),
    .A2(_05992_),
    .A3(_05994_),
    .B1(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__a31o_2 _13207_ (.A1(net8217),
    .A2(_06374_),
    .A3(_06375_),
    .B1(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__nor2_1 _13208_ (.A(net8261),
    .B(_06266_),
    .Y(_06379_));
 sky130_fd_sc_hd__a311o_1 _13209_ (.A1(_06266_),
    .A2(_05987_),
    .A3(_05988_),
    .B1(_06379_),
    .C1(net8217),
    .X(_06380_));
 sky130_fd_sc_hd__o211a_1 _13210_ (.A1(_06306_),
    .A2(_06370_),
    .B1(_06378_),
    .C1(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__a21o_1 _13211_ (.A1(_06303_),
    .A2(_06304_),
    .B1(_06306_),
    .X(_06382_));
 sky130_fd_sc_hd__a211o_4 _13212_ (.A1(net8035),
    .A2(net8051),
    .B1(_04491_),
    .C1(_06263_),
    .X(_06383_));
 sky130_fd_sc_hd__and2_1 _13213_ (.A(_06382_),
    .B(_06383_),
    .X(_06384_));
 sky130_fd_sc_hd__clkbuf_4 _13214_ (.A(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__a41o_1 _13215_ (.A1(_06308_),
    .A2(_06310_),
    .A3(_06367_),
    .A4(_06381_),
    .B1(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__o21a_1 _13216_ (.A1(net8015),
    .A2(_06266_),
    .B1(_06264_),
    .X(_06387_));
 sky130_fd_sc_hd__or2_2 _13217_ (.A(_06307_),
    .B(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__xnor2_2 _13218_ (.A(_06386_),
    .B(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__a22o_1 _13219_ (.A1(_06356_),
    .A2(_06357_),
    .B1(_06361_),
    .B2(net8217),
    .X(_06390_));
 sky130_fd_sc_hd__o2bb2a_4 _13220_ (.A1_N(_06382_),
    .A2_N(_06383_),
    .B1(_06365_),
    .B2(_06355_),
    .X(_06391_));
 sky130_fd_sc_hd__xor2_4 _13221_ (.A(_06390_),
    .B(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__o2bb2a_4 _13222_ (.A1_N(_06382_),
    .A2_N(_06383_),
    .B1(_06355_),
    .B2(_06366_),
    .X(_06393_));
 sky130_fd_sc_hd__xnor2_4 _13223_ (.A(_06378_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__or2_4 _13224_ (.A(_06392_),
    .B(_06394_),
    .X(_06395_));
 sky130_fd_sc_hd__o21a_1 _13225_ (.A1(_06306_),
    .A2(_06370_),
    .B1(_06380_),
    .X(_06396_));
 sky130_fd_sc_hd__a21oi_1 _13226_ (.A1(_06378_),
    .A2(_06367_),
    .B1(_06385_),
    .Y(_06397_));
 sky130_fd_sc_hd__xnor2_2 _13227_ (.A(_06396_),
    .B(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__or2_4 _13228_ (.A(_06395_),
    .B(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__a31o_1 _13229_ (.A1(_06310_),
    .A2(_06367_),
    .A3(_06381_),
    .B1(_06385_),
    .X(_06400_));
 sky130_fd_sc_hd__xor2_2 _13230_ (.A(_06308_),
    .B(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__a21oi_2 _13231_ (.A1(_06367_),
    .A2(_06381_),
    .B1(_06385_),
    .Y(_06402_));
 sky130_fd_sc_hd__xnor2_4 _13232_ (.A(_06310_),
    .B(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2_4 _13233_ (.A(_06382_),
    .B(_06383_),
    .Y(_06404_));
 sky130_fd_sc_hd__and2_1 _13234_ (.A(_06404_),
    .B(_06355_),
    .X(_06405_));
 sky130_fd_sc_hd__xor2_2 _13235_ (.A(_06365_),
    .B(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__or4_4 _13236_ (.A(_06399_),
    .B(_06401_),
    .C(_06403_),
    .D(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__or2_1 _13237_ (.A(net8002),
    .B(_06266_),
    .X(_06408_));
 sky130_fd_sc_hd__a21o_1 _13238_ (.A1(_06264_),
    .A2(_06408_),
    .B1(_06307_),
    .X(_06409_));
 sky130_fd_sc_hd__and4_1 _13239_ (.A(_06308_),
    .B(_06310_),
    .C(_06367_),
    .D(_06381_),
    .X(_06410_));
 sky130_fd_sc_hd__nor2_1 _13240_ (.A(_06385_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__o21a_1 _13241_ (.A1(_06411_),
    .A2(_06388_),
    .B1(_06404_),
    .X(_06412_));
 sky130_fd_sc_hd__xnor2_1 _13242_ (.A(_06409_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__nor2_1 _13243_ (.A(net7837),
    .B(_06266_),
    .Y(_06414_));
 sky130_fd_sc_hd__o21a_1 _13244_ (.A1(_06263_),
    .A2(_06414_),
    .B1(_06306_),
    .X(_06415_));
 sky130_fd_sc_hd__and2_1 _13245_ (.A(_06303_),
    .B(_06304_),
    .X(_06416_));
 sky130_fd_sc_hd__a21oi_1 _13246_ (.A1(net8217),
    .A2(_06416_),
    .B1(_06415_),
    .Y(_06417_));
 sky130_fd_sc_hd__nor2_1 _13247_ (.A(_06387_),
    .B(_06409_),
    .Y(_06418_));
 sky130_fd_sc_hd__or2_1 _13248_ (.A(net8068),
    .B(_06266_),
    .X(_06419_));
 sky130_fd_sc_hd__a21o_1 _13249_ (.A1(_06264_),
    .A2(_06419_),
    .B1(_06307_),
    .X(_06420_));
 sky130_fd_sc_hd__o21a_1 _13250_ (.A1(net8275),
    .A2(_06266_),
    .B1(_06264_),
    .X(_06421_));
 sky130_fd_sc_hd__nor2_1 _13251_ (.A(_06420_),
    .B(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__a31o_1 _13252_ (.A1(_06410_),
    .A2(_06418_),
    .A3(_06422_),
    .B1(_06385_),
    .X(_06423_));
 sky130_fd_sc_hd__mux2_1 _13253_ (.A0(_06415_),
    .A1(_06417_),
    .S(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__and4b_1 _13254_ (.A_N(_06383_),
    .B(_06410_),
    .C(_06418_),
    .D(_06422_),
    .X(_06425_));
 sky130_fd_sc_hd__nand2_1 _13255_ (.A(_06414_),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__nor2_1 _13256_ (.A(_06307_),
    .B(_06421_),
    .Y(_06427_));
 sky130_fd_sc_hd__inv_2 _13257_ (.A(_06420_),
    .Y(_06428_));
 sky130_fd_sc_hd__a31o_1 _13258_ (.A1(_06410_),
    .A2(_06418_),
    .A3(_06428_),
    .B1(_06385_),
    .X(_06429_));
 sky130_fd_sc_hd__xnor2_2 _13259_ (.A(_06427_),
    .B(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__o21a_1 _13260_ (.A1(_06385_),
    .A2(_06418_),
    .B1(_06386_),
    .X(_06431_));
 sky130_fd_sc_hd__xnor2_2 _13261_ (.A(_06428_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__and4b_1 _13262_ (.A_N(_06424_),
    .B(_06426_),
    .C(_06430_),
    .D(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__or4bb_4 _13263_ (.A(_06389_),
    .B(_06407_),
    .C_N(_06413_),
    .D_N(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__buf_6 _13264_ (.A(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__buf_2 _13265_ (.A(net559),
    .X(_06436_));
 sky130_fd_sc_hd__nand2_2 _13266_ (.A(_06404_),
    .B(_06354_),
    .Y(_06437_));
 sky130_fd_sc_hd__xnor2_4 _13267_ (.A(_06319_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__a21o_1 _13268_ (.A1(net8217),
    .A2(_06314_),
    .B1(_06316_),
    .X(_06439_));
 sky130_fd_sc_hd__o21ai_2 _13269_ (.A1(_06354_),
    .A2(_06319_),
    .B1(_06404_),
    .Y(_06440_));
 sky130_fd_sc_hd__xnor2_4 _13270_ (.A(_06439_),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__or2_2 _13271_ (.A(_06438_),
    .B(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__and2_1 _13272_ (.A(_06335_),
    .B(_06337_),
    .X(_06443_));
 sky130_fd_sc_hd__nand2_1 _13273_ (.A(_06351_),
    .B(_06404_),
    .Y(_06444_));
 sky130_fd_sc_hd__xnor2_1 _13274_ (.A(_06443_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__and2_2 _13275_ (.A(_06404_),
    .B(_06353_),
    .X(_06446_));
 sky130_fd_sc_hd__xor2_4 _13276_ (.A(_06327_),
    .B(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__a21oi_2 _13277_ (.A1(net8217),
    .A2(_06321_),
    .B1(_06323_),
    .Y(_06448_));
 sky130_fd_sc_hd__o21a_1 _13278_ (.A1(_06353_),
    .A2(_06327_),
    .B1(_06404_),
    .X(_06449_));
 sky130_fd_sc_hd__xnor2_4 _13279_ (.A(_06448_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__o21ai_2 _13280_ (.A1(net8217),
    .A2(_06329_),
    .B1(_06332_),
    .Y(_06451_));
 sky130_fd_sc_hd__or2_2 _13281_ (.A(_06385_),
    .B(_06352_),
    .X(_06452_));
 sky130_fd_sc_hd__xnor2_2 _13282_ (.A(_06451_),
    .B(_06452_),
    .Y(_06453_));
 sky130_fd_sc_hd__or4_2 _13283_ (.A(_06445_),
    .B(_06447_),
    .C(_06450_),
    .D(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__or3_4 _13284_ (.A(_06435_),
    .B(_06442_),
    .C(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__a21o_2 _13285_ (.A1(_06306_),
    .A2(_06338_),
    .B1(_06341_),
    .X(_06456_));
 sky130_fd_sc_hd__nor2_1 _13286_ (.A(_06346_),
    .B(_06350_),
    .Y(_06457_));
 sky130_fd_sc_hd__nor2_2 _13287_ (.A(_06457_),
    .B(_06385_),
    .Y(_06458_));
 sky130_fd_sc_hd__xor2_4 _13288_ (.A(_06456_),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__and2_1 _13289_ (.A(_06346_),
    .B(_06404_),
    .X(_06460_));
 sky130_fd_sc_hd__xnor2_4 _13290_ (.A(_06350_),
    .B(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__xnor2_2 _13291_ (.A(_06327_),
    .B(_06446_),
    .Y(_06462_));
 sky130_fd_sc_hd__or4_4 _13292_ (.A(_06435_),
    .B(_06442_),
    .C(_06462_),
    .D(_06450_),
    .X(_06463_));
 sky130_fd_sc_hd__o31ai_4 _13293_ (.A1(_06455_),
    .A2(_06459_),
    .A3(_06461_),
    .B1(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__nor4_1 _13294_ (.A(_06351_),
    .B(_06435_),
    .C(_06442_),
    .D(_06454_),
    .Y(_06465_));
 sky130_fd_sc_hd__inv_2 _13295_ (.A(_06403_),
    .Y(_06466_));
 sky130_fd_sc_hd__buf_2 _13296_ (.A(_06413_),
    .X(_06467_));
 sky130_fd_sc_hd__nor2_1 _13297_ (.A(_06389_),
    .B(_06401_),
    .Y(_06468_));
 sky130_fd_sc_hd__and3_2 _13298_ (.A(_06467_),
    .B(_06433_),
    .C(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__xnor2_1 _13299_ (.A(_06365_),
    .B(_06405_),
    .Y(_06470_));
 sky130_fd_sc_hd__nor2_1 _13300_ (.A(_06399_),
    .B(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__inv_2 _13301_ (.A(_06438_),
    .Y(_06472_));
 sky130_fd_sc_hd__nor2_1 _13302_ (.A(_06398_),
    .B(_06403_),
    .Y(_06473_));
 sky130_fd_sc_hd__nor3_1 _13303_ (.A(net570),
    .B(_06406_),
    .C(_06441_),
    .Y(_06474_));
 sky130_fd_sc_hd__and4_1 _13304_ (.A(_06472_),
    .B(_06450_),
    .C(_06473_),
    .D(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__and4_1 _13305_ (.A(_06467_),
    .B(net574),
    .C(_06468_),
    .D(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__a31o_1 _13306_ (.A1(_06466_),
    .A2(_06469_),
    .A3(_06471_),
    .B1(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__xor2_1 _13307_ (.A(_06386_),
    .B(_06388_),
    .X(_06478_));
 sky130_fd_sc_hd__nor2_1 _13308_ (.A(_06438_),
    .B(_06454_),
    .Y(_06479_));
 sky130_fd_sc_hd__and2_1 _13309_ (.A(_06473_),
    .B(_06474_),
    .X(_06480_));
 sky130_fd_sc_hd__xor2_1 _13310_ (.A(_06378_),
    .B(_06393_),
    .X(_06481_));
 sky130_fd_sc_hd__a31o_1 _13311_ (.A1(_06392_),
    .A2(_06481_),
    .A3(_06473_),
    .B1(_06401_),
    .X(_06482_));
 sky130_fd_sc_hd__a31o_1 _13312_ (.A1(_06459_),
    .A2(_06479_),
    .A3(_06480_),
    .B1(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__and4_1 _13313_ (.A(_06478_),
    .B(_06467_),
    .C(net574),
    .D(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__and4_1 _13314_ (.A(_06467_),
    .B(_06433_),
    .C(_06403_),
    .D(_06468_),
    .X(_06485_));
 sky130_fd_sc_hd__nand2_1 _13315_ (.A(_06430_),
    .B(_06432_),
    .Y(_06486_));
 sky130_fd_sc_hd__and3b_1 _13316_ (.A_N(_06424_),
    .B(_06426_),
    .C(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__or2_1 _13317_ (.A(_06485_),
    .B(_06487_),
    .X(_06488_));
 sky130_fd_sc_hd__or4_2 _13318_ (.A(_06465_),
    .B(_06477_),
    .C(_06484_),
    .D(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__nor2_1 _13319_ (.A(net82),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__buf_6 _13320_ (.A(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__buf_6 _13321_ (.A(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__buf_4 _13322_ (.A(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__clkbuf_1 _13323_ (.A(net7810),
    .X(_06494_));
 sky130_fd_sc_hd__or4_4 _13324_ (.A(_06351_),
    .B(_06434_),
    .C(_06442_),
    .D(_06454_),
    .X(_06495_));
 sky130_fd_sc_hd__inv_2 _13325_ (.A(_06343_),
    .Y(_06496_));
 sky130_fd_sc_hd__nand2_2 _13326_ (.A(_06343_),
    .B(_06404_),
    .Y(_06497_));
 sky130_fd_sc_hd__xnor2_4 _13327_ (.A(_06345_),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__xnor2_1 _13328_ (.A(_06456_),
    .B(_06458_),
    .Y(_06499_));
 sky130_fd_sc_hd__nand2_1 _13329_ (.A(_06499_),
    .B(_06461_),
    .Y(_06500_));
 sky130_fd_sc_hd__or3_1 _13330_ (.A(_06496_),
    .B(_06498_),
    .C(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__or4_4 _13331_ (.A(_06434_),
    .B(_06442_),
    .C(_06454_),
    .D(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__nand2_4 _13332_ (.A(_06495_),
    .B(net554),
    .Y(_06503_));
 sky130_fd_sc_hd__and4b_1 _13333_ (.A_N(_06407_),
    .B(_06467_),
    .C(_06478_),
    .D(_06433_),
    .X(_06504_));
 sky130_fd_sc_hd__clkbuf_4 _13334_ (.A(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__nor2_1 _13335_ (.A(_06472_),
    .B(_06441_),
    .Y(_06506_));
 sky130_fd_sc_hd__and2_1 _13336_ (.A(_06468_),
    .B(_06473_),
    .X(_06507_));
 sky130_fd_sc_hd__and3b_1 _13337_ (.A_N(net570),
    .B(_06470_),
    .C(_06441_),
    .X(_06508_));
 sky130_fd_sc_hd__and4_1 _13338_ (.A(_06467_),
    .B(net574),
    .C(_06507_),
    .D(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__a21oi_1 _13339_ (.A1(_06505_),
    .A2(_06506_),
    .B1(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__nand2_4 _13340_ (.A(_06463_),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__and4b_1 _13341_ (.A_N(_06500_),
    .B(_06507_),
    .C(_06474_),
    .D(_06498_),
    .X(_06512_));
 sky130_fd_sc_hd__nand2_1 _13342_ (.A(_06467_),
    .B(_06468_),
    .Y(_06513_));
 sky130_fd_sc_hd__a211o_1 _13343_ (.A1(_06479_),
    .A2(_06512_),
    .B1(_06475_),
    .C1(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__a21o_1 _13344_ (.A1(net574),
    .A2(_06514_),
    .B1(_06485_),
    .X(_06515_));
 sky130_fd_sc_hd__nor3_4 _13345_ (.A(_06503_),
    .B(_06511_),
    .C(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__and4bb_1 _13346_ (.A_N(_06424_),
    .B_N(_06432_),
    .C(_06426_),
    .D(_06430_),
    .X(_06517_));
 sky130_fd_sc_hd__a311o_1 _13347_ (.A1(_06389_),
    .A2(_06467_),
    .A3(_06433_),
    .B1(_06517_),
    .C1(_06424_),
    .X(_06518_));
 sky130_fd_sc_hd__a211o_1 _13348_ (.A1(_06505_),
    .A2(_06506_),
    .B1(_06485_),
    .C1(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__nor2_1 _13349_ (.A(_06481_),
    .B(_06398_),
    .Y(_06520_));
 sky130_fd_sc_hd__o211a_1 _13350_ (.A1(_06471_),
    .A2(_06520_),
    .B1(_06466_),
    .C1(_06469_),
    .X(_06521_));
 sky130_fd_sc_hd__xor2_2 _13351_ (.A(_06443_),
    .B(_06444_),
    .X(_06522_));
 sky130_fd_sc_hd__or4_1 _13352_ (.A(_06522_),
    .B(_06447_),
    .C(_06450_),
    .D(_06453_),
    .X(_06523_));
 sky130_fd_sc_hd__or3_1 _13353_ (.A(_06435_),
    .B(_06442_),
    .C(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__or4bb_4 _13354_ (.A(_06519_),
    .B(_06521_),
    .C_N(net554),
    .D_N(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__a21o_1 _13355_ (.A1(_06489_),
    .A2(_06525_),
    .B1(net82),
    .X(_06526_));
 sky130_fd_sc_hd__xnor2_1 _13356_ (.A(_06516_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__nor2_2 _13357_ (.A(net82),
    .B(_06525_),
    .Y(_06528_));
 sky130_fd_sc_hd__xnor2_4 _13358_ (.A(_06491_),
    .B(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__o31a_1 _13359_ (.A1(_06455_),
    .A2(_06459_),
    .A3(_06461_),
    .B1(_06463_),
    .X(_06530_));
 sky130_fd_sc_hd__buf_6 _13360_ (.A(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__and4bb_2 _13361_ (.A_N(_06519_),
    .B_N(_06521_),
    .C(_06502_),
    .D(_06524_),
    .X(_06532_));
 sky130_fd_sc_hd__buf_6 _13362_ (.A(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__a21oi_1 _13363_ (.A1(net561),
    .A2(net560),
    .B1(_06498_),
    .Y(_06534_));
 sky130_fd_sc_hd__a21oi_1 _13364_ (.A1(_06496_),
    .A2(_06528_),
    .B1(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__and3_1 _13365_ (.A(_06527_),
    .B(_06529_),
    .C(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__or3_1 _13366_ (.A(_06503_),
    .B(_06511_),
    .C(_06515_),
    .X(_06537_));
 sky130_fd_sc_hd__clkbuf_4 _13367_ (.A(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__a311oi_4 _13368_ (.A1(_06399_),
    .A2(_06466_),
    .A3(_06469_),
    .B1(_06477_),
    .C1(_06511_),
    .Y(_06539_));
 sky130_fd_sc_hd__xnor2_4 _13369_ (.A(_06538_),
    .B(net81),
    .Y(_06540_));
 sky130_fd_sc_hd__and2_1 _13370_ (.A(_06516_),
    .B(net562),
    .X(_06541_));
 sky130_fd_sc_hd__nand3_2 _13371_ (.A(_06466_),
    .B(_06469_),
    .C(_06471_),
    .Y(_06542_));
 sky130_fd_sc_hd__o21ai_4 _13372_ (.A1(_06540_),
    .A2(_06541_),
    .B1(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__nor2_2 _13373_ (.A(net7833),
    .B(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__o21a_2 _13374_ (.A1(_06540_),
    .A2(_06541_),
    .B1(_06542_),
    .X(_06545_));
 sky130_fd_sc_hd__nor2_2 _13375_ (.A(net559),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__clkbuf_4 _13376_ (.A(_06527_),
    .X(_06547_));
 sky130_fd_sc_hd__xor2_1 _13377_ (.A(_06451_),
    .B(_06452_),
    .X(_06548_));
 sky130_fd_sc_hd__nand2_4 _13378_ (.A(_06531_),
    .B(_06533_),
    .Y(_06549_));
 sky130_fd_sc_hd__or2_2 _13379_ (.A(net82),
    .B(_06489_),
    .X(_06550_));
 sky130_fd_sc_hd__buf_6 _13380_ (.A(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__mux4_2 _13381_ (.A0(_06522_),
    .A1(_06499_),
    .A2(_06461_),
    .A3(_06548_),
    .S0(_06549_),
    .S1(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__clkbuf_2 _13382_ (.A(_06549_),
    .X(_06553_));
 sky130_fd_sc_hd__mux4_1 _13383_ (.A0(_06438_),
    .A1(_06447_),
    .A2(_06450_),
    .A3(_06441_),
    .S0(_06551_),
    .S1(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__nand2_1 _13384_ (.A(_06547_),
    .B(_06554_),
    .Y(_06555_));
 sky130_fd_sc_hd__o21ai_2 _13385_ (.A1(_06547_),
    .A2(_06552_),
    .B1(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__buf_2 _13386_ (.A(_06538_),
    .X(_06557_));
 sky130_fd_sc_hd__buf_2 _13387_ (.A(_06528_),
    .X(_06558_));
 sky130_fd_sc_hd__or3_1 _13388_ (.A(_06406_),
    .B(_06464_),
    .C(_06525_),
    .X(_06559_));
 sky130_fd_sc_hd__o211a_1 _13389_ (.A1(_06441_),
    .A2(_06558_),
    .B1(_06559_),
    .C1(_06550_),
    .X(_06560_));
 sky130_fd_sc_hd__or3_1 _13390_ (.A(_06394_),
    .B(net82),
    .C(_06525_),
    .X(_06561_));
 sky130_fd_sc_hd__o211a_1 _13391_ (.A1(_06392_),
    .A2(_06558_),
    .B1(_06561_),
    .C1(_06491_),
    .X(_06562_));
 sky130_fd_sc_hd__or3_1 _13392_ (.A(_06557_),
    .B(_06560_),
    .C(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__buf_2 _13393_ (.A(_06516_),
    .X(_06564_));
 sky130_fd_sc_hd__mux2_1 _13394_ (.A0(_06389_),
    .A1(_06401_),
    .S(_06549_),
    .X(_06565_));
 sky130_fd_sc_hd__mux2_1 _13395_ (.A0(_06398_),
    .A1(_06403_),
    .S(_06528_),
    .X(_06566_));
 sky130_fd_sc_hd__mux2_1 _13396_ (.A0(_06565_),
    .A1(_06566_),
    .S(_06551_),
    .X(_06567_));
 sky130_fd_sc_hd__nand2_2 _13397_ (.A(_06516_),
    .B(_06539_),
    .Y(_06568_));
 sky130_fd_sc_hd__o21a_1 _13398_ (.A1(_06564_),
    .A2(_06567_),
    .B1(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__nor2_1 _13399_ (.A(_06430_),
    .B(_06551_),
    .Y(_06570_));
 sky130_fd_sc_hd__buf_2 _13400_ (.A(_06528_),
    .X(_06571_));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(_06467_),
    .A1(_06432_),
    .S(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__nor2_1 _13402_ (.A(_06493_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__a211o_1 _13403_ (.A1(_06563_),
    .A2(_06569_),
    .B1(_06570_),
    .C1(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__a221oi_4 _13404_ (.A1(net73),
    .A2(_06544_),
    .B1(_06546_),
    .B2(_06556_),
    .C1(_06574_),
    .Y(_06575_));
 sky130_fd_sc_hd__clkbuf_4 _13405_ (.A(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__inv_2 _13406_ (.A(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__a21oi_1 _13407_ (.A1(net561),
    .A2(net560),
    .B1(_06453_),
    .Y(_06578_));
 sky130_fd_sc_hd__a211o_1 _13408_ (.A1(_06462_),
    .A2(_06558_),
    .B1(_06578_),
    .C1(_06491_),
    .X(_06579_));
 sky130_fd_sc_hd__a21oi_1 _13409_ (.A1(_06531_),
    .A2(_06533_),
    .B1(_06450_),
    .Y(_06580_));
 sky130_fd_sc_hd__a211o_1 _13410_ (.A1(_06472_),
    .A2(_06558_),
    .B1(_06580_),
    .C1(_06550_),
    .X(_06581_));
 sky130_fd_sc_hd__a21o_1 _13411_ (.A1(_06579_),
    .A2(_06581_),
    .B1(_06516_),
    .X(_06582_));
 sky130_fd_sc_hd__a211o_1 _13412_ (.A1(_06461_),
    .A2(_06558_),
    .B1(_06534_),
    .C1(_06491_),
    .X(_06583_));
 sky130_fd_sc_hd__and3_1 _13413_ (.A(_06522_),
    .B(_06531_),
    .C(_06533_),
    .X(_06584_));
 sky130_fd_sc_hd__a21oi_1 _13414_ (.A1(net561),
    .A2(net560),
    .B1(_06459_),
    .Y(_06585_));
 sky130_fd_sc_hd__or3_4 _13415_ (.A(_06550_),
    .B(_06584_),
    .C(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__a21o_1 _13416_ (.A1(_06583_),
    .A2(_06586_),
    .B1(_06538_),
    .X(_06587_));
 sky130_fd_sc_hd__o31ai_1 _13417_ (.A1(_06568_),
    .A2(_06560_),
    .A3(_06562_),
    .B1(net559),
    .Y(_06588_));
 sky130_fd_sc_hd__a31o_4 _13418_ (.A1(_06540_),
    .A2(_06582_),
    .A3(_06587_),
    .B1(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__or3b_4 _13419_ (.A(_06435_),
    .B(_06545_),
    .C_N(_06536_),
    .X(_06590_));
 sky130_fd_sc_hd__a21oi_1 _13420_ (.A1(net561),
    .A2(net560),
    .B1(_06496_),
    .Y(_06591_));
 sky130_fd_sc_hd__a211o_1 _13421_ (.A1(_06498_),
    .A2(_06571_),
    .B1(_06591_),
    .C1(_06492_),
    .X(_06592_));
 sky130_fd_sc_hd__and3_1 _13422_ (.A(_06459_),
    .B(_06463_),
    .C(_06532_),
    .X(_06593_));
 sky130_fd_sc_hd__a21oi_1 _13423_ (.A1(_06530_),
    .A2(_06532_),
    .B1(_06461_),
    .Y(_06594_));
 sky130_fd_sc_hd__or3_1 _13424_ (.A(_06550_),
    .B(_06593_),
    .C(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__a21o_1 _13425_ (.A1(_06592_),
    .A2(_06595_),
    .B1(_06557_),
    .X(_06596_));
 sky130_fd_sc_hd__or3_1 _13426_ (.A(_06450_),
    .B(net82),
    .C(_06525_),
    .X(_06597_));
 sky130_fd_sc_hd__a21o_1 _13427_ (.A1(_06531_),
    .A2(_06533_),
    .B1(_06447_),
    .X(_06598_));
 sky130_fd_sc_hd__and3_1 _13428_ (.A(_06491_),
    .B(_06597_),
    .C(_06598_),
    .X(_06599_));
 sky130_fd_sc_hd__a21o_1 _13429_ (.A1(_06530_),
    .A2(_06532_),
    .B1(_06522_),
    .X(_06600_));
 sky130_fd_sc_hd__or3_1 _13430_ (.A(_06548_),
    .B(_06464_),
    .C(_06525_),
    .X(_06601_));
 sky130_fd_sc_hd__a21oi_1 _13431_ (.A1(_06600_),
    .A2(_06601_),
    .B1(_06492_),
    .Y(_06602_));
 sky130_fd_sc_hd__or3_1 _13432_ (.A(_06516_),
    .B(_06599_),
    .C(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__or2_1 _13433_ (.A(_06516_),
    .B(_06539_),
    .X(_06604_));
 sky130_fd_sc_hd__nand2_1 _13434_ (.A(_06568_),
    .B(_06604_),
    .Y(_06605_));
 sky130_fd_sc_hd__clkbuf_2 _13435_ (.A(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__a21oi_2 _13436_ (.A1(_06596_),
    .A2(_06603_),
    .B1(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__mux2_1 _13437_ (.A0(_06401_),
    .A1(_06403_),
    .S(_06549_),
    .X(_06608_));
 sky130_fd_sc_hd__or3_1 _13438_ (.A(_06398_),
    .B(net82),
    .C(_06525_),
    .X(_06609_));
 sky130_fd_sc_hd__o211a_1 _13439_ (.A1(_06394_),
    .A2(_06558_),
    .B1(_06609_),
    .C1(_06550_),
    .X(_06610_));
 sky130_fd_sc_hd__a211o_1 _13440_ (.A1(_06492_),
    .A2(_06608_),
    .B1(_06610_),
    .C1(_06564_),
    .X(_06611_));
 sky130_fd_sc_hd__or3_1 _13441_ (.A(_06392_),
    .B(net82),
    .C(_06525_),
    .X(_06612_));
 sky130_fd_sc_hd__a21o_1 _13442_ (.A1(net561),
    .A2(net560),
    .B1(_06406_),
    .X(_06613_));
 sky130_fd_sc_hd__a21o_1 _13443_ (.A1(_06531_),
    .A2(_06533_),
    .B1(_06438_),
    .X(_06614_));
 sky130_fd_sc_hd__o211a_1 _13444_ (.A1(_06441_),
    .A2(_06549_),
    .B1(_06614_),
    .C1(_06550_),
    .X(_06615_));
 sky130_fd_sc_hd__a311o_1 _13445_ (.A1(_06492_),
    .A2(_06612_),
    .A3(_06613_),
    .B1(_06615_),
    .C1(_06538_),
    .X(_06616_));
 sky130_fd_sc_hd__a21oi_2 _13446_ (.A1(_06611_),
    .A2(_06616_),
    .B1(_06540_),
    .Y(_06617_));
 sky130_fd_sc_hd__a211o_4 _13447_ (.A1(_06589_),
    .A2(_06590_),
    .B1(_06607_),
    .C1(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__o211a_1 _13448_ (.A1(_06441_),
    .A2(_06549_),
    .B1(_06614_),
    .C1(_06491_),
    .X(_06619_));
 sky130_fd_sc_hd__a31oi_2 _13449_ (.A1(_06551_),
    .A2(_06597_),
    .A3(_06598_),
    .B1(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__and3_1 _13450_ (.A(_06491_),
    .B(_06600_),
    .C(_06601_),
    .X(_06621_));
 sky130_fd_sc_hd__or3_1 _13451_ (.A(_06490_),
    .B(_06593_),
    .C(_06594_),
    .X(_06622_));
 sky130_fd_sc_hd__or3b_1 _13452_ (.A(_06538_),
    .B(_06621_),
    .C_N(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__o211a_1 _13453_ (.A1(_06564_),
    .A2(_06620_),
    .B1(_06623_),
    .C1(_06540_),
    .X(_06624_));
 sky130_fd_sc_hd__o21a_1 _13454_ (.A1(_06394_),
    .A2(_06528_),
    .B1(_06609_),
    .X(_06625_));
 sky130_fd_sc_hd__and3_1 _13455_ (.A(_06550_),
    .B(_06612_),
    .C(_06613_),
    .X(_06626_));
 sky130_fd_sc_hd__a21oi_1 _13456_ (.A1(_06492_),
    .A2(_06625_),
    .B1(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__a21o_1 _13457_ (.A1(_06564_),
    .A2(_06627_),
    .B1(_06505_),
    .X(_06628_));
 sky130_fd_sc_hd__a21o_1 _13458_ (.A1(_06498_),
    .A2(_06558_),
    .B1(_06594_),
    .X(_06629_));
 sky130_fd_sc_hd__a22o_1 _13459_ (.A1(_06492_),
    .A2(_06591_),
    .B1(_06629_),
    .B2(_06529_),
    .X(_06630_));
 sky130_fd_sc_hd__nand2_1 _13460_ (.A(_06547_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_2 _13461_ (.A(_06505_),
    .B(_06543_),
    .Y(_06632_));
 sky130_fd_sc_hd__o22a_1 _13462_ (.A1(_06624_),
    .A2(_06628_),
    .B1(_06631_),
    .B2(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__clkbuf_8 _13463_ (.A(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__a311o_1 _13464_ (.A1(_06492_),
    .A2(_06612_),
    .A3(_06613_),
    .B1(_06615_),
    .C1(_06564_),
    .X(_06635_));
 sky130_fd_sc_hd__or3_1 _13465_ (.A(_06538_),
    .B(_06599_),
    .C(_06602_),
    .X(_06636_));
 sky130_fd_sc_hd__a21o_1 _13466_ (.A1(_06635_),
    .A2(_06636_),
    .B1(_06606_),
    .X(_06637_));
 sky130_fd_sc_hd__a211o_1 _13467_ (.A1(_06493_),
    .A2(_06608_),
    .B1(_06610_),
    .C1(_06568_),
    .X(_06638_));
 sky130_fd_sc_hd__inv_2 _13468_ (.A(_06461_),
    .Y(_06639_));
 sky130_fd_sc_hd__mux4_1 _13469_ (.A0(_06445_),
    .A1(_06498_),
    .A2(_06639_),
    .A3(_06459_),
    .S0(_06528_),
    .S1(_06491_),
    .X(_06640_));
 sky130_fd_sc_hd__a32o_1 _13470_ (.A1(_06538_),
    .A2(_06551_),
    .A3(_06591_),
    .B1(_06640_),
    .B2(_06527_),
    .X(_06641_));
 sky130_fd_sc_hd__and2_1 _13471_ (.A(_06505_),
    .B(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__a31oi_2 _13472_ (.A1(_06436_),
    .A2(_06637_),
    .A3(_06638_),
    .B1(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__mux4_2 _13473_ (.A0(_06343_),
    .A1(_06459_),
    .A2(_06639_),
    .A3(_06498_),
    .S0(_06549_),
    .S1(_06492_),
    .X(_06644_));
 sky130_fd_sc_hd__o21a_1 _13474_ (.A1(_06441_),
    .A2(_06558_),
    .B1(_06559_),
    .X(_06645_));
 sky130_fd_sc_hd__a21oi_1 _13475_ (.A1(_06472_),
    .A2(_06558_),
    .B1(_06580_),
    .Y(_06646_));
 sky130_fd_sc_hd__mux2_1 _13476_ (.A0(_06645_),
    .A1(_06646_),
    .S(_06551_),
    .X(_06647_));
 sky130_fd_sc_hd__a211o_1 _13477_ (.A1(_06462_),
    .A2(_06571_),
    .B1(_06578_),
    .C1(_06551_),
    .X(_06648_));
 sky130_fd_sc_hd__or3_1 _13478_ (.A(_06491_),
    .B(_06584_),
    .C(_06585_),
    .X(_06649_));
 sky130_fd_sc_hd__a21oi_1 _13479_ (.A1(_06648_),
    .A2(_06649_),
    .B1(_06538_),
    .Y(_06650_));
 sky130_fd_sc_hd__a211o_1 _13480_ (.A1(_06557_),
    .A2(_06647_),
    .B1(_06650_),
    .C1(_06605_),
    .X(_06651_));
 sky130_fd_sc_hd__o21a_1 _13481_ (.A1(_06392_),
    .A2(_06558_),
    .B1(_06561_),
    .X(_06652_));
 sky130_fd_sc_hd__mux2_1 _13482_ (.A0(_06652_),
    .A1(_06566_),
    .S(_06492_),
    .X(_06653_));
 sky130_fd_sc_hd__o21a_1 _13483_ (.A1(_06568_),
    .A2(_06653_),
    .B1(net559),
    .X(_06654_));
 sky130_fd_sc_hd__a32oi_4 _13484_ (.A1(_06547_),
    .A2(_06546_),
    .A3(_06644_),
    .B1(_06651_),
    .B2(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__or3_1 _13485_ (.A(_06564_),
    .B(_06560_),
    .C(_06562_),
    .X(_06656_));
 sky130_fd_sc_hd__nand3_1 _13486_ (.A(_06564_),
    .B(_06579_),
    .C(_06581_),
    .Y(_06657_));
 sky130_fd_sc_hd__a21o_1 _13487_ (.A1(_06656_),
    .A2(_06657_),
    .B1(_06606_),
    .X(_06658_));
 sky130_fd_sc_hd__o21a_1 _13488_ (.A1(_06568_),
    .A2(_06567_),
    .B1(net559),
    .X(_06659_));
 sky130_fd_sc_hd__nand2_1 _13489_ (.A(_06529_),
    .B(_06535_),
    .Y(_06660_));
 sky130_fd_sc_hd__mux2_1 _13490_ (.A0(_06660_),
    .A1(_06552_),
    .S(_06547_),
    .X(_06661_));
 sky130_fd_sc_hd__o2bb2a_2 _13491_ (.A1_N(_06658_),
    .A2_N(_06659_),
    .B1(_06632_),
    .B2(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__a2111o_4 _13492_ (.A1(_06618_),
    .A2(_06634_),
    .B1(net79),
    .C1(net80),
    .D1(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__mux4_1 _13493_ (.A0(_06522_),
    .A1(_06462_),
    .A2(_06548_),
    .A3(_06499_),
    .S0(_06551_),
    .S1(_06571_),
    .X(_06664_));
 sky130_fd_sc_hd__o211a_1 _13494_ (.A1(_06547_),
    .A2(_06630_),
    .B1(_06543_),
    .C1(_06505_),
    .X(_06665_));
 sky130_fd_sc_hd__a21bo_1 _13495_ (.A1(_06547_),
    .A2(_06664_),
    .B1_N(_06665_),
    .X(_06666_));
 sky130_fd_sc_hd__mux2_1 _13496_ (.A0(_06620_),
    .A1(_06627_),
    .S(_06557_),
    .X(_06667_));
 sky130_fd_sc_hd__or2_1 _13497_ (.A(_06606_),
    .B(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__mux2_1 _13498_ (.A0(_06478_),
    .A1(_06467_),
    .S(_06571_),
    .X(_06669_));
 sky130_fd_sc_hd__nor2_1 _13499_ (.A(_06493_),
    .B(_06608_),
    .Y(_06670_));
 sky130_fd_sc_hd__a211o_1 _13500_ (.A1(_06493_),
    .A2(_06669_),
    .B1(_06670_),
    .C1(_06557_),
    .X(_06671_));
 sky130_fd_sc_hd__and3_1 _13501_ (.A(_06666_),
    .B(_06668_),
    .C(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__buf_4 _13502_ (.A(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__mux4_1 _13503_ (.A0(_06445_),
    .A1(_06447_),
    .A2(_06450_),
    .A3(_06453_),
    .S0(_06493_),
    .S1(_06553_),
    .X(_06674_));
 sky130_fd_sc_hd__mux2_1 _13504_ (.A0(_06644_),
    .A1(_06674_),
    .S(_06547_),
    .X(_06675_));
 sky130_fd_sc_hd__buf_1 _13505_ (.A(_06540_),
    .X(_06676_));
 sky130_fd_sc_hd__mux2_1 _13506_ (.A0(_06647_),
    .A1(_06653_),
    .S(_06557_),
    .X(_06677_));
 sky130_fd_sc_hd__nand2_1 _13507_ (.A(_06493_),
    .B(_06572_),
    .Y(_06678_));
 sky130_fd_sc_hd__o21ai_1 _13508_ (.A1(_06493_),
    .A2(_06565_),
    .B1(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__a21bo_1 _13509_ (.A1(_06676_),
    .A2(_06677_),
    .B1_N(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__a21o_1 _13510_ (.A1(_06546_),
    .A2(_06675_),
    .B1(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__a21bo_1 _13511_ (.A1(_06663_),
    .A2(_06673_),
    .B1_N(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__buf_6 _13512_ (.A(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__nand3_1 _13513_ (.A(_06676_),
    .B(_06611_),
    .C(_06616_),
    .Y(_06684_));
 sky130_fd_sc_hd__mux2_1 _13514_ (.A0(_06430_),
    .A1(_06432_),
    .S(_06553_),
    .X(_06685_));
 sky130_fd_sc_hd__mux2_1 _13515_ (.A0(_06669_),
    .A1(_06685_),
    .S(_06493_),
    .X(_06686_));
 sky130_fd_sc_hd__nand2_1 _13516_ (.A(_06505_),
    .B(_06545_),
    .Y(_06687_));
 sky130_fd_sc_hd__and3_1 _13517_ (.A(_06343_),
    .B(_06564_),
    .C(net562),
    .X(_06688_));
 sky130_fd_sc_hd__mux4_1 _13518_ (.A0(_06438_),
    .A1(_06447_),
    .A2(_06453_),
    .A3(_06450_),
    .S0(_06493_),
    .S1(_06571_),
    .X(_06689_));
 sky130_fd_sc_hd__mux2_1 _13519_ (.A0(_06640_),
    .A1(_06689_),
    .S(_06547_),
    .X(_06690_));
 sky130_fd_sc_hd__o22ai_1 _13520_ (.A1(_06687_),
    .A2(_06688_),
    .B1(_06690_),
    .B2(_06632_),
    .Y(_06691_));
 sky130_fd_sc_hd__a31o_4 _13521_ (.A1(_06436_),
    .A2(_06684_),
    .A3(_06686_),
    .B1(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__buf_2 _13522_ (.A(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__nor2_8 _13523_ (.A(_06683_),
    .B(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__a21o_2 _13524_ (.A1(_06577_),
    .A2(_06694_),
    .B1(net83),
    .X(_06695_));
 sky130_fd_sc_hd__clkbuf_4 _13525_ (.A(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__xnor2_4 _13526_ (.A(_06576_),
    .B(_06694_),
    .Y(_06697_));
 sky130_fd_sc_hd__buf_2 _13527_ (.A(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__buf_2 _13528_ (.A(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__or2_1 _13529_ (.A(_06607_),
    .B(_06617_),
    .X(_06700_));
 sky130_fd_sc_hd__buf_2 _13530_ (.A(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__buf_2 _13531_ (.A(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_4 _13532_ (.A(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__and2_1 _13533_ (.A(_06589_),
    .B(_06590_),
    .X(_06704_));
 sky130_fd_sc_hd__clkbuf_4 _13534_ (.A(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__clkbuf_4 _13535_ (.A(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__or4_4 _13536_ (.A(_06703_),
    .B(_06706_),
    .C(_06697_),
    .D(_06695_),
    .X(_06707_));
 sky130_fd_sc_hd__clkbuf_4 _13537_ (.A(_06634_),
    .X(_06708_));
 sky130_fd_sc_hd__nor2_1 _13538_ (.A(_06708_),
    .B(_06697_),
    .Y(_06709_));
 sky130_fd_sc_hd__nor2_1 _13539_ (.A(_06706_),
    .B(_06695_),
    .Y(_06710_));
 sky130_fd_sc_hd__xnor2_1 _13540_ (.A(_06709_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__nor2_1 _13541_ (.A(_06707_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__nand2_1 _13542_ (.A(_06709_),
    .B(_06710_),
    .Y(_06713_));
 sky130_fd_sc_hd__or2_1 _13543_ (.A(_06708_),
    .B(_06695_),
    .X(_06714_));
 sky130_fd_sc_hd__buf_2 _13544_ (.A(net80),
    .X(_06715_));
 sky130_fd_sc_hd__nor2_1 _13545_ (.A(_06715_),
    .B(_06697_),
    .Y(_06716_));
 sky130_fd_sc_hd__xnor2_1 _13546_ (.A(_06714_),
    .B(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__xnor2_1 _13547_ (.A(_06713_),
    .B(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__clkbuf_4 _13548_ (.A(_06662_),
    .X(_06719_));
 sky130_fd_sc_hd__a211o_2 _13549_ (.A1(net567),
    .A2(_06634_),
    .B1(net79),
    .C1(net80),
    .X(_06720_));
 sky130_fd_sc_hd__nor2_2 _13550_ (.A(_06719_),
    .B(_06720_),
    .Y(_06721_));
 sky130_fd_sc_hd__a211oi_4 _13551_ (.A1(_06589_),
    .A2(_06590_),
    .B1(_06607_),
    .C1(_06617_),
    .Y(_06722_));
 sky130_fd_sc_hd__nand2_1 _13552_ (.A(net80),
    .B(_06634_),
    .Y(_06723_));
 sky130_fd_sc_hd__a21o_4 _13553_ (.A1(_06618_),
    .A2(_06634_),
    .B1(net80),
    .X(_06724_));
 sky130_fd_sc_hd__o21ai_4 _13554_ (.A1(_06722_),
    .A2(_06723_),
    .B1(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__xnor2_4 _13555_ (.A(_06724_),
    .B(net576),
    .Y(_06726_));
 sky130_fd_sc_hd__nand3_4 _13556_ (.A(_06666_),
    .B(_06668_),
    .C(_06671_),
    .Y(_06727_));
 sky130_fd_sc_hd__a22o_1 _13557_ (.A1(_06681_),
    .A2(_06725_),
    .B1(_06726_),
    .B2(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_4 _13558_ (.A(net555),
    .X(_06729_));
 sky130_fd_sc_hd__nand4_1 _13559_ (.A(_06729_),
    .B(_06727_),
    .C(_06725_),
    .D(_06726_),
    .Y(_06730_));
 sky130_fd_sc_hd__a21boi_1 _13560_ (.A1(_06721_),
    .A2(_06728_),
    .B1_N(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__xor2_2 _13561_ (.A(_06683_),
    .B(_06692_),
    .X(_06732_));
 sky130_fd_sc_hd__nor2_1 _13562_ (.A(net80),
    .B(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__xnor2_4 _13563_ (.A(_06663_),
    .B(_06673_),
    .Y(_06734_));
 sky130_fd_sc_hd__nor2_1 _13564_ (.A(_06719_),
    .B(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__or3b_4 _13565_ (.A(_06681_),
    .B(_06727_),
    .C_N(_06663_),
    .X(_06736_));
 sky130_fd_sc_hd__buf_4 _13566_ (.A(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__a21oi_1 _13567_ (.A1(_06683_),
    .A2(_06737_),
    .B1(net79),
    .Y(_06738_));
 sky130_fd_sc_hd__xnor2_1 _13568_ (.A(_06735_),
    .B(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__xnor2_1 _13569_ (.A(_06733_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__and2b_1 _13570_ (.A_N(_06731_),
    .B(_06740_),
    .X(_06741_));
 sky130_fd_sc_hd__nor2_1 _13571_ (.A(net79),
    .B(_06734_),
    .Y(_06742_));
 sky130_fd_sc_hd__a21oi_1 _13572_ (.A1(_06683_),
    .A2(_06737_),
    .B1(net80),
    .Y(_06743_));
 sky130_fd_sc_hd__or2_4 _13573_ (.A(_06634_),
    .B(_06732_),
    .X(_06744_));
 sky130_fd_sc_hd__xnor2_2 _13574_ (.A(_06742_),
    .B(_06743_),
    .Y(_06745_));
 sky130_fd_sc_hd__nor2_1 _13575_ (.A(net582),
    .B(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__a21o_1 _13576_ (.A1(_06742_),
    .A2(_06743_),
    .B1(_06746_),
    .X(_06747_));
 sky130_fd_sc_hd__xnor2_1 _13577_ (.A(_06731_),
    .B(_06740_),
    .Y(_06748_));
 sky130_fd_sc_hd__and2_1 _13578_ (.A(_06747_),
    .B(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__or3_1 _13579_ (.A(_06718_),
    .B(_06741_),
    .C(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__o21a_1 _13580_ (.A1(_06741_),
    .A2(_06749_),
    .B1(_06718_),
    .X(_06751_));
 sky130_fd_sc_hd__a21o_1 _13581_ (.A1(_06712_),
    .A2(_06750_),
    .B1(_06751_),
    .X(_06752_));
 sky130_fd_sc_hd__xor2_1 _13582_ (.A(_06701_),
    .B(_06705_),
    .X(_06753_));
 sky130_fd_sc_hd__clkbuf_4 _13583_ (.A(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__xnor2_4 _13584_ (.A(_06618_),
    .B(_06634_),
    .Y(_06755_));
 sky130_fd_sc_hd__or4_2 _13585_ (.A(net83),
    .B(_06576_),
    .C(_06754_),
    .D(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__buf_2 _13586_ (.A(_06495_),
    .X(_06757_));
 sky130_fd_sc_hd__xnor2_4 _13587_ (.A(_06701_),
    .B(_06705_),
    .Y(_06758_));
 sky130_fd_sc_hd__xnor2_4 _13588_ (.A(net78),
    .B(_06634_),
    .Y(_06759_));
 sky130_fd_sc_hd__a22o_1 _13589_ (.A1(_06757_),
    .A2(_06758_),
    .B1(_06759_),
    .B2(_06577_),
    .X(_06760_));
 sky130_fd_sc_hd__nand2_1 _13590_ (.A(_06756_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__or3_1 _13591_ (.A(_06575_),
    .B(_06702_),
    .C(_06754_),
    .X(_06762_));
 sky130_fd_sc_hd__nor2_1 _13592_ (.A(_06692_),
    .B(_06755_),
    .Y(_06763_));
 sky130_fd_sc_hd__o21ai_1 _13593_ (.A1(_06576_),
    .A2(_06754_),
    .B1(_06702_),
    .Y(_06764_));
 sky130_fd_sc_hd__nand3_1 _13594_ (.A(_06762_),
    .B(_06763_),
    .C(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__nand2_1 _13595_ (.A(_06762_),
    .B(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__xor2_1 _13596_ (.A(_06761_),
    .B(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__inv_2 _13597_ (.A(_06662_),
    .Y(_06768_));
 sky130_fd_sc_hd__xnor2_2 _13598_ (.A(_06768_),
    .B(_06720_),
    .Y(_06769_));
 sky130_fd_sc_hd__or2_1 _13599_ (.A(_06673_),
    .B(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__o21a_2 _13600_ (.A1(_06722_),
    .A2(_06723_),
    .B1(_06724_),
    .X(_06771_));
 sky130_fd_sc_hd__or2_1 _13601_ (.A(_06693_),
    .B(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__nand2_1 _13602_ (.A(_06729_),
    .B(_06726_),
    .Y(_06773_));
 sky130_fd_sc_hd__xor2_1 _13603_ (.A(_06772_),
    .B(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__xnor2_1 _13604_ (.A(_06770_),
    .B(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__xnor2_1 _13605_ (.A(_06767_),
    .B(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__and3_1 _13606_ (.A(_06721_),
    .B(_06730_),
    .C(_06728_),
    .X(_06777_));
 sky130_fd_sc_hd__a21o_1 _13607_ (.A1(_06762_),
    .A2(_06764_),
    .B1(_06763_),
    .X(_06778_));
 sky130_fd_sc_hd__nand2_1 _13608_ (.A(_06765_),
    .B(_06778_),
    .Y(_06779_));
 sky130_fd_sc_hd__or4_1 _13609_ (.A(_06575_),
    .B(_06702_),
    .C(_06692_),
    .D(_06753_),
    .X(_06780_));
 sky130_fd_sc_hd__and2_1 _13610_ (.A(net555),
    .B(_06759_),
    .X(_06781_));
 sky130_fd_sc_hd__o22ai_1 _13611_ (.A1(_06575_),
    .A2(_06702_),
    .B1(_06692_),
    .B2(_06754_),
    .Y(_06782_));
 sky130_fd_sc_hd__nand3_1 _13612_ (.A(_06780_),
    .B(_06781_),
    .C(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__and2_1 _13613_ (.A(_06780_),
    .B(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__xnor2_1 _13614_ (.A(_06779_),
    .B(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__a21oi_1 _13615_ (.A1(_06730_),
    .A2(_06728_),
    .B1(_06721_),
    .Y(_06786_));
 sky130_fd_sc_hd__o32a_1 _13616_ (.A1(_06777_),
    .A2(_06785_),
    .A3(_06786_),
    .B1(_06779_),
    .B2(_06784_),
    .X(_06787_));
 sky130_fd_sc_hd__xnor2_1 _13617_ (.A(_06776_),
    .B(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__xor2_1 _13618_ (.A(_06747_),
    .B(_06748_),
    .X(_06789_));
 sky130_fd_sc_hd__or2b_1 _13619_ (.A(_06787_),
    .B_N(_06776_),
    .X(_06790_));
 sky130_fd_sc_hd__a21bo_1 _13620_ (.A1(_06788_),
    .A2(_06789_),
    .B1_N(_06790_),
    .X(_06791_));
 sky130_fd_sc_hd__nand2_1 _13621_ (.A(_06759_),
    .B(_06756_),
    .Y(_06792_));
 sky130_fd_sc_hd__inv_2 _13622_ (.A(_06769_),
    .Y(_06793_));
 sky130_fd_sc_hd__nand2_1 _13623_ (.A(_06729_),
    .B(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__a31o_2 _13624_ (.A1(_06436_),
    .A2(_06637_),
    .A3(_06638_),
    .B1(_06642_),
    .X(_06795_));
 sky130_fd_sc_hd__xnor2_4 _13625_ (.A(_06724_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__or2_1 _13626_ (.A(_06693_),
    .B(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__nor2_1 _13627_ (.A(_06576_),
    .B(_06771_),
    .Y(_06798_));
 sky130_fd_sc_hd__xnor2_1 _13628_ (.A(_06797_),
    .B(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__xnor2_1 _13629_ (.A(_06794_),
    .B(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__xnor2_1 _13630_ (.A(_06792_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__or2b_1 _13631_ (.A(_06766_),
    .B_N(_06761_),
    .X(_06802_));
 sky130_fd_sc_hd__and3_1 _13632_ (.A(_06756_),
    .B(_06760_),
    .C(_06766_),
    .X(_06803_));
 sky130_fd_sc_hd__a21o_1 _13633_ (.A1(_06802_),
    .A2(_06775_),
    .B1(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__and2_1 _13634_ (.A(_06801_),
    .B(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__nor2_1 _13635_ (.A(_06801_),
    .B(_06804_),
    .Y(_06806_));
 sky130_fd_sc_hd__nor2_1 _13636_ (.A(_06805_),
    .B(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__buf_6 _13637_ (.A(_06732_),
    .X(_06808_));
 sky130_fd_sc_hd__or3_1 _13638_ (.A(_06715_),
    .B(net544),
    .C(_06739_),
    .X(_06809_));
 sky130_fd_sc_hd__a21bo_1 _13639_ (.A1(_06735_),
    .A2(_06738_),
    .B1_N(_06809_),
    .X(_06810_));
 sky130_fd_sc_hd__and3_1 _13640_ (.A(_06727_),
    .B(_06793_),
    .C(_06774_),
    .X(_06811_));
 sky130_fd_sc_hd__o21bai_1 _13641_ (.A1(_06772_),
    .A2(_06773_),
    .B1_N(_06811_),
    .Y(_06812_));
 sky130_fd_sc_hd__buf_2 _13642_ (.A(net79),
    .X(_06813_));
 sky130_fd_sc_hd__or2_1 _13643_ (.A(_06813_),
    .B(net540),
    .X(_06814_));
 sky130_fd_sc_hd__and2_4 _13644_ (.A(_06683_),
    .B(_06737_),
    .X(_06815_));
 sky130_fd_sc_hd__nor2_2 _13645_ (.A(_06719_),
    .B(net572),
    .Y(_06816_));
 sky130_fd_sc_hd__nor2_1 _13646_ (.A(_06721_),
    .B(_06673_),
    .Y(_06817_));
 sky130_fd_sc_hd__xor2_2 _13647_ (.A(_06816_),
    .B(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__xnor2_2 _13648_ (.A(_06814_),
    .B(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__xnor2_1 _13649_ (.A(_06812_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__xnor2_1 _13650_ (.A(_06810_),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__xnor2_1 _13651_ (.A(_06807_),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__xor2_1 _13652_ (.A(_06791_),
    .B(_06822_),
    .X(_06823_));
 sky130_fd_sc_hd__and2b_1 _13653_ (.A_N(_06751_),
    .B(_06750_),
    .X(_06824_));
 sky130_fd_sc_hd__xnor2_1 _13654_ (.A(_06712_),
    .B(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__or2b_1 _13655_ (.A(_06822_),
    .B_N(_06791_),
    .X(_06826_));
 sky130_fd_sc_hd__o21ai_1 _13656_ (.A1(_06823_),
    .A2(_06825_),
    .B1(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__a21o_1 _13657_ (.A1(_06807_),
    .A2(_06821_),
    .B1(_06805_),
    .X(_06828_));
 sky130_fd_sc_hd__nand2_1 _13658_ (.A(_06577_),
    .B(_06726_),
    .Y(_06829_));
 sky130_fd_sc_hd__o21ai_1 _13659_ (.A1(net83),
    .A2(_06771_),
    .B1(_06829_),
    .Y(_06830_));
 sky130_fd_sc_hd__o21a_1 _13660_ (.A1(_06771_),
    .A2(_06829_),
    .B1(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__buf_4 _13661_ (.A(_06769_),
    .X(_06832_));
 sky130_fd_sc_hd__nor2_1 _13662_ (.A(_06693_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__xnor2_1 _13663_ (.A(_06831_),
    .B(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__a21boi_1 _13664_ (.A1(_06759_),
    .A2(_06800_),
    .B1_N(_06756_),
    .Y(_06835_));
 sky130_fd_sc_hd__nor2_1 _13665_ (.A(_06834_),
    .B(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__and2_1 _13666_ (.A(_06834_),
    .B(_06835_),
    .X(_06837_));
 sky130_fd_sc_hd__nor2_1 _13667_ (.A(_06836_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__inv_2 _13668_ (.A(net541),
    .Y(_06839_));
 sky130_fd_sc_hd__and2_1 _13669_ (.A(_06816_),
    .B(_06817_),
    .X(_06840_));
 sky130_fd_sc_hd__a31oi_2 _13670_ (.A1(_06795_),
    .A2(_06839_),
    .A3(_06818_),
    .B1(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__and2b_1 _13671_ (.A_N(_06797_),
    .B(_06798_),
    .X(_06842_));
 sky130_fd_sc_hd__and3_1 _13672_ (.A(_06729_),
    .B(_06793_),
    .C(_06799_),
    .X(_06843_));
 sky130_fd_sc_hd__o2bb2a_1 _13673_ (.A1_N(_06729_),
    .A2_N(_06721_),
    .B1(net540),
    .B2(_06719_),
    .X(_06844_));
 sky130_fd_sc_hd__a31oi_2 _13674_ (.A1(_06729_),
    .A2(_06721_),
    .A3(_06839_),
    .B1(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__o21a_1 _13675_ (.A1(_06842_),
    .A2(_06843_),
    .B1(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__nor3_1 _13676_ (.A(_06842_),
    .B(_06843_),
    .C(_06845_),
    .Y(_06847_));
 sky130_fd_sc_hd__nor2_1 _13677_ (.A(_06846_),
    .B(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__xnor2_1 _13678_ (.A(_06841_),
    .B(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__xor2_1 _13679_ (.A(_06838_),
    .B(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__xnor2_1 _13680_ (.A(_06828_),
    .B(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__or2b_1 _13681_ (.A(_06713_),
    .B_N(_06717_),
    .X(_06852_));
 sky130_fd_sc_hd__and2b_1 _13682_ (.A_N(_06820_),
    .B(_06810_),
    .X(_06853_));
 sky130_fd_sc_hd__a21o_1 _13683_ (.A1(_06812_),
    .A2(_06819_),
    .B1(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__or3_1 _13684_ (.A(_06715_),
    .B(_06698_),
    .C(_06714_),
    .X(_06855_));
 sky130_fd_sc_hd__or2_1 _13685_ (.A(_06715_),
    .B(_06695_),
    .X(_06856_));
 sky130_fd_sc_hd__or3_1 _13686_ (.A(_06813_),
    .B(_06698_),
    .C(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__o21ai_1 _13687_ (.A1(_06813_),
    .A2(_06698_),
    .B1(_06856_),
    .Y(_06858_));
 sky130_fd_sc_hd__and2_1 _13688_ (.A(_06857_),
    .B(_06858_),
    .X(_06859_));
 sky130_fd_sc_hd__xnor2_1 _13689_ (.A(_06855_),
    .B(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__xnor2_1 _13690_ (.A(_06854_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__xnor2_1 _13691_ (.A(_06852_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__xor2_1 _13692_ (.A(_06851_),
    .B(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__xnor2_1 _13693_ (.A(_06827_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__xnor2_2 _13694_ (.A(_06752_),
    .B(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__xnor2_4 _13695_ (.A(_06744_),
    .B(_06745_),
    .Y(_06866_));
 sky130_fd_sc_hd__or4_4 _13696_ (.A(_06662_),
    .B(_06673_),
    .C(_06771_),
    .D(_06796_),
    .X(_06867_));
 sky130_fd_sc_hd__or2_1 _13697_ (.A(net79),
    .B(_06769_),
    .X(_06868_));
 sky130_fd_sc_hd__a22o_1 _13698_ (.A1(_06727_),
    .A2(_06725_),
    .B1(_06726_),
    .B2(_06768_),
    .X(_06869_));
 sky130_fd_sc_hd__nand3b_1 _13699_ (.A_N(_06868_),
    .B(_06867_),
    .C(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__nand2_1 _13700_ (.A(_06867_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__and2b_1 _13701_ (.A_N(_06866_),
    .B(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__nor2_2 _13702_ (.A(_06705_),
    .B(_06808_),
    .Y(_06873_));
 sky130_fd_sc_hd__or2_1 _13703_ (.A(net80),
    .B(_06734_),
    .X(_06874_));
 sky130_fd_sc_hd__a21oi_1 _13704_ (.A1(_06683_),
    .A2(_06737_),
    .B1(_06634_),
    .Y(_06875_));
 sky130_fd_sc_hd__xnor2_1 _13705_ (.A(_06874_),
    .B(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__or3_4 _13706_ (.A(_06708_),
    .B(_06815_),
    .C(_06874_),
    .X(_06877_));
 sky130_fd_sc_hd__a21bo_1 _13707_ (.A1(_06873_),
    .A2(_06876_),
    .B1_N(_06877_),
    .X(_06878_));
 sky130_fd_sc_hd__xnor2_2 _13708_ (.A(_06871_),
    .B(_06866_),
    .Y(_06879_));
 sky130_fd_sc_hd__and2_1 _13709_ (.A(_06878_),
    .B(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__xor2_1 _13710_ (.A(_06707_),
    .B(_06711_),
    .X(_06881_));
 sky130_fd_sc_hd__o21ai_2 _13711_ (.A1(_06872_),
    .A2(_06880_),
    .B1(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__inv_2 _13712_ (.A(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__or2_1 _13713_ (.A(_06777_),
    .B(_06786_),
    .X(_06884_));
 sky130_fd_sc_hd__xnor2_1 _13714_ (.A(_06785_),
    .B(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__a21o_1 _13715_ (.A1(_06780_),
    .A2(_06782_),
    .B1(_06781_),
    .X(_06886_));
 sky130_fd_sc_hd__nor2_1 _13716_ (.A(_06673_),
    .B(_06755_),
    .Y(_06887_));
 sky130_fd_sc_hd__a2bb2o_1 _13717_ (.A1_N(_06702_),
    .A2_N(_06692_),
    .B1(_06758_),
    .B2(net555),
    .X(_06888_));
 sky130_fd_sc_hd__or4b_1 _13718_ (.A(_06702_),
    .B(_06692_),
    .C(_06705_),
    .D_N(net556),
    .X(_06889_));
 sky130_fd_sc_hd__a21bo_1 _13719_ (.A1(_06887_),
    .A2(_06888_),
    .B1_N(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__and3_1 _13720_ (.A(_06783_),
    .B(_06886_),
    .C(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__a21oi_1 _13721_ (.A1(_06783_),
    .A2(_06886_),
    .B1(_06890_),
    .Y(_06892_));
 sky130_fd_sc_hd__nor2_1 _13722_ (.A(_06891_),
    .B(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__a21bo_1 _13723_ (.A1(_06867_),
    .A2(_06869_),
    .B1_N(_06868_),
    .X(_06894_));
 sky130_fd_sc_hd__and2_1 _13724_ (.A(_06870_),
    .B(_06894_),
    .X(_06895_));
 sky130_fd_sc_hd__a21o_1 _13725_ (.A1(_06893_),
    .A2(_06895_),
    .B1(_06891_),
    .X(_06896_));
 sky130_fd_sc_hd__xnor2_2 _13726_ (.A(_06885_),
    .B(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__xor2_1 _13727_ (.A(net551),
    .B(_06879_),
    .X(_06898_));
 sky130_fd_sc_hd__and2b_1 _13728_ (.A_N(_06885_),
    .B(_06896_),
    .X(_06899_));
 sky130_fd_sc_hd__a21oi_2 _13729_ (.A1(_06897_),
    .A2(net539),
    .B1(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__xnor2_1 _13730_ (.A(_06788_),
    .B(_06789_),
    .Y(_06901_));
 sky130_fd_sc_hd__xnor2_1 _13731_ (.A(_06900_),
    .B(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__or3_1 _13732_ (.A(_06872_),
    .B(_06880_),
    .C(_06881_),
    .X(_06903_));
 sky130_fd_sc_hd__and2_1 _13733_ (.A(_06882_),
    .B(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__or2b_1 _13734_ (.A(net558),
    .B_N(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__o21a_1 _13735_ (.A1(net545),
    .A2(_06901_),
    .B1(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__xor2_1 _13736_ (.A(_06823_),
    .B(_06825_),
    .X(_06907_));
 sky130_fd_sc_hd__xnor2_2 _13737_ (.A(_06906_),
    .B(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__and2b_1 _13738_ (.A_N(_06906_),
    .B(_06907_),
    .X(_06909_));
 sky130_fd_sc_hd__a21oi_2 _13739_ (.A1(_06883_),
    .A2(_06908_),
    .B1(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__xor2_2 _13740_ (.A(_06865_),
    .B(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__xnor2_1 _13741_ (.A(_06873_),
    .B(_06876_),
    .Y(_06912_));
 sky130_fd_sc_hd__xnor2_1 _13742_ (.A(net546),
    .B(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__buf_4 _13743_ (.A(net571),
    .X(_06914_));
 sky130_fd_sc_hd__nor2_1 _13744_ (.A(_06706_),
    .B(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__nor2_1 _13745_ (.A(_06708_),
    .B(net3607),
    .Y(_06916_));
 sky130_fd_sc_hd__nor2_1 _13746_ (.A(_06703_),
    .B(_06808_),
    .Y(_06917_));
 sky130_fd_sc_hd__a21o_1 _13747_ (.A1(_06683_),
    .A2(_06737_),
    .B1(_06705_),
    .X(_06918_));
 sky130_fd_sc_hd__xnor2_1 _13748_ (.A(_06918_),
    .B(_06916_),
    .Y(_06919_));
 sky130_fd_sc_hd__a22o_1 _13749_ (.A1(_06915_),
    .A2(_06916_),
    .B1(_06917_),
    .B2(_06919_),
    .X(_06920_));
 sky130_fd_sc_hd__or2b_1 _13750_ (.A(net3513),
    .B_N(_06920_),
    .X(_06921_));
 sky130_fd_sc_hd__o21ai_1 _13751_ (.A1(net547),
    .A2(_06912_),
    .B1(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__xnor2_1 _13752_ (.A(_06577_),
    .B(net579),
    .Y(_06923_));
 sky130_fd_sc_hd__inv_2 _13753_ (.A(_06706_),
    .Y(_06924_));
 sky130_fd_sc_hd__a2bb2o_1 _13754_ (.A1_N(_06703_),
    .A2_N(_06695_),
    .B1(_06923_),
    .B2(_06924_),
    .X(_06925_));
 sky130_fd_sc_hd__and3_1 _13755_ (.A(_06707_),
    .B(_06922_),
    .C(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__xor2_1 _13756_ (.A(_06893_),
    .B(_06895_),
    .X(_06927_));
 sky130_fd_sc_hd__nand3_1 _13757_ (.A(_06889_),
    .B(_06887_),
    .C(_06888_),
    .Y(_06928_));
 sky130_fd_sc_hd__a21o_1 _13758_ (.A1(_06889_),
    .A2(_06888_),
    .B1(_06887_),
    .X(_06929_));
 sky130_fd_sc_hd__nor2_1 _13759_ (.A(_06719_),
    .B(_06755_),
    .Y(_06930_));
 sky130_fd_sc_hd__inv_2 _13760_ (.A(_06702_),
    .Y(_06931_));
 sky130_fd_sc_hd__a22o_1 _13761_ (.A1(net556),
    .A2(_06931_),
    .B1(_06727_),
    .B2(_06758_),
    .X(_06932_));
 sky130_fd_sc_hd__nand4_2 _13762_ (.A(_06729_),
    .B(_06931_),
    .C(_06727_),
    .D(_06758_),
    .Y(_06933_));
 sky130_fd_sc_hd__a21bo_1 _13763_ (.A1(_06930_),
    .A2(_06932_),
    .B1_N(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__and3_1 _13764_ (.A(_06928_),
    .B(_06929_),
    .C(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__a21oi_1 _13765_ (.A1(_06928_),
    .A2(_06929_),
    .B1(_06934_),
    .Y(_06936_));
 sky130_fd_sc_hd__nor2_1 _13766_ (.A(_06935_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__o2bb2a_1 _13767_ (.A1_N(_06719_),
    .A2_N(_06715_),
    .B1(_06725_),
    .B2(_06793_),
    .X(_06938_));
 sky130_fd_sc_hd__a21oi_1 _13768_ (.A1(_06937_),
    .A2(_06938_),
    .B1(_06935_),
    .Y(_06939_));
 sky130_fd_sc_hd__xnor2_1 _13769_ (.A(_06927_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__xnor2_1 _13770_ (.A(_06920_),
    .B(_06913_),
    .Y(_06941_));
 sky130_fd_sc_hd__and2b_1 _13771_ (.A_N(_06939_),
    .B(_06927_),
    .X(_06942_));
 sky130_fd_sc_hd__a21oi_1 _13772_ (.A1(_06940_),
    .A2(_06941_),
    .B1(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__xor2_1 _13773_ (.A(_06897_),
    .B(_06898_),
    .X(_06944_));
 sky130_fd_sc_hd__xnor2_2 _13774_ (.A(_06943_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__nand2_1 _13775_ (.A(_06707_),
    .B(_06925_),
    .Y(_06946_));
 sky130_fd_sc_hd__xnor2_1 _13776_ (.A(_06922_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__and2b_1 _13777_ (.A_N(_06943_),
    .B(net538),
    .X(_06948_));
 sky130_fd_sc_hd__a21o_1 _13778_ (.A1(net549),
    .A2(_06947_),
    .B1(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__xnor2_2 _13779_ (.A(_06902_),
    .B(_06904_),
    .Y(_06950_));
 sky130_fd_sc_hd__xor2_2 _13780_ (.A(_06949_),
    .B(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__xnor2_2 _13781_ (.A(_06926_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__xnor2_1 _13782_ (.A(_06917_),
    .B(_06919_),
    .Y(_06953_));
 sky130_fd_sc_hd__nor2_1 _13783_ (.A(_06720_),
    .B(net577),
    .Y(_06954_));
 sky130_fd_sc_hd__xor2_1 _13784_ (.A(_06720_),
    .B(_06953_),
    .X(_06955_));
 sky130_fd_sc_hd__nor2_1 _13785_ (.A(_06706_),
    .B(net3634),
    .Y(_06956_));
 sky130_fd_sc_hd__nor2_1 _13786_ (.A(_06703_),
    .B(_06914_),
    .Y(_06957_));
 sky130_fd_sc_hd__and3_1 _13787_ (.A(_06955_),
    .B(_06956_),
    .C(_06957_),
    .X(_06958_));
 sky130_fd_sc_hd__nor2_1 _13788_ (.A(_06703_),
    .B(_06698_),
    .Y(_06959_));
 sky130_fd_sc_hd__o21a_1 _13789_ (.A1(_06954_),
    .A2(_06958_),
    .B1(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__xnor2_1 _13790_ (.A(_06937_),
    .B(_06938_),
    .Y(_06961_));
 sky130_fd_sc_hd__nand3_1 _13791_ (.A(_06933_),
    .B(_06930_),
    .C(_06932_),
    .Y(_06962_));
 sky130_fd_sc_hd__a21o_1 _13792_ (.A1(_06933_),
    .A2(_06932_),
    .B1(_06930_),
    .X(_06963_));
 sky130_fd_sc_hd__nor2_1 _13793_ (.A(net575),
    .B(_06755_),
    .Y(_06964_));
 sky130_fd_sc_hd__a22o_1 _13794_ (.A1(_06931_),
    .A2(_06727_),
    .B1(_06758_),
    .B2(_06768_),
    .X(_06965_));
 sky130_fd_sc_hd__and4_1 _13795_ (.A(_06768_),
    .B(_06931_),
    .C(_06727_),
    .D(_06758_),
    .X(_06966_));
 sky130_fd_sc_hd__a21o_1 _13796_ (.A1(_06964_),
    .A2(_06965_),
    .B1(_06966_),
    .X(_06967_));
 sky130_fd_sc_hd__nand3_1 _13797_ (.A(_06962_),
    .B(_06963_),
    .C(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__a21o_1 _13798_ (.A1(_06962_),
    .A2(_06963_),
    .B1(_06967_),
    .X(_06969_));
 sky130_fd_sc_hd__or2_1 _13799_ (.A(net80),
    .B(net79),
    .X(_06970_));
 sky130_fd_sc_hd__nand2_1 _13800_ (.A(_06715_),
    .B(_06813_),
    .Y(_06971_));
 sky130_fd_sc_hd__nor2_1 _13801_ (.A(_06708_),
    .B(_06832_),
    .Y(_06972_));
 sky130_fd_sc_hd__a41o_1 _13802_ (.A1(net568),
    .A2(_06708_),
    .A3(_06970_),
    .A4(_06971_),
    .B1(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__nand3_1 _13803_ (.A(_06968_),
    .B(_06969_),
    .C(_06973_),
    .Y(_06974_));
 sky130_fd_sc_hd__nand2_1 _13804_ (.A(_06968_),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__xnor2_1 _13805_ (.A(_06961_),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__nand2_1 _13806_ (.A(_06956_),
    .B(_06957_),
    .Y(_06977_));
 sky130_fd_sc_hd__xnor2_1 _13807_ (.A(_06955_),
    .B(_06977_),
    .Y(_06978_));
 sky130_fd_sc_hd__and2b_1 _13808_ (.A_N(_06961_),
    .B(_06975_),
    .X(_06979_));
 sky130_fd_sc_hd__a21oi_1 _13809_ (.A1(_06976_),
    .A2(_06978_),
    .B1(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__xor2_1 _13810_ (.A(_06940_),
    .B(_06941_),
    .X(_06981_));
 sky130_fd_sc_hd__xnor2_2 _13811_ (.A(net578),
    .B(net534),
    .Y(_06982_));
 sky130_fd_sc_hd__nor3_1 _13812_ (.A(_06954_),
    .B(_06958_),
    .C(_06959_),
    .Y(_06983_));
 sky130_fd_sc_hd__nor2_1 _13813_ (.A(_06960_),
    .B(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__or2b_1 _13814_ (.A(_06981_),
    .B_N(_06980_),
    .X(_06985_));
 sky130_fd_sc_hd__a21bo_1 _13815_ (.A1(_06982_),
    .A2(_06984_),
    .B1_N(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__xnor2_2 _13816_ (.A(_06945_),
    .B(_06947_),
    .Y(_06987_));
 sky130_fd_sc_hd__xnor2_2 _13817_ (.A(_06986_),
    .B(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__or2b_1 _13818_ (.A(net537),
    .B_N(_06986_),
    .X(_06989_));
 sky130_fd_sc_hd__a21boi_4 _13819_ (.A1(net3526),
    .A2(net566),
    .B1_N(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__nor2_1 _13820_ (.A(net552),
    .B(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__inv_2 _13821_ (.A(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__xnor2_2 _13822_ (.A(_06882_),
    .B(_06908_),
    .Y(_06993_));
 sky130_fd_sc_hd__nand2_1 _13823_ (.A(_06949_),
    .B(_06950_),
    .Y(_06994_));
 sky130_fd_sc_hd__a21bo_1 _13824_ (.A1(_06926_),
    .A2(net533),
    .B1_N(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__xnor2_2 _13825_ (.A(_06993_),
    .B(_06995_),
    .Y(_06996_));
 sky130_fd_sc_hd__or2_4 _13826_ (.A(_06992_),
    .B(_06996_),
    .X(_06997_));
 sky130_fd_sc_hd__xnor2_1 _13827_ (.A(_06956_),
    .B(_06957_),
    .Y(_06998_));
 sky130_fd_sc_hd__nor2_1 _13828_ (.A(_06706_),
    .B(_06832_),
    .Y(_06999_));
 sky130_fd_sc_hd__nor2_1 _13829_ (.A(net567),
    .B(_06715_),
    .Y(_07000_));
 sky130_fd_sc_hd__mux2_1 _13830_ (.A0(_06813_),
    .A1(_07000_),
    .S(_06708_),
    .X(_07001_));
 sky130_fd_sc_hd__or3_1 _13831_ (.A(_06715_),
    .B(_06708_),
    .C(_06813_),
    .X(_07002_));
 sky130_fd_sc_hd__a21bo_1 _13832_ (.A1(_06999_),
    .A2(_07001_),
    .B1_N(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__nand2b_1 _13833_ (.A_N(_06998_),
    .B(_07003_),
    .Y(_07004_));
 sky130_fd_sc_hd__or2b_1 _13834_ (.A(_07003_),
    .B_N(_06998_),
    .X(_07005_));
 sky130_fd_sc_hd__nand2_1 _13835_ (.A(_07004_),
    .B(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__a21o_1 _13836_ (.A1(_06968_),
    .A2(_06969_),
    .B1(_06973_),
    .X(_07007_));
 sky130_fd_sc_hd__or2b_1 _13837_ (.A(_06966_),
    .B_N(_06965_),
    .X(_07008_));
 sky130_fd_sc_hd__xnor2_2 _13838_ (.A(_06964_),
    .B(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__nor2_1 _13839_ (.A(_06715_),
    .B(_06755_),
    .Y(_07010_));
 sky130_fd_sc_hd__a22o_1 _13840_ (.A1(_06768_),
    .A2(_06931_),
    .B1(_06795_),
    .B2(_06758_),
    .X(_07011_));
 sky130_fd_sc_hd__or4_1 _13841_ (.A(_06719_),
    .B(_06702_),
    .C(_06705_),
    .D(net79),
    .X(_07012_));
 sky130_fd_sc_hd__a21bo_1 _13842_ (.A1(_07010_),
    .A2(_07011_),
    .B1_N(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__xnor2_1 _13843_ (.A(_06999_),
    .B(_07001_),
    .Y(_07014_));
 sky130_fd_sc_hd__xnor2_1 _13844_ (.A(_07009_),
    .B(_07013_),
    .Y(_07015_));
 sky130_fd_sc_hd__nor2_1 _13845_ (.A(_07014_),
    .B(_07015_),
    .Y(_07016_));
 sky130_fd_sc_hd__a21o_1 _13846_ (.A1(_07009_),
    .A2(_07013_),
    .B1(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__a21oi_1 _13847_ (.A1(_06974_),
    .A2(_07007_),
    .B1(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__and3_1 _13848_ (.A(_06974_),
    .B(_07007_),
    .C(_07017_),
    .X(_07019_));
 sky130_fd_sc_hd__o21bai_1 _13849_ (.A1(_07006_),
    .A2(_07018_),
    .B1_N(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__xor2_1 _13850_ (.A(_06976_),
    .B(net548),
    .X(_07021_));
 sky130_fd_sc_hd__nor2_1 _13851_ (.A(_07020_),
    .B(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__and2_1 _13852_ (.A(_07020_),
    .B(_07021_),
    .X(_07023_));
 sky130_fd_sc_hd__o21ba_1 _13853_ (.A1(_07004_),
    .A2(_07022_),
    .B1_N(_07023_),
    .X(_07024_));
 sky130_fd_sc_hd__xor2_2 _13854_ (.A(_06982_),
    .B(_06984_),
    .X(_07025_));
 sky130_fd_sc_hd__xor2_1 _13855_ (.A(_06960_),
    .B(_06988_),
    .X(_07026_));
 sky130_fd_sc_hd__nand3b_2 _13856_ (.A_N(_07024_),
    .B(_07025_),
    .C(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__xor2_2 _13857_ (.A(_06952_),
    .B(_06990_),
    .X(_07028_));
 sky130_fd_sc_hd__or2b_4 _13858_ (.A(_07028_),
    .B_N(_07027_),
    .X(_07029_));
 sky130_fd_sc_hd__xnor2_2 _13859_ (.A(_07027_),
    .B(net529),
    .Y(_07030_));
 sky130_fd_sc_hd__xnor2_1 _13860_ (.A(_07025_),
    .B(_07024_),
    .Y(_07031_));
 sky130_fd_sc_hd__nand2_1 _13861_ (.A(net536),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__clkbuf_4 _13862_ (.A(net3579),
    .X(_07033_));
 sky130_fd_sc_hd__nor2_1 _13863_ (.A(_06703_),
    .B(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__or2_1 _13864_ (.A(net80),
    .B(_06708_),
    .X(_07035_));
 sky130_fd_sc_hd__or3_1 _13865_ (.A(_06706_),
    .B(_07035_),
    .C(_06813_),
    .X(_07036_));
 sky130_fd_sc_hd__o21ai_1 _13866_ (.A1(_06706_),
    .A2(_06796_),
    .B1(_07035_),
    .Y(_07037_));
 sky130_fd_sc_hd__nand2_1 _13867_ (.A(_07036_),
    .B(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__o31ai_2 _13868_ (.A1(_06703_),
    .A2(_06832_),
    .A3(_07038_),
    .B1(_07036_),
    .Y(_07039_));
 sky130_fd_sc_hd__and2_1 _13869_ (.A(_07034_),
    .B(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__and2_1 _13870_ (.A(_07012_),
    .B(_07011_),
    .X(_07041_));
 sky130_fd_sc_hd__xnor2_1 _13871_ (.A(_07010_),
    .B(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__or2_1 _13872_ (.A(_06702_),
    .B(_06813_),
    .X(_07043_));
 sky130_fd_sc_hd__or2_1 _13873_ (.A(_06715_),
    .B(_06754_),
    .X(_07044_));
 sky130_fd_sc_hd__nand2_1 _13874_ (.A(_07043_),
    .B(_07044_),
    .Y(_07045_));
 sky130_fd_sc_hd__nor2_1 _13875_ (.A(net77),
    .B(_06708_),
    .Y(_07046_));
 sky130_fd_sc_hd__nor2_1 _13876_ (.A(_07043_),
    .B(_07044_),
    .Y(_07047_));
 sky130_fd_sc_hd__a21oi_1 _13877_ (.A1(_07045_),
    .A2(_07046_),
    .B1(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__nor2_1 _13878_ (.A(_07042_),
    .B(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__nor2_1 _13879_ (.A(_06703_),
    .B(_06832_),
    .Y(_07050_));
 sky130_fd_sc_hd__xnor2_1 _13880_ (.A(_07038_),
    .B(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__and2_1 _13881_ (.A(_07042_),
    .B(_07048_),
    .X(_07052_));
 sky130_fd_sc_hd__nor2_1 _13882_ (.A(_07049_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__and2_1 _13883_ (.A(_07051_),
    .B(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__and2_1 _13884_ (.A(_07014_),
    .B(_07015_),
    .X(_07055_));
 sky130_fd_sc_hd__nor2_1 _13885_ (.A(_07016_),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__o21a_1 _13886_ (.A1(_07049_),
    .A2(_07054_),
    .B1(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__xnor2_1 _13887_ (.A(_07034_),
    .B(_07039_),
    .Y(_07058_));
 sky130_fd_sc_hd__nor3_1 _13888_ (.A(_07056_),
    .B(_07049_),
    .C(_07054_),
    .Y(_07059_));
 sky130_fd_sc_hd__or2_1 _13889_ (.A(_07057_),
    .B(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__nor2_1 _13890_ (.A(_07058_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__nor2_1 _13891_ (.A(_07019_),
    .B(_07018_),
    .Y(_07062_));
 sky130_fd_sc_hd__xnor2_1 _13892_ (.A(_07006_),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__o21a_1 _13893_ (.A1(_07057_),
    .A2(_07061_),
    .B1(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__nor3_1 _13894_ (.A(_07063_),
    .B(_07057_),
    .C(_07061_),
    .Y(_07065_));
 sky130_fd_sc_hd__nor2_1 _13895_ (.A(_07064_),
    .B(_07065_),
    .Y(_07066_));
 sky130_fd_sc_hd__a21o_1 _13896_ (.A1(_07040_),
    .A2(_07066_),
    .B1(_07064_),
    .X(_07067_));
 sky130_fd_sc_hd__nor2_1 _13897_ (.A(_07023_),
    .B(_07022_),
    .Y(_07068_));
 sky130_fd_sc_hd__xnor2_1 _13898_ (.A(_07004_),
    .B(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__and3b_1 _13899_ (.A_N(_07032_),
    .B(_07067_),
    .C(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__xnor2_2 _13900_ (.A(_07030_),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__clkbuf_4 _13901_ (.A(_06703_),
    .X(_07072_));
 sky130_fd_sc_hd__nor2_1 _13902_ (.A(_07051_),
    .B(_07053_),
    .Y(_07073_));
 sky130_fd_sc_hd__or2_1 _13903_ (.A(_07054_),
    .B(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__o22a_1 _13904_ (.A1(_06706_),
    .A2(_06771_),
    .B1(_06796_),
    .B2(_06703_),
    .X(_07075_));
 sky130_fd_sc_hd__or2_1 _13905_ (.A(_07047_),
    .B(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__or2_1 _13906_ (.A(_07045_),
    .B(_07046_),
    .X(_07077_));
 sky130_fd_sc_hd__a21oi_1 _13907_ (.A1(_07048_),
    .A2(_07077_),
    .B1(_07000_),
    .Y(_07078_));
 sky130_fd_sc_hd__or3_1 _13908_ (.A(_07074_),
    .B(_07076_),
    .C(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__o21ai_1 _13909_ (.A1(_07076_),
    .A2(_07078_),
    .B1(_07074_),
    .Y(_07080_));
 sky130_fd_sc_hd__and2_1 _13910_ (.A(_07079_),
    .B(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__a2bb2o_1 _13911_ (.A1_N(_07047_),
    .A2_N(_07081_),
    .B1(_06706_),
    .B2(_07035_),
    .X(_07082_));
 sky130_fd_sc_hd__nand2_1 _13912_ (.A(_07058_),
    .B(_07060_),
    .Y(_07083_));
 sky130_fd_sc_hd__or2b_1 _13913_ (.A(_07061_),
    .B_N(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__o21a_1 _13914_ (.A1(_07072_),
    .A2(_07082_),
    .B1(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__nand2_1 _13915_ (.A(_07000_),
    .B(_06813_),
    .Y(_07086_));
 sky130_fd_sc_hd__a2bb2o_1 _13916_ (.A1_N(_07040_),
    .A2_N(_07066_),
    .B1(_07086_),
    .B2(_07079_),
    .X(_07087_));
 sky130_fd_sc_hd__nor2_1 _13917_ (.A(_07067_),
    .B(_07069_),
    .Y(_07088_));
 sky130_fd_sc_hd__or4_4 _13918_ (.A(_07032_),
    .B(_07085_),
    .C(_07087_),
    .D(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__nand2_1 _13919_ (.A(_07030_),
    .B(_07070_),
    .Y(_07090_));
 sky130_fd_sc_hd__o21ai_4 _13920_ (.A1(_07071_),
    .A2(_07089_),
    .B1(_07090_),
    .Y(_07091_));
 sky130_fd_sc_hd__and2_4 _13921_ (.A(_06992_),
    .B(_07029_),
    .X(_07092_));
 sky130_fd_sc_hd__xor2_2 _13922_ (.A(_06996_),
    .B(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__a2bb2o_4 _13923_ (.A1_N(net3503),
    .A2_N(_07029_),
    .B1(_07091_),
    .B2(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__nand2_1 _13924_ (.A(_06993_),
    .B(_06995_),
    .Y(_07095_));
 sky130_fd_sc_hd__nand2_2 _13925_ (.A(_07095_),
    .B(_06997_),
    .Y(_07096_));
 sky130_fd_sc_hd__xnor2_2 _13926_ (.A(_06911_),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__a2bb2o_4 _13927_ (.A1_N(_06911_),
    .A2_N(_06997_),
    .B1(_07094_),
    .B2(_07097_),
    .X(_07098_));
 sky130_fd_sc_hd__or2_1 _13928_ (.A(_06852_),
    .B(_06861_),
    .X(_07099_));
 sky130_fd_sc_hd__a21bo_1 _13929_ (.A1(_06854_),
    .A2(_06860_),
    .B1_N(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__nor2_1 _13930_ (.A(_06851_),
    .B(_06862_),
    .Y(_07101_));
 sky130_fd_sc_hd__a21oi_1 _13931_ (.A1(_06828_),
    .A2(_06850_),
    .B1(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__a21o_1 _13932_ (.A1(_06838_),
    .A2(_06849_),
    .B1(_06836_),
    .X(_07103_));
 sky130_fd_sc_hd__clkbuf_2 _13933_ (.A(net83),
    .X(_07104_));
 sky130_fd_sc_hd__nor2_1 _13934_ (.A(_07104_),
    .B(_06796_),
    .Y(_07105_));
 sky130_fd_sc_hd__nor2_1 _13935_ (.A(_06576_),
    .B(_06832_),
    .Y(_07106_));
 sky130_fd_sc_hd__xor2_1 _13936_ (.A(_07105_),
    .B(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__a2bb2o_1 _13937_ (.A1_N(_06771_),
    .A2_N(_06829_),
    .B1(_06830_),
    .B2(_06833_),
    .X(_07108_));
 sky130_fd_sc_hd__inv_2 _13938_ (.A(net3533),
    .Y(_07109_));
 sky130_fd_sc_hd__o22a_1 _13939_ (.A1(_06727_),
    .A2(net541),
    .B1(_07109_),
    .B2(_06693_),
    .X(_07110_));
 sky130_fd_sc_hd__xor2_1 _13940_ (.A(_07108_),
    .B(_07110_),
    .X(_07111_));
 sky130_fd_sc_hd__a21oi_1 _13941_ (.A1(_06721_),
    .A2(_06693_),
    .B1(_06683_),
    .Y(_07112_));
 sky130_fd_sc_hd__xor2_1 _13942_ (.A(_07111_),
    .B(_07112_),
    .X(_07113_));
 sky130_fd_sc_hd__nand2_1 _13943_ (.A(_07107_),
    .B(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__or2_1 _13944_ (.A(_07107_),
    .B(_07113_),
    .X(_07115_));
 sky130_fd_sc_hd__nand2_1 _13945_ (.A(_07114_),
    .B(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__xor2_1 _13946_ (.A(_07103_),
    .B(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__or2b_1 _13947_ (.A(_06855_),
    .B_N(_06859_),
    .X(_07118_));
 sky130_fd_sc_hd__and2b_1 _13948_ (.A_N(_06841_),
    .B(_06848_),
    .X(_07119_));
 sky130_fd_sc_hd__or2_1 _13949_ (.A(_06846_),
    .B(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__or2_1 _13950_ (.A(_06813_),
    .B(_06695_),
    .X(_07121_));
 sky130_fd_sc_hd__or3_1 _13951_ (.A(_06719_),
    .B(_06698_),
    .C(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__o21ai_1 _13952_ (.A1(_06719_),
    .A2(_06698_),
    .B1(_07121_),
    .Y(_07123_));
 sky130_fd_sc_hd__and2_1 _13953_ (.A(_07122_),
    .B(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__xnor2_1 _13954_ (.A(_06857_),
    .B(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__xnor2_2 _13955_ (.A(_07120_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__xnor2_1 _13956_ (.A(_07118_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__or2_1 _13957_ (.A(_07117_),
    .B(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__nand2_1 _13958_ (.A(_07117_),
    .B(_07127_),
    .Y(_07129_));
 sky130_fd_sc_hd__and2_1 _13959_ (.A(_07128_),
    .B(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__xnor2_2 _13960_ (.A(_07102_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__xnor2_1 _13961_ (.A(_07100_),
    .B(_07131_),
    .Y(_07132_));
 sky130_fd_sc_hd__or2b_1 _13962_ (.A(_06864_),
    .B_N(_06752_),
    .X(_07133_));
 sky130_fd_sc_hd__a21boi_1 _13963_ (.A1(_06827_),
    .A2(_06863_),
    .B1_N(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__nor2_2 _13964_ (.A(_07134_),
    .B(_07132_),
    .Y(_07135_));
 sky130_fd_sc_hd__nand2_1 _13965_ (.A(_07132_),
    .B(_07134_),
    .Y(_07136_));
 sky130_fd_sc_hd__and2b_1 _13966_ (.A_N(_07135_),
    .B(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__and2b_1 _13967_ (.A_N(_06910_),
    .B(_06865_),
    .X(_07138_));
 sky130_fd_sc_hd__nor2_1 _13968_ (.A(_06911_),
    .B(_07095_),
    .Y(_07139_));
 sky130_fd_sc_hd__nor2_1 _13969_ (.A(_07138_),
    .B(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__xnor2_1 _13970_ (.A(_07137_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__xnor2_1 _13971_ (.A(_07098_),
    .B(_07141_),
    .Y(_07142_));
 sky130_fd_sc_hd__xor2_1 _13972_ (.A(_07094_),
    .B(_07097_),
    .X(_07143_));
 sky130_fd_sc_hd__xnor2_2 _13973_ (.A(net3498),
    .B(_07093_),
    .Y(_07144_));
 sky130_fd_sc_hd__xnor2_4 _13974_ (.A(net535),
    .B(_07089_),
    .Y(_07145_));
 sky130_fd_sc_hd__nor2_2 _13975_ (.A(_07144_),
    .B(_07145_),
    .Y(_07146_));
 sky130_fd_sc_hd__nor2_2 _13976_ (.A(_07143_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__nand2_2 _13977_ (.A(_07142_),
    .B(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__or2b_1 _13978_ (.A(_07102_),
    .B_N(_07130_),
    .X(_07149_));
 sky130_fd_sc_hd__nand2_1 _13979_ (.A(_07100_),
    .B(_07131_),
    .Y(_07150_));
 sky130_fd_sc_hd__or2b_1 _13980_ (.A(_07116_),
    .B_N(_07103_),
    .X(_07151_));
 sky130_fd_sc_hd__nand2_1 _13981_ (.A(_07105_),
    .B(_07106_),
    .Y(_07152_));
 sky130_fd_sc_hd__nand2_1 _13982_ (.A(_06729_),
    .B(_06839_),
    .Y(_07153_));
 sky130_fd_sc_hd__and4bb_1 _13983_ (.A_N(_06693_),
    .B_N(net573),
    .C(_07109_),
    .D(_06577_),
    .X(_07154_));
 sky130_fd_sc_hd__o22a_1 _13984_ (.A1(_06576_),
    .A2(net3533),
    .B1(net571),
    .B2(_06693_),
    .X(_07155_));
 sky130_fd_sc_hd__nor2_1 _13985_ (.A(_07154_),
    .B(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__xnor2_2 _13986_ (.A(_07153_),
    .B(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__xnor2_2 _13987_ (.A(_07152_),
    .B(_07157_),
    .Y(_07158_));
 sky130_fd_sc_hd__xnor2_1 _13988_ (.A(net581),
    .B(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__and3b_1 _13989_ (.A_N(_07159_),
    .B(_06793_),
    .C(_06757_),
    .X(_07160_));
 sky130_fd_sc_hd__o21a_1 _13990_ (.A1(_07104_),
    .A2(_06832_),
    .B1(_07159_),
    .X(_07161_));
 sky130_fd_sc_hd__or2_1 _13991_ (.A(_07160_),
    .B(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__xnor2_1 _13992_ (.A(_07114_),
    .B(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__and2b_1 _13993_ (.A_N(_06857_),
    .B(_07124_),
    .X(_07164_));
 sky130_fd_sc_hd__and2_1 _13994_ (.A(_07108_),
    .B(_07110_),
    .X(_07165_));
 sky130_fd_sc_hd__and2_1 _13995_ (.A(_07111_),
    .B(_07112_),
    .X(_07166_));
 sky130_fd_sc_hd__or2_1 _13996_ (.A(_06719_),
    .B(_06695_),
    .X(_07167_));
 sky130_fd_sc_hd__or3_1 _13997_ (.A(_06673_),
    .B(_06698_),
    .C(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__o21ai_1 _13998_ (.A1(_06673_),
    .A2(_06698_),
    .B1(_07167_),
    .Y(_07169_));
 sky130_fd_sc_hd__and2_1 _13999_ (.A(_07168_),
    .B(_07169_),
    .X(_07170_));
 sky130_fd_sc_hd__xnor2_1 _14000_ (.A(_07122_),
    .B(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__o21a_1 _14001_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__nor3_1 _14002_ (.A(_07165_),
    .B(_07166_),
    .C(_07171_),
    .Y(_07173_));
 sky130_fd_sc_hd__nor2_1 _14003_ (.A(_07172_),
    .B(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__xnor2_1 _14004_ (.A(_07164_),
    .B(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__xnor2_1 _14005_ (.A(_07163_),
    .B(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__a21o_1 _14006_ (.A1(_07151_),
    .A2(_07128_),
    .B1(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__nand3_1 _14007_ (.A(_07151_),
    .B(_07128_),
    .C(_07176_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_1 _14008_ (.A(_07177_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__nand2_1 _14009_ (.A(_07120_),
    .B(_07125_),
    .Y(_07180_));
 sky130_fd_sc_hd__o21a_1 _14010_ (.A1(_07118_),
    .A2(_07126_),
    .B1(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__xnor2_1 _14011_ (.A(_07179_),
    .B(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__a21oi_2 _14012_ (.A1(_07149_),
    .A2(_07150_),
    .B1(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__and3_1 _14013_ (.A(_07149_),
    .B(_07150_),
    .C(_07182_),
    .X(_07184_));
 sky130_fd_sc_hd__or2_1 _14014_ (.A(_07183_),
    .B(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__inv_2 _14015_ (.A(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__a21oi_1 _14016_ (.A1(_07138_),
    .A2(_07136_),
    .B1(_07135_),
    .Y(_07187_));
 sky130_fd_sc_hd__xnor2_1 _14017_ (.A(_07186_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__a22o_1 _14018_ (.A1(_07137_),
    .A2(_07139_),
    .B1(_07141_),
    .B2(_07098_),
    .X(_07189_));
 sky130_fd_sc_hd__xor2_1 _14019_ (.A(_07188_),
    .B(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__or2_4 _14020_ (.A(_07148_),
    .B(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__nand2_1 _14021_ (.A(_07148_),
    .B(_07190_),
    .Y(_07192_));
 sky130_fd_sc_hd__nand2_2 _14022_ (.A(_07191_),
    .B(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__clkbuf_4 _14023_ (.A(_07193_),
    .X(_07194_));
 sky130_fd_sc_hd__or2_1 _14024_ (.A(_06699_),
    .B(_07194_),
    .X(_07195_));
 sky130_fd_sc_hd__or2_1 _14025_ (.A(_07142_),
    .B(_07147_),
    .X(_07196_));
 sky130_fd_sc_hd__nand2_2 _14026_ (.A(_07148_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__clkbuf_4 _14027_ (.A(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__or3_1 _14028_ (.A(_06696_),
    .B(_07195_),
    .C(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__a32o_2 _14029_ (.A1(_07138_),
    .A2(_07137_),
    .A3(_07186_),
    .B1(_07188_),
    .B2(_07189_),
    .X(_07200_));
 sky130_fd_sc_hd__or2_1 _14030_ (.A(_07179_),
    .B(_07181_),
    .X(_07201_));
 sky130_fd_sc_hd__or2_1 _14031_ (.A(_07163_),
    .B(_07175_),
    .X(_07202_));
 sky130_fd_sc_hd__o21ai_1 _14032_ (.A1(_07114_),
    .A2(_07162_),
    .B1(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__or3_1 _14033_ (.A(_06576_),
    .B(net3579),
    .C(_06914_),
    .X(_07204_));
 sky130_fd_sc_hd__o21ai_1 _14034_ (.A1(_06576_),
    .A2(_06914_),
    .B1(net3579),
    .Y(_07205_));
 sky130_fd_sc_hd__and2_1 _14035_ (.A(_07204_),
    .B(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__nand2_1 _14036_ (.A(_07160_),
    .B(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__or2_1 _14037_ (.A(_07160_),
    .B(_07206_),
    .X(_07208_));
 sky130_fd_sc_hd__nand2_1 _14038_ (.A(_07207_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__or2b_1 _14039_ (.A(_07122_),
    .B_N(_07170_),
    .X(_07210_));
 sky130_fd_sc_hd__a32o_1 _14040_ (.A1(_07105_),
    .A2(_07106_),
    .A3(_07157_),
    .B1(_07158_),
    .B2(_06694_),
    .X(_07211_));
 sky130_fd_sc_hd__or2_1 _14041_ (.A(_06673_),
    .B(_06695_),
    .X(_07212_));
 sky130_fd_sc_hd__nand2_1 _14042_ (.A(_06729_),
    .B(_06923_),
    .Y(_07213_));
 sky130_fd_sc_hd__xor2_1 _14043_ (.A(_07212_),
    .B(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__xnor2_1 _14044_ (.A(_07168_),
    .B(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__nand2_1 _14045_ (.A(_07211_),
    .B(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__or2_1 _14046_ (.A(_07211_),
    .B(_07215_),
    .X(_07217_));
 sky130_fd_sc_hd__nand2_1 _14047_ (.A(_07216_),
    .B(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__xor2_1 _14048_ (.A(_07210_),
    .B(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__xnor2_1 _14049_ (.A(_07209_),
    .B(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__xnor2_1 _14050_ (.A(_07203_),
    .B(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__a21oi_1 _14051_ (.A1(_07164_),
    .A2(_07174_),
    .B1(_07172_),
    .Y(_07222_));
 sky130_fd_sc_hd__xnor2_1 _14052_ (.A(_07221_),
    .B(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__a21oi_1 _14053_ (.A1(_07177_),
    .A2(_07201_),
    .B1(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__and3_1 _14054_ (.A(_07177_),
    .B(_07201_),
    .C(_07223_),
    .X(_07225_));
 sky130_fd_sc_hd__nor2_2 _14055_ (.A(_07224_),
    .B(_07225_),
    .Y(_07226_));
 sky130_fd_sc_hd__xor2_1 _14056_ (.A(_07183_),
    .B(_07226_),
    .X(_07227_));
 sky130_fd_sc_hd__nand3_1 _14057_ (.A(_07135_),
    .B(_07186_),
    .C(_07227_),
    .Y(_07228_));
 sky130_fd_sc_hd__a21o_1 _14058_ (.A1(_07135_),
    .A2(_07186_),
    .B1(_07227_),
    .X(_07229_));
 sky130_fd_sc_hd__and2_4 _14059_ (.A(_07228_),
    .B(_07229_),
    .X(_07230_));
 sky130_fd_sc_hd__xor2_2 _14060_ (.A(_07200_),
    .B(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__xnor2_1 _14061_ (.A(_07191_),
    .B(_07231_),
    .Y(_07232_));
 sky130_fd_sc_hd__buf_4 _14062_ (.A(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__nor2_1 _14063_ (.A(_06699_),
    .B(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__nor2_1 _14064_ (.A(_06696_),
    .B(_07194_),
    .Y(_07235_));
 sky130_fd_sc_hd__xnor2_1 _14065_ (.A(_07234_),
    .B(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__or2_1 _14066_ (.A(_07199_),
    .B(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__nand2_1 _14067_ (.A(_07199_),
    .B(_07236_),
    .Y(_07238_));
 sky130_fd_sc_hd__nand2_1 _14068_ (.A(_07237_),
    .B(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__clkbuf_4 _14069_ (.A(net543),
    .X(_07240_));
 sky130_fd_sc_hd__or2_1 _14070_ (.A(_07240_),
    .B(_07194_),
    .X(_07241_));
 sky130_fd_sc_hd__clkbuf_4 _14071_ (.A(_06914_),
    .X(_07242_));
 sky130_fd_sc_hd__nor2_4 _14072_ (.A(_07191_),
    .B(_07231_),
    .Y(_07243_));
 sky130_fd_sc_hd__a21boi_4 _14073_ (.A1(_07200_),
    .A2(_07230_),
    .B1_N(_07228_),
    .Y(_07244_));
 sky130_fd_sc_hd__nand2_2 _14074_ (.A(_07183_),
    .B(_07226_),
    .Y(_07245_));
 sky130_fd_sc_hd__nand2_1 _14075_ (.A(_07203_),
    .B(_07220_),
    .Y(_07246_));
 sky130_fd_sc_hd__or2_1 _14076_ (.A(_07221_),
    .B(_07222_),
    .X(_07247_));
 sky130_fd_sc_hd__or2b_1 _14077_ (.A(_07209_),
    .B_N(_07219_),
    .X(_07248_));
 sky130_fd_sc_hd__nand2_1 _14078_ (.A(net580),
    .B(_07206_),
    .Y(_07249_));
 sky130_fd_sc_hd__or4_1 _14079_ (.A(_07104_),
    .B(_06576_),
    .C(net541),
    .D(_06914_),
    .X(_07250_));
 sky130_fd_sc_hd__inv_2 _14080_ (.A(_06914_),
    .Y(_07251_));
 sky130_fd_sc_hd__a22o_1 _14081_ (.A1(_06577_),
    .A2(_06839_),
    .B1(_07251_),
    .B2(net5902),
    .X(_07252_));
 sky130_fd_sc_hd__nand2_1 _14082_ (.A(_07250_),
    .B(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__a21oi_1 _14083_ (.A1(_07204_),
    .A2(_07249_),
    .B1(_07253_),
    .Y(_07254_));
 sky130_fd_sc_hd__and3_1 _14084_ (.A(_07204_),
    .B(_07249_),
    .C(_07253_),
    .X(_07255_));
 sky130_fd_sc_hd__or2_1 _14085_ (.A(_07254_),
    .B(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__or2b_1 _14086_ (.A(_07168_),
    .B_N(_07214_),
    .X(_07257_));
 sky130_fd_sc_hd__or2_1 _14087_ (.A(_07212_),
    .B(_07213_),
    .X(_07258_));
 sky130_fd_sc_hd__and2b_1 _14088_ (.A_N(_06695_),
    .B(_06729_),
    .X(_07259_));
 sky130_fd_sc_hd__or2_1 _14089_ (.A(_06693_),
    .B(_06698_),
    .X(_07260_));
 sky130_fd_sc_hd__xnor2_1 _14090_ (.A(_07259_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__nand2_1 _14091_ (.A(net580),
    .B(_07249_),
    .Y(_07262_));
 sky130_fd_sc_hd__and3_1 _14092_ (.A(_07258_),
    .B(_07261_),
    .C(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__xnor2_1 _14093_ (.A(_07257_),
    .B(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__xor2_1 _14094_ (.A(_07256_),
    .B(_07264_),
    .X(_07265_));
 sky130_fd_sc_hd__a21oi_1 _14095_ (.A1(_07207_),
    .A2(_07248_),
    .B1(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__and3_1 _14096_ (.A(_07207_),
    .B(_07248_),
    .C(_07265_),
    .X(_07267_));
 sky130_fd_sc_hd__nor2_1 _14097_ (.A(_07266_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__o21a_1 _14098_ (.A1(_07210_),
    .A2(_07218_),
    .B1(_07216_),
    .X(_07269_));
 sky130_fd_sc_hd__inv_2 _14099_ (.A(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__xnor2_1 _14100_ (.A(_07268_),
    .B(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__a21o_1 _14101_ (.A1(_07246_),
    .A2(_07247_),
    .B1(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__nand3_1 _14102_ (.A(_07246_),
    .B(_07247_),
    .C(_07271_),
    .Y(_07273_));
 sky130_fd_sc_hd__and2_1 _14103_ (.A(_07272_),
    .B(_07273_),
    .X(_07274_));
 sky130_fd_sc_hd__nand2_1 _14104_ (.A(_07224_),
    .B(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__or2_1 _14105_ (.A(_07224_),
    .B(_07274_),
    .X(_07276_));
 sky130_fd_sc_hd__nand2_2 _14106_ (.A(_07275_),
    .B(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__xnor2_4 _14107_ (.A(_07245_),
    .B(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__xnor2_4 _14108_ (.A(_07244_),
    .B(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__xnor2_4 _14109_ (.A(_07243_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__clkbuf_4 _14110_ (.A(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__o22a_1 _14111_ (.A1(_07242_),
    .A2(_07233_),
    .B1(_07281_),
    .B2(_07033_),
    .X(_07282_));
 sky130_fd_sc_hd__nor2_2 _14112_ (.A(_07241_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__clkbuf_4 _14113_ (.A(_06832_),
    .X(_07284_));
 sky130_fd_sc_hd__a21oi_1 _14114_ (.A1(_07268_),
    .A2(_07270_),
    .B1(_07266_),
    .Y(_07285_));
 sky130_fd_sc_hd__or2b_1 _14115_ (.A(_07256_),
    .B_N(_07264_),
    .X(_07286_));
 sky130_fd_sc_hd__a211o_1 _14116_ (.A1(_06577_),
    .A2(_07251_),
    .B1(net542),
    .C1(_07104_),
    .X(_07287_));
 sky130_fd_sc_hd__inv_2 _14117_ (.A(_07254_),
    .Y(_07288_));
 sky130_fd_sc_hd__a21o_1 _14118_ (.A1(_06923_),
    .A2(_07259_),
    .B1(_06693_),
    .X(_07289_));
 sky130_fd_sc_hd__nor2_1 _14119_ (.A(_07288_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__and2_1 _14120_ (.A(_07288_),
    .B(_07289_),
    .X(_07291_));
 sky130_fd_sc_hd__o21ai_1 _14121_ (.A1(_07290_),
    .A2(_07291_),
    .B1(_07258_),
    .Y(_07292_));
 sky130_fd_sc_hd__xnor2_1 _14122_ (.A(_07287_),
    .B(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__xnor2_1 _14123_ (.A(_07286_),
    .B(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__inv_2 _14124_ (.A(_07263_),
    .Y(_07295_));
 sky130_fd_sc_hd__o21a_1 _14125_ (.A1(_07257_),
    .A2(_07295_),
    .B1(_07262_),
    .X(_07296_));
 sky130_fd_sc_hd__xnor2_1 _14126_ (.A(_07294_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__xnor2_1 _14127_ (.A(_07285_),
    .B(_07297_),
    .Y(_07298_));
 sky130_fd_sc_hd__xnor2_1 _14128_ (.A(_07272_),
    .B(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__nand2_1 _14129_ (.A(_07200_),
    .B(_07230_),
    .Y(_07300_));
 sky130_fd_sc_hd__a21o_1 _14130_ (.A1(_07245_),
    .A2(_07228_),
    .B1(_07277_),
    .X(_07301_));
 sky130_fd_sc_hd__o211a_1 _14131_ (.A1(_07300_),
    .A2(_07278_),
    .B1(_07301_),
    .C1(_07275_),
    .X(_07302_));
 sky130_fd_sc_hd__a22o_4 _14132_ (.A1(_07243_),
    .A2(_07279_),
    .B1(_07299_),
    .B2(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__buf_6 _14133_ (.A(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__buf_2 _14134_ (.A(_07304_),
    .X(_07305_));
 sky130_fd_sc_hd__clkbuf_4 _14135_ (.A(_06771_),
    .X(_07306_));
 sky130_fd_sc_hd__nor2_2 _14136_ (.A(_07306_),
    .B(_07303_),
    .Y(_07307_));
 sky130_fd_sc_hd__clkbuf_4 _14137_ (.A(_06796_),
    .X(_07308_));
 sky130_fd_sc_hd__nor2_2 _14138_ (.A(_07308_),
    .B(_07303_),
    .Y(_07309_));
 sky130_fd_sc_hd__xnor2_4 _14139_ (.A(_07307_),
    .B(_07309_),
    .Y(_07310_));
 sky130_fd_sc_hd__nand2_1 _14140_ (.A(_07307_),
    .B(_07309_),
    .Y(_07311_));
 sky130_fd_sc_hd__o31a_1 _14141_ (.A1(_07284_),
    .A2(_07305_),
    .A3(_07310_),
    .B1(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__nor2_1 _14142_ (.A(_07240_),
    .B(_07233_),
    .Y(_07313_));
 sky130_fd_sc_hd__nor2_2 _14143_ (.A(_07033_),
    .B(net569),
    .Y(_07314_));
 sky130_fd_sc_hd__nor2_1 _14144_ (.A(_07242_),
    .B(_07281_),
    .Y(_07315_));
 sky130_fd_sc_hd__xor2_1 _14145_ (.A(_07314_),
    .B(_07315_),
    .X(_07316_));
 sky130_fd_sc_hd__and2_1 _14146_ (.A(_07313_),
    .B(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__nor2_1 _14147_ (.A(_07313_),
    .B(_07316_),
    .Y(_07318_));
 sky130_fd_sc_hd__or2_1 _14148_ (.A(_07317_),
    .B(_07318_),
    .X(_07319_));
 sky130_fd_sc_hd__xor2_2 _14149_ (.A(_07312_),
    .B(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__nor2_1 _14150_ (.A(_07312_),
    .B(_07319_),
    .Y(_07321_));
 sky130_fd_sc_hd__a21oi_2 _14151_ (.A1(_07283_),
    .A2(_07320_),
    .B1(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__or2_1 _14152_ (.A(_06699_),
    .B(_07198_),
    .X(_07323_));
 sky130_fd_sc_hd__and2_1 _14153_ (.A(_07143_),
    .B(_07146_),
    .X(_07324_));
 sky130_fd_sc_hd__or2_1 _14154_ (.A(_07147_),
    .B(_07324_),
    .X(_07325_));
 sky130_fd_sc_hd__clkbuf_2 _14155_ (.A(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__clkbuf_4 _14156_ (.A(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__or3_1 _14157_ (.A(_06696_),
    .B(_07323_),
    .C(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__nor2_1 _14158_ (.A(_06696_),
    .B(_07198_),
    .Y(_07329_));
 sky130_fd_sc_hd__xnor2_1 _14159_ (.A(_07195_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__and2b_1 _14160_ (.A_N(_07328_),
    .B(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__xor2_1 _14161_ (.A(_07239_),
    .B(_07322_),
    .X(_07332_));
 sky130_fd_sc_hd__nand2_1 _14162_ (.A(_07331_),
    .B(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__o21ai_2 _14163_ (.A1(_07239_),
    .A2(_07322_),
    .B1(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__nand2_1 _14164_ (.A(_07234_),
    .B(_07235_),
    .Y(_07335_));
 sky130_fd_sc_hd__nor2_1 _14165_ (.A(_06699_),
    .B(_07281_),
    .Y(_07336_));
 sky130_fd_sc_hd__nor2_1 _14166_ (.A(_06696_),
    .B(_07233_),
    .Y(_07337_));
 sky130_fd_sc_hd__xnor2_1 _14167_ (.A(_07336_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__or2_1 _14168_ (.A(_07335_),
    .B(_07338_),
    .X(_07339_));
 sky130_fd_sc_hd__nand2_1 _14169_ (.A(_07335_),
    .B(_07338_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2_1 _14170_ (.A(_07339_),
    .B(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__and2_4 _14171_ (.A(net5902),
    .B(_07304_),
    .X(_07342_));
 sky130_fd_sc_hd__a21oi_1 _14172_ (.A1(_06725_),
    .A2(_07342_),
    .B1(_07309_),
    .Y(_07343_));
 sky130_fd_sc_hd__nor2_1 _14173_ (.A(_07284_),
    .B(_07305_),
    .Y(_07344_));
 sky130_fd_sc_hd__nor2b_1 _14174_ (.A(_07343_),
    .B_N(_07344_),
    .Y(_07345_));
 sky130_fd_sc_hd__nor2_1 _14175_ (.A(_07242_),
    .B(net569),
    .Y(_07346_));
 sky130_fd_sc_hd__xor2_2 _14176_ (.A(_07314_),
    .B(_07346_),
    .X(_07347_));
 sky130_fd_sc_hd__nor2_1 _14177_ (.A(_07240_),
    .B(_07281_),
    .Y(_07348_));
 sky130_fd_sc_hd__xor2_1 _14178_ (.A(_07347_),
    .B(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__xnor2_1 _14179_ (.A(_07345_),
    .B(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__a21oi_1 _14180_ (.A1(_07314_),
    .A2(_07315_),
    .B1(_07317_),
    .Y(_07351_));
 sky130_fd_sc_hd__nor2_1 _14181_ (.A(_07350_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__a21oi_1 _14182_ (.A1(_07345_),
    .A2(_07349_),
    .B1(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__xor2_1 _14183_ (.A(_07341_),
    .B(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__xnor2_1 _14184_ (.A(_07237_),
    .B(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__and2_1 _14185_ (.A(_07350_),
    .B(_07351_),
    .X(_07356_));
 sky130_fd_sc_hd__or2_1 _14186_ (.A(_07352_),
    .B(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__a211o_1 _14187_ (.A1(_06726_),
    .A2(_07342_),
    .B1(_07344_),
    .C1(net8355),
    .X(_07358_));
 sky130_fd_sc_hd__or2b_1 _14188_ (.A(_07357_),
    .B_N(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__inv_2 _14189_ (.A(_07342_),
    .Y(_07360_));
 sky130_fd_sc_hd__nand2_1 _14190_ (.A(_07314_),
    .B(_07346_),
    .Y(_07361_));
 sky130_fd_sc_hd__nand2_1 _14191_ (.A(_07347_),
    .B(_07348_),
    .Y(_07362_));
 sky130_fd_sc_hd__nor2_1 _14192_ (.A(_07240_),
    .B(_07305_),
    .Y(_07363_));
 sky130_fd_sc_hd__xnor2_1 _14193_ (.A(_07347_),
    .B(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__a31o_1 _14194_ (.A1(_07361_),
    .A2(_07362_),
    .A3(_07364_),
    .B1(_07290_),
    .X(_07365_));
 sky130_fd_sc_hd__o211a_1 _14195_ (.A1(_07284_),
    .A2(_07360_),
    .B1(_07365_),
    .C1(net5902),
    .X(_07366_));
 sky130_fd_sc_hd__xor2_1 _14196_ (.A(_07359_),
    .B(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__nand2_1 _14197_ (.A(_07355_),
    .B(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__or2_1 _14198_ (.A(_07355_),
    .B(_07367_),
    .X(_07369_));
 sky130_fd_sc_hd__nand2_1 _14199_ (.A(_07368_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__or2_1 _14200_ (.A(_07331_),
    .B(_07332_),
    .X(_07371_));
 sky130_fd_sc_hd__nand2_1 _14201_ (.A(_07333_),
    .B(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__and2b_1 _14202_ (.A_N(_07344_),
    .B(_07343_),
    .X(_07373_));
 sky130_fd_sc_hd__nor2_1 _14203_ (.A(_07345_),
    .B(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__xor2_2 _14204_ (.A(_07283_),
    .B(_07320_),
    .X(_07375_));
 sky130_fd_sc_hd__xnor2_1 _14205_ (.A(_07358_),
    .B(_07357_),
    .Y(_07376_));
 sky130_fd_sc_hd__a21oi_1 _14206_ (.A1(_07374_),
    .A2(_07375_),
    .B1(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__and3_1 _14207_ (.A(_07374_),
    .B(_07375_),
    .C(_07376_),
    .X(_07378_));
 sky130_fd_sc_hd__o21ba_1 _14208_ (.A1(_07372_),
    .A2(_07377_),
    .B1_N(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__nor2_1 _14209_ (.A(_07370_),
    .B(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__and2_1 _14210_ (.A(_07370_),
    .B(_07379_),
    .X(_07381_));
 sky130_fd_sc_hd__nor2_1 _14211_ (.A(_07380_),
    .B(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__xnor2_1 _14212_ (.A(_07334_),
    .B(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__or2_1 _14213_ (.A(_07378_),
    .B(_07377_),
    .X(_07384_));
 sky130_fd_sc_hd__xnor2_1 _14214_ (.A(_07372_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__o21ai_1 _14215_ (.A1(_06696_),
    .A2(_07327_),
    .B1(_07323_),
    .Y(_07386_));
 sky130_fd_sc_hd__and2_1 _14216_ (.A(_07328_),
    .B(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__or2_1 _14217_ (.A(_06699_),
    .B(_07327_),
    .X(_07388_));
 sky130_fd_sc_hd__and2_1 _14218_ (.A(_07144_),
    .B(_07145_),
    .X(_07389_));
 sky130_fd_sc_hd__nor2_2 _14219_ (.A(_07146_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__clkbuf_4 _14220_ (.A(_07390_),
    .X(_07391_));
 sky130_fd_sc_hd__nor2_1 _14221_ (.A(_06696_),
    .B(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__and2b_1 _14222_ (.A_N(_07388_),
    .B(_07392_),
    .X(_07393_));
 sky130_fd_sc_hd__o21ai_2 _14223_ (.A1(net8355),
    .A2(_07387_),
    .B1(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__xor2_1 _14224_ (.A(_07328_),
    .B(_07330_),
    .X(_07395_));
 sky130_fd_sc_hd__or3_1 _14225_ (.A(_07284_),
    .B(_07310_),
    .C(_07281_),
    .X(_07396_));
 sky130_fd_sc_hd__and2_1 _14226_ (.A(_07241_),
    .B(_07282_),
    .X(_07397_));
 sky130_fd_sc_hd__or2_1 _14227_ (.A(_07283_),
    .B(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__a21o_1 _14228_ (.A1(_07311_),
    .A2(_07396_),
    .B1(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__nand3_1 _14229_ (.A(_07311_),
    .B(_07396_),
    .C(_07398_),
    .Y(_07400_));
 sky130_fd_sc_hd__nand2_2 _14230_ (.A(_07399_),
    .B(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__nor2_1 _14231_ (.A(_07240_),
    .B(_07198_),
    .Y(_07402_));
 sky130_fd_sc_hd__or2_1 _14232_ (.A(_07033_),
    .B(_07232_),
    .X(_07403_));
 sky130_fd_sc_hd__nor2_1 _14233_ (.A(_06914_),
    .B(_07193_),
    .Y(_07404_));
 sky130_fd_sc_hd__xnor2_2 _14234_ (.A(_07403_),
    .B(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__or3_1 _14235_ (.A(_07242_),
    .B(_07194_),
    .C(_07403_),
    .X(_07406_));
 sky130_fd_sc_hd__a21boi_4 _14236_ (.A1(_07402_),
    .A2(_07405_),
    .B1_N(_07406_),
    .Y(_07407_));
 sky130_fd_sc_hd__o21a_1 _14237_ (.A1(_07401_),
    .A2(_07407_),
    .B1(_07399_),
    .X(_07408_));
 sky130_fd_sc_hd__xor2_1 _14238_ (.A(_07395_),
    .B(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__xnor2_1 _14239_ (.A(_07394_),
    .B(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__xnor2_1 _14240_ (.A(_07374_),
    .B(_07375_),
    .Y(_07411_));
 sky130_fd_sc_hd__xor2_4 _14241_ (.A(_07401_),
    .B(_07407_),
    .X(_07412_));
 sky130_fd_sc_hd__clkbuf_4 _14242_ (.A(_06755_),
    .X(_07413_));
 sky130_fd_sc_hd__xor2_1 _14243_ (.A(_07310_),
    .B(_07344_),
    .X(_07414_));
 sky130_fd_sc_hd__o211a_1 _14244_ (.A1(_07413_),
    .A2(_07360_),
    .B1(_07414_),
    .C1(net5902),
    .X(_07415_));
 sky130_fd_sc_hd__nor2_2 _14245_ (.A(_07284_),
    .B(_07281_),
    .Y(_07416_));
 sky130_fd_sc_hd__xnor2_4 _14246_ (.A(_07310_),
    .B(_07416_),
    .Y(_07417_));
 sky130_fd_sc_hd__and3b_1 _14247_ (.A_N(net569),
    .B(_06758_),
    .C(_06759_),
    .X(_07418_));
 sky130_fd_sc_hd__nor2_1 _14248_ (.A(_07413_),
    .B(_07305_),
    .Y(_07419_));
 sky130_fd_sc_hd__a21oi_1 _14249_ (.A1(_06758_),
    .A2(_07342_),
    .B1(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__nor2_2 _14250_ (.A(_07418_),
    .B(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__a21oi_1 _14251_ (.A1(_07417_),
    .A2(_07421_),
    .B1(_07418_),
    .Y(_07422_));
 sky130_fd_sc_hd__nand2_1 _14252_ (.A(_07415_),
    .B(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__nor2_1 _14253_ (.A(_07415_),
    .B(_07422_),
    .Y(_07424_));
 sky130_fd_sc_hd__a21oi_2 _14254_ (.A1(_07412_),
    .A2(_07423_),
    .B1(_07424_),
    .Y(_07425_));
 sky130_fd_sc_hd__xor2_1 _14255_ (.A(_07411_),
    .B(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__nor2_1 _14256_ (.A(_07411_),
    .B(_07425_),
    .Y(_07427_));
 sky130_fd_sc_hd__a21oi_1 _14257_ (.A1(_07410_),
    .A2(_07426_),
    .B1(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__xnor2_1 _14258_ (.A(_07385_),
    .B(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__or2b_1 _14259_ (.A(_07394_),
    .B_N(_07409_),
    .X(_07430_));
 sky130_fd_sc_hd__o21ai_1 _14260_ (.A1(_07395_),
    .A2(_07408_),
    .B1(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__or2b_1 _14261_ (.A(_07429_),
    .B_N(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__o21a_1 _14262_ (.A1(_07385_),
    .A2(_07428_),
    .B1(_07432_),
    .X(_07433_));
 sky130_fd_sc_hd__nor2_2 _14263_ (.A(_07383_),
    .B(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__or2b_1 _14264_ (.A(_07237_),
    .B_N(_07354_),
    .X(_07435_));
 sky130_fd_sc_hd__o21ai_1 _14265_ (.A1(_07341_),
    .A2(_07353_),
    .B1(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__a211o_1 _14266_ (.A1(_07109_),
    .A2(_07342_),
    .B1(_07346_),
    .C1(_07363_),
    .X(_07437_));
 sky130_fd_sc_hd__a21bo_1 _14267_ (.A1(_07347_),
    .A2(_07363_),
    .B1_N(_07361_),
    .X(_07438_));
 sky130_fd_sc_hd__or3_2 _14268_ (.A(_07240_),
    .B(_07242_),
    .C(_07305_),
    .X(_07439_));
 sky130_fd_sc_hd__nand2_1 _14269_ (.A(_07438_),
    .B(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__a21o_1 _14270_ (.A1(_07437_),
    .A2(_07440_),
    .B1(net8355),
    .X(_07441_));
 sky130_fd_sc_hd__or2_1 _14271_ (.A(_06699_),
    .B(_07305_),
    .X(_07442_));
 sky130_fd_sc_hd__nor3b_1 _14272_ (.A(_06696_),
    .B(_07281_),
    .C_N(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__a21o_1 _14273_ (.A1(_07336_),
    .A2(_07337_),
    .B1(_07290_),
    .X(_07444_));
 sky130_fd_sc_hd__o21a_1 _14274_ (.A1(_07443_),
    .A2(_07444_),
    .B1(_07339_),
    .X(_07445_));
 sky130_fd_sc_hd__xnor2_1 _14275_ (.A(_07441_),
    .B(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__o21a_1 _14276_ (.A1(_07359_),
    .A2(_07366_),
    .B1(_07368_),
    .X(_07447_));
 sky130_fd_sc_hd__xnor2_1 _14277_ (.A(_07446_),
    .B(_07447_),
    .Y(_07448_));
 sky130_fd_sc_hd__xor2_1 _14278_ (.A(_07436_),
    .B(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__a21oi_1 _14279_ (.A1(_07334_),
    .A2(_07382_),
    .B1(_07380_),
    .Y(_07450_));
 sky130_fd_sc_hd__nor2_1 _14280_ (.A(_07449_),
    .B(_07450_),
    .Y(_07451_));
 sky130_fd_sc_hd__and2_1 _14281_ (.A(_07449_),
    .B(_07450_),
    .X(_07452_));
 sky130_fd_sc_hd__nor2_1 _14282_ (.A(_07451_),
    .B(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__xor2_2 _14283_ (.A(_07434_),
    .B(_07453_),
    .X(_07454_));
 sky130_fd_sc_hd__xor2_1 _14284_ (.A(_07431_),
    .B(_07429_),
    .X(_07455_));
 sky130_fd_sc_hd__xnor2_1 _14285_ (.A(_07410_),
    .B(_07426_),
    .Y(_07456_));
 sky130_fd_sc_hd__clkbuf_4 _14286_ (.A(_07145_),
    .X(_07457_));
 sky130_fd_sc_hd__or2_1 _14287_ (.A(_06696_),
    .B(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__nor3_2 _14288_ (.A(_06699_),
    .B(_07391_),
    .C(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__xnor2_2 _14289_ (.A(_07388_),
    .B(_07392_),
    .Y(_07460_));
 sky130_fd_sc_hd__nand2_2 _14290_ (.A(_07459_),
    .B(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__or3_1 _14291_ (.A(net8355),
    .B(_07393_),
    .C(_07387_),
    .X(_07462_));
 sky130_fd_sc_hd__nand2_1 _14292_ (.A(_07394_),
    .B(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__or4_4 _14293_ (.A(_07306_),
    .B(_06796_),
    .C(_07303_),
    .D(_07280_),
    .X(_07464_));
 sky130_fd_sc_hd__o22ai_1 _14294_ (.A1(_07306_),
    .A2(_07304_),
    .B1(_07280_),
    .B2(_07308_),
    .Y(_07465_));
 sky130_fd_sc_hd__nor2_1 _14295_ (.A(_06832_),
    .B(_07233_),
    .Y(_07466_));
 sky130_fd_sc_hd__nand3_1 _14296_ (.A(_07464_),
    .B(_07465_),
    .C(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__xnor2_1 _14297_ (.A(_07402_),
    .B(_07405_),
    .Y(_07468_));
 sky130_fd_sc_hd__a21o_1 _14298_ (.A1(_07464_),
    .A2(_07467_),
    .B1(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__nand3_1 _14299_ (.A(_07464_),
    .B(_07467_),
    .C(_07468_),
    .Y(_07470_));
 sky130_fd_sc_hd__nand2_2 _14300_ (.A(_07469_),
    .B(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nor2_1 _14301_ (.A(_07240_),
    .B(_07326_),
    .Y(_07472_));
 sky130_fd_sc_hd__or2_1 _14302_ (.A(_07033_),
    .B(_07193_),
    .X(_07473_));
 sky130_fd_sc_hd__nor2_1 _14303_ (.A(_06914_),
    .B(_07197_),
    .Y(_07474_));
 sky130_fd_sc_hd__xnor2_2 _14304_ (.A(_07473_),
    .B(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__or3_1 _14305_ (.A(_07242_),
    .B(_07198_),
    .C(_07473_),
    .X(_07476_));
 sky130_fd_sc_hd__a21boi_4 _14306_ (.A1(_07472_),
    .A2(_07475_),
    .B1_N(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__o21a_1 _14307_ (.A1(_07471_),
    .A2(_07477_),
    .B1(_07469_),
    .X(_07478_));
 sky130_fd_sc_hd__nor2_1 _14308_ (.A(_07463_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__and2_1 _14309_ (.A(_07463_),
    .B(_07478_),
    .X(_07480_));
 sky130_fd_sc_hd__nor2_2 _14310_ (.A(_07479_),
    .B(_07480_),
    .Y(_07481_));
 sky130_fd_sc_hd__xnor2_4 _14311_ (.A(_07461_),
    .B(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__and2b_1 _14312_ (.A_N(_07424_),
    .B(_07423_),
    .X(_07483_));
 sky130_fd_sc_hd__xnor2_4 _14313_ (.A(_07412_),
    .B(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__xor2_4 _14314_ (.A(_07471_),
    .B(_07477_),
    .X(_07485_));
 sky130_fd_sc_hd__xnor2_4 _14315_ (.A(_07417_),
    .B(_07421_),
    .Y(_07486_));
 sky130_fd_sc_hd__a21o_1 _14316_ (.A1(_07464_),
    .A2(_07465_),
    .B1(_07466_),
    .X(_07487_));
 sky130_fd_sc_hd__and2_4 _14317_ (.A(_07467_),
    .B(_07487_),
    .X(_07488_));
 sky130_fd_sc_hd__clkbuf_4 _14318_ (.A(_06754_),
    .X(_07489_));
 sky130_fd_sc_hd__a2bb2o_1 _14319_ (.A1_N(_07489_),
    .A2_N(_07305_),
    .B1(_07342_),
    .B2(_06931_),
    .X(_07490_));
 sky130_fd_sc_hd__or3_1 _14320_ (.A(_07072_),
    .B(_06754_),
    .C(_07303_),
    .X(_07491_));
 sky130_fd_sc_hd__or3_4 _14321_ (.A(_06924_),
    .B(_06755_),
    .C(_07303_),
    .X(_07492_));
 sky130_fd_sc_hd__a21o_1 _14322_ (.A1(_07491_),
    .A2(_07492_),
    .B1(_07418_),
    .X(_07493_));
 sky130_fd_sc_hd__o21a_4 _14323_ (.A1(_07419_),
    .A2(_07490_),
    .B1(_07493_),
    .X(_07494_));
 sky130_fd_sc_hd__a21boi_4 _14324_ (.A1(_07488_),
    .A2(_07494_),
    .B1_N(_07493_),
    .Y(_07495_));
 sky130_fd_sc_hd__xor2_4 _14325_ (.A(_07486_),
    .B(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__nor2_1 _14326_ (.A(_07486_),
    .B(_07495_),
    .Y(_07497_));
 sky130_fd_sc_hd__a21oi_4 _14327_ (.A1(_07485_),
    .A2(_07496_),
    .B1(_07497_),
    .Y(_07498_));
 sky130_fd_sc_hd__xor2_4 _14328_ (.A(_07484_),
    .B(_07498_),
    .X(_07499_));
 sky130_fd_sc_hd__nor2_1 _14329_ (.A(_07484_),
    .B(_07498_),
    .Y(_07500_));
 sky130_fd_sc_hd__a21oi_1 _14330_ (.A1(_07482_),
    .A2(_07499_),
    .B1(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__xnor2_1 _14331_ (.A(_07456_),
    .B(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__a31o_1 _14332_ (.A1(_07459_),
    .A2(_07460_),
    .A3(_07481_),
    .B1(_07479_),
    .X(_07503_));
 sky130_fd_sc_hd__or2b_1 _14333_ (.A(_07502_),
    .B_N(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__o21a_1 _14334_ (.A1(_07456_),
    .A2(_07501_),
    .B1(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__nor2_1 _14335_ (.A(_07455_),
    .B(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__and2_1 _14336_ (.A(_07383_),
    .B(_07433_),
    .X(_07507_));
 sky130_fd_sc_hd__nor2_2 _14337_ (.A(_07434_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__and2_1 _14338_ (.A(_07506_),
    .B(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__xor2_2 _14339_ (.A(_07454_),
    .B(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__inv_2 _14340_ (.A(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__xor2_1 _14341_ (.A(_07503_),
    .B(_07502_),
    .X(_07512_));
 sky130_fd_sc_hd__nor2_1 _14342_ (.A(_07308_),
    .B(_07233_),
    .Y(_07513_));
 sky130_fd_sc_hd__or3b_4 _14343_ (.A(_07306_),
    .B(_07280_),
    .C_N(_07513_),
    .X(_07514_));
 sky130_fd_sc_hd__o21bai_1 _14344_ (.A1(_07306_),
    .A2(_07281_),
    .B1_N(_07513_),
    .Y(_07515_));
 sky130_fd_sc_hd__nor2_1 _14345_ (.A(_06832_),
    .B(_07194_),
    .Y(_07516_));
 sky130_fd_sc_hd__nand3_1 _14346_ (.A(_07514_),
    .B(_07515_),
    .C(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__xnor2_1 _14347_ (.A(_07472_),
    .B(_07475_),
    .Y(_07518_));
 sky130_fd_sc_hd__a21o_1 _14348_ (.A1(_07514_),
    .A2(_07517_),
    .B1(_07518_),
    .X(_07519_));
 sky130_fd_sc_hd__nand3_1 _14349_ (.A(_07514_),
    .B(_07517_),
    .C(_07518_),
    .Y(_07520_));
 sky130_fd_sc_hd__nand2_2 _14350_ (.A(_07519_),
    .B(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__nor2_1 _14351_ (.A(_07240_),
    .B(_07390_),
    .Y(_07522_));
 sky130_fd_sc_hd__or2_1 _14352_ (.A(_07033_),
    .B(_07197_),
    .X(_07523_));
 sky130_fd_sc_hd__nor2_1 _14353_ (.A(_07242_),
    .B(_07326_),
    .Y(_07524_));
 sky130_fd_sc_hd__xnor2_2 _14354_ (.A(_07523_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__or3_1 _14355_ (.A(_07242_),
    .B(_07327_),
    .C(_07523_),
    .X(_07526_));
 sky130_fd_sc_hd__a21boi_4 _14356_ (.A1(_07522_),
    .A2(_07525_),
    .B1_N(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__or2_1 _14357_ (.A(_07521_),
    .B(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__or2_1 _14358_ (.A(_07459_),
    .B(_07460_),
    .X(_07529_));
 sky130_fd_sc_hd__nand2_1 _14359_ (.A(_07461_),
    .B(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__a21oi_4 _14360_ (.A1(_07519_),
    .A2(_07528_),
    .B1(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__xnor2_4 _14361_ (.A(_07482_),
    .B(_07499_),
    .Y(_07532_));
 sky130_fd_sc_hd__and3_1 _14362_ (.A(_07519_),
    .B(_07528_),
    .C(_07530_),
    .X(_07533_));
 sky130_fd_sc_hd__nor2_2 _14363_ (.A(_07531_),
    .B(_07533_),
    .Y(_07534_));
 sky130_fd_sc_hd__xnor2_4 _14364_ (.A(_07485_),
    .B(_07496_),
    .Y(_07535_));
 sky130_fd_sc_hd__xor2_4 _14365_ (.A(_07521_),
    .B(_07527_),
    .X(_07536_));
 sky130_fd_sc_hd__xnor2_4 _14366_ (.A(_07488_),
    .B(_07494_),
    .Y(_07537_));
 sky130_fd_sc_hd__a21oi_2 _14367_ (.A1(_06924_),
    .A2(_07413_),
    .B1(net569),
    .Y(_07538_));
 sky130_fd_sc_hd__nor2_1 _14368_ (.A(_06924_),
    .B(_07304_),
    .Y(_07539_));
 sky130_fd_sc_hd__nor2_1 _14369_ (.A(_07413_),
    .B(_07280_),
    .Y(_07540_));
 sky130_fd_sc_hd__a21bo_2 _14370_ (.A1(_07539_),
    .A2(_07540_),
    .B1_N(_07491_),
    .X(_07541_));
 sky130_fd_sc_hd__a21o_1 _14371_ (.A1(_07514_),
    .A2(_07515_),
    .B1(_07516_),
    .X(_07542_));
 sky130_fd_sc_hd__and2_2 _14372_ (.A(_07517_),
    .B(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__nand2_2 _14373_ (.A(_07492_),
    .B(_07538_),
    .Y(_07544_));
 sky130_fd_sc_hd__xnor2_4 _14374_ (.A(_07544_),
    .B(_07541_),
    .Y(_07545_));
 sky130_fd_sc_hd__a32oi_4 _14375_ (.A1(_07492_),
    .A2(_07538_),
    .A3(_07541_),
    .B1(_07543_),
    .B2(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__xor2_4 _14376_ (.A(_07537_),
    .B(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__or2_1 _14377_ (.A(_07537_),
    .B(_07546_),
    .X(_07548_));
 sky130_fd_sc_hd__a21boi_4 _14378_ (.A1(_07536_),
    .A2(_07547_),
    .B1_N(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__xor2_4 _14379_ (.A(_07535_),
    .B(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__nor2_1 _14380_ (.A(_07535_),
    .B(_07549_),
    .Y(_07551_));
 sky130_fd_sc_hd__a21oi_4 _14381_ (.A1(_07534_),
    .A2(_07550_),
    .B1(_07551_),
    .Y(_07552_));
 sky130_fd_sc_hd__xor2_4 _14382_ (.A(_07532_),
    .B(_07552_),
    .X(_07553_));
 sky130_fd_sc_hd__nor2_1 _14383_ (.A(_07532_),
    .B(_07552_),
    .Y(_07554_));
 sky130_fd_sc_hd__a21oi_1 _14384_ (.A1(_07531_),
    .A2(_07553_),
    .B1(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__nor2_1 _14385_ (.A(_07512_),
    .B(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__and2_1 _14386_ (.A(_07455_),
    .B(_07505_),
    .X(_07557_));
 sky130_fd_sc_hd__nor2_1 _14387_ (.A(_07506_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__and2_1 _14388_ (.A(_07556_),
    .B(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__xnor2_4 _14389_ (.A(_07531_),
    .B(_07553_),
    .Y(_07560_));
 sky130_fd_sc_hd__or2_1 _14390_ (.A(_06771_),
    .B(_07232_),
    .X(_07561_));
 sky130_fd_sc_hd__or3_1 _14391_ (.A(_07308_),
    .B(_07194_),
    .C(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__nor2_1 _14392_ (.A(_07308_),
    .B(_07193_),
    .Y(_07563_));
 sky130_fd_sc_hd__xnor2_1 _14393_ (.A(_07561_),
    .B(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__nor2_1 _14394_ (.A(_07284_),
    .B(_07198_),
    .Y(_07565_));
 sky130_fd_sc_hd__nand2_1 _14395_ (.A(_07564_),
    .B(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__xnor2_1 _14396_ (.A(_07522_),
    .B(_07525_),
    .Y(_07567_));
 sky130_fd_sc_hd__a21o_1 _14397_ (.A1(_07562_),
    .A2(_07566_),
    .B1(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__nand3_1 _14398_ (.A(_07562_),
    .B(_07566_),
    .C(_07567_),
    .Y(_07569_));
 sky130_fd_sc_hd__nand2_1 _14399_ (.A(_07568_),
    .B(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__or2_1 _14400_ (.A(_07033_),
    .B(_07326_),
    .X(_07571_));
 sky130_fd_sc_hd__nor2_1 _14401_ (.A(_07240_),
    .B(_07145_),
    .Y(_07572_));
 sky130_fd_sc_hd__nor2_1 _14402_ (.A(_06914_),
    .B(_07390_),
    .Y(_07573_));
 sky130_fd_sc_hd__xnor2_1 _14403_ (.A(_07571_),
    .B(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__nand2_1 _14404_ (.A(_07572_),
    .B(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__o31a_1 _14405_ (.A1(_07242_),
    .A2(_07391_),
    .A3(_07571_),
    .B1(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__or2_1 _14406_ (.A(_07570_),
    .B(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__o21a_1 _14407_ (.A1(_06699_),
    .A2(_07391_),
    .B1(_07458_),
    .X(_07578_));
 sky130_fd_sc_hd__or2_1 _14408_ (.A(_07459_),
    .B(_07578_),
    .X(_07579_));
 sky130_fd_sc_hd__a21oi_2 _14409_ (.A1(_07568_),
    .A2(_07577_),
    .B1(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__xnor2_2 _14410_ (.A(_07534_),
    .B(_07550_),
    .Y(_07581_));
 sky130_fd_sc_hd__and3_1 _14411_ (.A(_07568_),
    .B(_07577_),
    .C(_07579_),
    .X(_07582_));
 sky130_fd_sc_hd__nor2_1 _14412_ (.A(_07580_),
    .B(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__xnor2_2 _14413_ (.A(_07536_),
    .B(_07547_),
    .Y(_07584_));
 sky130_fd_sc_hd__xor2_2 _14414_ (.A(_07570_),
    .B(_07576_),
    .X(_07585_));
 sky130_fd_sc_hd__xnor2_2 _14415_ (.A(_07543_),
    .B(_07545_),
    .Y(_07586_));
 sky130_fd_sc_hd__or2_1 _14416_ (.A(_07564_),
    .B(_07565_),
    .X(_07587_));
 sky130_fd_sc_hd__and2_1 _14417_ (.A(_07566_),
    .B(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__xnor2_2 _14418_ (.A(_07539_),
    .B(_07540_),
    .Y(_07589_));
 sky130_fd_sc_hd__nor2_1 _14419_ (.A(_07413_),
    .B(_07233_),
    .Y(_07590_));
 sky130_fd_sc_hd__o22ai_2 _14420_ (.A1(_07072_),
    .A2(net569),
    .B1(_07281_),
    .B2(_06754_),
    .Y(_07591_));
 sky130_fd_sc_hd__or4_4 _14421_ (.A(_07072_),
    .B(_06754_),
    .C(_07304_),
    .D(_07280_),
    .X(_07592_));
 sky130_fd_sc_hd__a21bo_4 _14422_ (.A1(_07590_),
    .A2(_07591_),
    .B1_N(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__xnor2_2 _14423_ (.A(_07589_),
    .B(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__and2b_1 _14424_ (.A_N(_07589_),
    .B(_07593_),
    .X(_07595_));
 sky130_fd_sc_hd__a21oi_2 _14425_ (.A1(_07588_),
    .A2(_07594_),
    .B1(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__xor2_2 _14426_ (.A(_07586_),
    .B(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__nor2_1 _14427_ (.A(_07586_),
    .B(_07596_),
    .Y(_07598_));
 sky130_fd_sc_hd__a21oi_2 _14428_ (.A1(_07585_),
    .A2(_07597_),
    .B1(_07598_),
    .Y(_07599_));
 sky130_fd_sc_hd__xor2_2 _14429_ (.A(_07584_),
    .B(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__nor2_1 _14430_ (.A(_07584_),
    .B(_07599_),
    .Y(_07601_));
 sky130_fd_sc_hd__a21oi_2 _14431_ (.A1(_07583_),
    .A2(_07600_),
    .B1(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__xor2_2 _14432_ (.A(_07581_),
    .B(_07602_),
    .X(_07603_));
 sky130_fd_sc_hd__nor2_1 _14433_ (.A(_07581_),
    .B(_07602_),
    .Y(_07604_));
 sky130_fd_sc_hd__a21oi_2 _14434_ (.A1(_07580_),
    .A2(_07603_),
    .B1(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__nor2_1 _14435_ (.A(_07560_),
    .B(_07605_),
    .Y(_07606_));
 sky130_fd_sc_hd__and2_1 _14436_ (.A(_07512_),
    .B(_07555_),
    .X(_07607_));
 sky130_fd_sc_hd__nor2_2 _14437_ (.A(_07556_),
    .B(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__xor2_4 _14438_ (.A(_07560_),
    .B(_07605_),
    .X(_07609_));
 sky130_fd_sc_hd__xnor2_2 _14439_ (.A(_07580_),
    .B(_07603_),
    .Y(_07610_));
 sky130_fd_sc_hd__nor2_1 _14440_ (.A(_07308_),
    .B(_07197_),
    .Y(_07611_));
 sky130_fd_sc_hd__a31o_1 _14441_ (.A1(_06725_),
    .A2(_07191_),
    .A3(_07192_),
    .B1(_07611_),
    .X(_07612_));
 sky130_fd_sc_hd__nor2_1 _14442_ (.A(_07284_),
    .B(_07326_),
    .Y(_07613_));
 sky130_fd_sc_hd__or3b_1 _14443_ (.A(_07306_),
    .B(_07193_),
    .C_N(_07611_),
    .X(_07614_));
 sky130_fd_sc_hd__a21bo_1 _14444_ (.A1(_07612_),
    .A2(_07613_),
    .B1_N(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__xnor2_1 _14445_ (.A(_07572_),
    .B(_07574_),
    .Y(_07616_));
 sky130_fd_sc_hd__or2b_1 _14446_ (.A(_07615_),
    .B_N(_07616_),
    .X(_07617_));
 sky130_fd_sc_hd__nor2_1 _14447_ (.A(_07033_),
    .B(_07391_),
    .Y(_07618_));
 sky130_fd_sc_hd__nor2_1 _14448_ (.A(_07242_),
    .B(_07457_),
    .Y(_07619_));
 sky130_fd_sc_hd__and2_1 _14449_ (.A(_07618_),
    .B(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__and2b_1 _14450_ (.A_N(_07616_),
    .B(_07615_),
    .X(_07621_));
 sky130_fd_sc_hd__a21oi_1 _14451_ (.A1(_07617_),
    .A2(_07620_),
    .B1(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__nor2_1 _14452_ (.A(_06699_),
    .B(_07457_),
    .Y(_07623_));
 sky130_fd_sc_hd__nor2b_1 _14453_ (.A(_07622_),
    .B_N(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__xnor2_2 _14454_ (.A(_07583_),
    .B(_07600_),
    .Y(_07625_));
 sky130_fd_sc_hd__and2b_1 _14455_ (.A_N(_07623_),
    .B(_07622_),
    .X(_07626_));
 sky130_fd_sc_hd__nor2_1 _14456_ (.A(_07624_),
    .B(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__xnor2_2 _14457_ (.A(_07585_),
    .B(_07597_),
    .Y(_07628_));
 sky130_fd_sc_hd__or2b_1 _14458_ (.A(_07621_),
    .B_N(_07617_),
    .X(_07629_));
 sky130_fd_sc_hd__xnor2_1 _14459_ (.A(_07629_),
    .B(_07620_),
    .Y(_07630_));
 sky130_fd_sc_hd__xnor2_2 _14460_ (.A(_07588_),
    .B(_07594_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_1 _14461_ (.A(_07614_),
    .B(_07612_),
    .Y(_07632_));
 sky130_fd_sc_hd__xnor2_2 _14462_ (.A(_07632_),
    .B(_07613_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand3_1 _14463_ (.A(_07592_),
    .B(_07590_),
    .C(_07591_),
    .Y(_07634_));
 sky130_fd_sc_hd__a21o_1 _14464_ (.A1(_07592_),
    .A2(_07591_),
    .B1(_07590_),
    .X(_07635_));
 sky130_fd_sc_hd__nor2_1 _14465_ (.A(_07413_),
    .B(_07194_),
    .Y(_07636_));
 sky130_fd_sc_hd__o22ai_2 _14466_ (.A1(_07489_),
    .A2(_07233_),
    .B1(_07281_),
    .B2(_07072_),
    .Y(_07637_));
 sky130_fd_sc_hd__or4_1 _14467_ (.A(_07072_),
    .B(_06754_),
    .C(_07233_),
    .D(_07280_),
    .X(_07638_));
 sky130_fd_sc_hd__a21bo_1 _14468_ (.A1(_07636_),
    .A2(_07637_),
    .B1_N(_07638_),
    .X(_07639_));
 sky130_fd_sc_hd__a21o_1 _14469_ (.A1(_07634_),
    .A2(_07635_),
    .B1(_07639_),
    .X(_07640_));
 sky130_fd_sc_hd__nand3_1 _14470_ (.A(_07634_),
    .B(_07635_),
    .C(_07639_),
    .Y(_07641_));
 sky130_fd_sc_hd__a21boi_2 _14471_ (.A1(_07633_),
    .A2(_07640_),
    .B1_N(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__xor2_2 _14472_ (.A(_07631_),
    .B(_07642_),
    .X(_07643_));
 sky130_fd_sc_hd__nor2_1 _14473_ (.A(_07631_),
    .B(_07642_),
    .Y(_07644_));
 sky130_fd_sc_hd__a21oi_2 _14474_ (.A1(_07630_),
    .A2(_07643_),
    .B1(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__xor2_2 _14475_ (.A(_07628_),
    .B(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__nor2_1 _14476_ (.A(_07628_),
    .B(_07645_),
    .Y(_07647_));
 sky130_fd_sc_hd__a21oi_2 _14477_ (.A1(_07627_),
    .A2(_07646_),
    .B1(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__xor2_2 _14478_ (.A(_07625_),
    .B(_07648_),
    .X(_07649_));
 sky130_fd_sc_hd__nor2_1 _14479_ (.A(_07625_),
    .B(_07648_),
    .Y(_07650_));
 sky130_fd_sc_hd__a21oi_2 _14480_ (.A1(_07624_),
    .A2(_07649_),
    .B1(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__nor2_1 _14481_ (.A(_07610_),
    .B(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__and2_1 _14482_ (.A(_07609_),
    .B(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__nor2_1 _14483_ (.A(_07606_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__xnor2_2 _14484_ (.A(_07608_),
    .B(_07654_),
    .Y(_07655_));
 sky130_fd_sc_hd__xor2_2 _14485_ (.A(_07610_),
    .B(_07651_),
    .X(_07656_));
 sky130_fd_sc_hd__or2_1 _14486_ (.A(_07306_),
    .B(_07197_),
    .X(_07657_));
 sky130_fd_sc_hd__or3_1 _14487_ (.A(_07308_),
    .B(_07327_),
    .C(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__nor2_1 _14488_ (.A(_07308_),
    .B(_07326_),
    .Y(_07659_));
 sky130_fd_sc_hd__xnor2_1 _14489_ (.A(_07657_),
    .B(_07659_),
    .Y(_07660_));
 sky130_fd_sc_hd__nor2_1 _14490_ (.A(_07284_),
    .B(_07390_),
    .Y(_07661_));
 sky130_fd_sc_hd__nand2_1 _14491_ (.A(_07660_),
    .B(_07661_),
    .Y(_07662_));
 sky130_fd_sc_hd__nor2_1 _14492_ (.A(_07618_),
    .B(_07619_),
    .Y(_07663_));
 sky130_fd_sc_hd__or2_1 _14493_ (.A(_07620_),
    .B(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__a21oi_2 _14494_ (.A1(_07658_),
    .A2(_07662_),
    .B1(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__xnor2_1 _14495_ (.A(_07630_),
    .B(_07643_),
    .Y(_07666_));
 sky130_fd_sc_hd__and3_1 _14496_ (.A(_07658_),
    .B(_07662_),
    .C(_07664_),
    .X(_07667_));
 sky130_fd_sc_hd__nor2_1 _14497_ (.A(_07665_),
    .B(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__nand3_1 _14498_ (.A(_07641_),
    .B(_07633_),
    .C(_07640_),
    .Y(_07669_));
 sky130_fd_sc_hd__a21o_1 _14499_ (.A1(_07641_),
    .A2(_07640_),
    .B1(_07633_),
    .X(_07670_));
 sky130_fd_sc_hd__or2_1 _14500_ (.A(_07660_),
    .B(_07661_),
    .X(_07671_));
 sky130_fd_sc_hd__and2_1 _14501_ (.A(_07662_),
    .B(_07671_),
    .X(_07672_));
 sky130_fd_sc_hd__nand3_1 _14502_ (.A(_07638_),
    .B(_07636_),
    .C(_07637_),
    .Y(_07673_));
 sky130_fd_sc_hd__a21o_1 _14503_ (.A1(_07638_),
    .A2(_07637_),
    .B1(_07636_),
    .X(_07674_));
 sky130_fd_sc_hd__nor2_1 _14504_ (.A(_07413_),
    .B(_07198_),
    .Y(_07675_));
 sky130_fd_sc_hd__or2_1 _14505_ (.A(_07072_),
    .B(_07233_),
    .X(_07676_));
 sky130_fd_sc_hd__nor2_1 _14506_ (.A(_07489_),
    .B(_07194_),
    .Y(_07677_));
 sky130_fd_sc_hd__xnor2_1 _14507_ (.A(_07676_),
    .B(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__or3_1 _14508_ (.A(_07489_),
    .B(_07194_),
    .C(_07676_),
    .X(_07679_));
 sky130_fd_sc_hd__a21bo_1 _14509_ (.A1(_07675_),
    .A2(_07678_),
    .B1_N(_07679_),
    .X(_07680_));
 sky130_fd_sc_hd__a21o_1 _14510_ (.A1(_07673_),
    .A2(_07674_),
    .B1(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__and3_1 _14511_ (.A(_07673_),
    .B(_07674_),
    .C(_07680_),
    .X(_07682_));
 sky130_fd_sc_hd__a21o_1 _14512_ (.A1(_07672_),
    .A2(_07681_),
    .B1(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__a21o_1 _14513_ (.A1(_07669_),
    .A2(_07670_),
    .B1(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__and3_1 _14514_ (.A(_07669_),
    .B(_07670_),
    .C(_07683_),
    .X(_07685_));
 sky130_fd_sc_hd__a21oi_1 _14515_ (.A1(_07668_),
    .A2(_07684_),
    .B1(_07685_),
    .Y(_07686_));
 sky130_fd_sc_hd__nand2_1 _14516_ (.A(_07666_),
    .B(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__nor2_1 _14517_ (.A(_07666_),
    .B(_07686_),
    .Y(_07688_));
 sky130_fd_sc_hd__a21oi_1 _14518_ (.A1(_07665_),
    .A2(_07687_),
    .B1(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__xnor2_1 _14519_ (.A(_07627_),
    .B(_07646_),
    .Y(_07690_));
 sky130_fd_sc_hd__xor2_1 _14520_ (.A(_07624_),
    .B(_07649_),
    .X(_07691_));
 sky130_fd_sc_hd__nor3b_2 _14521_ (.A(_07689_),
    .B(_07690_),
    .C_N(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__and2_1 _14522_ (.A(_07656_),
    .B(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__xor2_1 _14523_ (.A(_07690_),
    .B(_07689_),
    .X(_07694_));
 sky130_fd_sc_hd__nand2_1 _14524_ (.A(_07691_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__xor2_2 _14525_ (.A(_07656_),
    .B(net76),
    .X(_07696_));
 sky130_fd_sc_hd__and2b_1 _14526_ (.A_N(_07688_),
    .B(_07687_),
    .X(_07697_));
 sky130_fd_sc_hd__xor2_1 _14527_ (.A(_07665_),
    .B(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__nor2_1 _14528_ (.A(_07306_),
    .B(_07327_),
    .Y(_07699_));
 sky130_fd_sc_hd__nor2_1 _14529_ (.A(_07308_),
    .B(_07391_),
    .Y(_07700_));
 sky130_fd_sc_hd__xnor2_1 _14530_ (.A(_07699_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__nand2_1 _14531_ (.A(_07699_),
    .B(_07700_),
    .Y(_07702_));
 sky130_fd_sc_hd__o31a_1 _14532_ (.A1(_07284_),
    .A2(_07457_),
    .A3(_07701_),
    .B1(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__or3_1 _14533_ (.A(_07033_),
    .B(_07457_),
    .C(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__o21ai_1 _14534_ (.A1(_07033_),
    .A2(_07457_),
    .B1(_07703_),
    .Y(_07705_));
 sky130_fd_sc_hd__and2_1 _14535_ (.A(_07704_),
    .B(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__and2b_1 _14536_ (.A_N(_07682_),
    .B(_07681_),
    .X(_07707_));
 sky130_fd_sc_hd__xnor2_1 _14537_ (.A(_07672_),
    .B(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__nor2_1 _14538_ (.A(_07284_),
    .B(_07457_),
    .Y(_07709_));
 sky130_fd_sc_hd__xnor2_1 _14539_ (.A(_07701_),
    .B(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__xnor2_1 _14540_ (.A(_07675_),
    .B(_07678_),
    .Y(_07711_));
 sky130_fd_sc_hd__nor2_1 _14541_ (.A(_07413_),
    .B(_07327_),
    .Y(_07712_));
 sky130_fd_sc_hd__or2_1 _14542_ (.A(_07072_),
    .B(_07194_),
    .X(_07713_));
 sky130_fd_sc_hd__nor2_1 _14543_ (.A(_07489_),
    .B(_07198_),
    .Y(_07714_));
 sky130_fd_sc_hd__xnor2_1 _14544_ (.A(_07713_),
    .B(_07714_),
    .Y(_07715_));
 sky130_fd_sc_hd__or3_1 _14545_ (.A(_07489_),
    .B(_07198_),
    .C(_07713_),
    .X(_07716_));
 sky130_fd_sc_hd__a21bo_1 _14546_ (.A1(_07712_),
    .A2(_07715_),
    .B1_N(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__xnor2_1 _14547_ (.A(_07711_),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__and2b_1 _14548_ (.A_N(_07711_),
    .B(_07717_),
    .X(_07719_));
 sky130_fd_sc_hd__a21oi_1 _14549_ (.A1(_07710_),
    .A2(_07718_),
    .B1(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__xor2_1 _14550_ (.A(_07708_),
    .B(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__nor2_1 _14551_ (.A(_07708_),
    .B(_07720_),
    .Y(_07722_));
 sky130_fd_sc_hd__a21oi_1 _14552_ (.A1(_07706_),
    .A2(_07721_),
    .B1(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__and2b_1 _14553_ (.A_N(_07685_),
    .B(_07684_),
    .X(_07724_));
 sky130_fd_sc_hd__xor2_1 _14554_ (.A(_07668_),
    .B(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__or2b_1 _14555_ (.A(_07723_),
    .B_N(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__or2b_1 _14556_ (.A(_07725_),
    .B_N(_07723_),
    .X(_07727_));
 sky130_fd_sc_hd__nand2_1 _14557_ (.A(_07726_),
    .B(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__or2_1 _14558_ (.A(_07704_),
    .B(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__nand2_1 _14559_ (.A(_07726_),
    .B(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__and4_1 _14560_ (.A(_07691_),
    .B(_07698_),
    .C(_07730_),
    .D(_07694_),
    .X(_07731_));
 sky130_fd_sc_hd__xnor2_2 _14561_ (.A(_07696_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__nand2_1 _14562_ (.A(_07704_),
    .B(_07728_),
    .Y(_07733_));
 sky130_fd_sc_hd__nor2_1 _14563_ (.A(_07306_),
    .B(_07391_),
    .Y(_07734_));
 sky130_fd_sc_hd__or2_1 _14564_ (.A(_07308_),
    .B(_07457_),
    .X(_07735_));
 sky130_fd_sc_hd__inv_2 _14565_ (.A(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__nand2_1 _14566_ (.A(_07734_),
    .B(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__or2_1 _14567_ (.A(_07734_),
    .B(_07736_),
    .X(_07738_));
 sky130_fd_sc_hd__nand2_1 _14568_ (.A(_07737_),
    .B(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__xnor2_1 _14569_ (.A(_07712_),
    .B(_07715_),
    .Y(_07740_));
 sky130_fd_sc_hd__nor2_1 _14570_ (.A(_07413_),
    .B(_07391_),
    .Y(_07741_));
 sky130_fd_sc_hd__or2_1 _14571_ (.A(_07072_),
    .B(_07198_),
    .X(_07742_));
 sky130_fd_sc_hd__nor2_1 _14572_ (.A(_07489_),
    .B(_07327_),
    .Y(_07743_));
 sky130_fd_sc_hd__xnor2_1 _14573_ (.A(_07742_),
    .B(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__or3_1 _14574_ (.A(_07489_),
    .B(_07327_),
    .C(_07742_),
    .X(_07745_));
 sky130_fd_sc_hd__a21boi_1 _14575_ (.A1(_07741_),
    .A2(_07744_),
    .B1_N(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__nor2_1 _14576_ (.A(_07740_),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__and2_1 _14577_ (.A(_07740_),
    .B(_07746_),
    .X(_07748_));
 sky130_fd_sc_hd__nor2_1 _14578_ (.A(_07747_),
    .B(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__xnor2_1 _14579_ (.A(_07739_),
    .B(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__xnor2_1 _14580_ (.A(_07741_),
    .B(_07744_),
    .Y(_07751_));
 sky130_fd_sc_hd__or2_1 _14581_ (.A(_07072_),
    .B(_07327_),
    .X(_07752_));
 sky130_fd_sc_hd__nor2_1 _14582_ (.A(_07413_),
    .B(_07457_),
    .Y(_07753_));
 sky130_fd_sc_hd__nor2_1 _14583_ (.A(_07489_),
    .B(_07391_),
    .Y(_07754_));
 sky130_fd_sc_hd__xnor2_1 _14584_ (.A(_07752_),
    .B(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__nand2_1 _14585_ (.A(_07753_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__o31a_1 _14586_ (.A1(_07489_),
    .A2(_07391_),
    .A3(_07752_),
    .B1(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__nor2_1 _14587_ (.A(_07306_),
    .B(_07457_),
    .Y(_07758_));
 sky130_fd_sc_hd__xor2_1 _14588_ (.A(_07751_),
    .B(_07757_),
    .X(_07759_));
 sky130_fd_sc_hd__nand2_1 _14589_ (.A(_07758_),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__o21ai_1 _14590_ (.A1(_07751_),
    .A2(_07757_),
    .B1(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__nand2_1 _14591_ (.A(_07750_),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__and3_1 _14592_ (.A(net77),
    .B(_07146_),
    .C(_07756_),
    .X(_07763_));
 sky130_fd_sc_hd__o211a_1 _14593_ (.A1(_07753_),
    .A2(_07755_),
    .B1(_07760_),
    .C1(_07763_),
    .X(_07764_));
 sky130_fd_sc_hd__o221ai_2 _14594_ (.A1(_07758_),
    .A2(_07759_),
    .B1(_07761_),
    .B2(_07750_),
    .C1(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__o21ba_1 _14595_ (.A1(_07739_),
    .A2(_07748_),
    .B1_N(_07747_),
    .X(_07766_));
 sky130_fd_sc_hd__xnor2_1 _14596_ (.A(_07710_),
    .B(_07718_),
    .Y(_07767_));
 sky130_fd_sc_hd__a32oi_1 _14597_ (.A1(_07737_),
    .A2(_07762_),
    .A3(_07765_),
    .B1(_07766_),
    .B2(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__nor2_1 _14598_ (.A(_07767_),
    .B(_07766_),
    .Y(_07769_));
 sky130_fd_sc_hd__a21oi_1 _14599_ (.A1(_07762_),
    .A2(_07765_),
    .B1(_07737_),
    .Y(_07770_));
 sky130_fd_sc_hd__or3_1 _14600_ (.A(_07768_),
    .B(_07769_),
    .C(_07770_),
    .X(_07771_));
 sky130_fd_sc_hd__xor2_1 _14601_ (.A(_07706_),
    .B(_07721_),
    .X(_07772_));
 sky130_fd_sc_hd__and4_1 _14602_ (.A(_07729_),
    .B(_07733_),
    .C(_07771_),
    .D(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__o21ai_2 _14603_ (.A1(_07698_),
    .A2(_07730_),
    .B1(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__nand2_1 _14604_ (.A(_07696_),
    .B(_07731_),
    .Y(_07775_));
 sky130_fd_sc_hd__o31ai_4 _14605_ (.A1(_07695_),
    .A2(_07732_),
    .A3(_07774_),
    .B1(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__nor2_2 _14606_ (.A(_07652_),
    .B(_07693_),
    .Y(_07777_));
 sky130_fd_sc_hd__xnor2_4 _14607_ (.A(_07609_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__a22o_1 _14608_ (.A1(_07609_),
    .A2(_07693_),
    .B1(_07776_),
    .B2(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__a22o_1 _14609_ (.A1(_07608_),
    .A2(_07653_),
    .B1(_07655_),
    .B2(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__a21o_1 _14610_ (.A1(_07606_),
    .A2(_07608_),
    .B1(_07556_),
    .X(_07781_));
 sky130_fd_sc_hd__xnor2_1 _14611_ (.A(_07558_),
    .B(_07781_),
    .Y(_07782_));
 sky130_fd_sc_hd__inv_2 _14612_ (.A(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__a32o_2 _14613_ (.A1(_07558_),
    .A2(_07606_),
    .A3(_07608_),
    .B1(_07780_),
    .B2(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__nor2_1 _14614_ (.A(_07506_),
    .B(_07559_),
    .Y(_07785_));
 sky130_fd_sc_hd__xnor2_2 _14615_ (.A(_07508_),
    .B(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__a22oi_4 _14616_ (.A1(_07508_),
    .A2(_07559_),
    .B1(_07784_),
    .B2(_07786_),
    .Y(_07787_));
 sky130_fd_sc_hd__and2_1 _14617_ (.A(_07454_),
    .B(_07509_),
    .X(_07788_));
 sky130_fd_sc_hd__o21bai_4 _14618_ (.A1(_07511_),
    .A2(_07787_),
    .B1_N(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__and2_2 _14619_ (.A(_07434_),
    .B(_07453_),
    .X(_07790_));
 sky130_fd_sc_hd__a21o_1 _14620_ (.A1(_07251_),
    .A2(_07342_),
    .B1(_07363_),
    .X(_07791_));
 sky130_fd_sc_hd__and3b_1 _14621_ (.A_N(_07305_),
    .B(_07339_),
    .C(_07440_),
    .X(_07792_));
 sky130_fd_sc_hd__a21oi_1 _14622_ (.A1(_07439_),
    .A2(_07791_),
    .B1(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__nand3_1 _14623_ (.A(_07439_),
    .B(_07792_),
    .C(_07791_),
    .Y(_07794_));
 sky130_fd_sc_hd__and3_1 _14624_ (.A(_07441_),
    .B(_07445_),
    .C(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__o21a_1 _14625_ (.A1(_07793_),
    .A2(_07795_),
    .B1(_07339_),
    .X(_07796_));
 sky130_fd_sc_hd__or2b_1 _14626_ (.A(_07448_),
    .B_N(_07436_),
    .X(_07797_));
 sky130_fd_sc_hd__o21a_1 _14627_ (.A1(_07446_),
    .A2(_07447_),
    .B1(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__xor2_1 _14628_ (.A(_07796_),
    .B(_07798_),
    .X(_07799_));
 sky130_fd_sc_hd__and2_1 _14629_ (.A(_07451_),
    .B(_07799_),
    .X(_07800_));
 sky130_fd_sc_hd__nor2_1 _14630_ (.A(_07451_),
    .B(_07799_),
    .Y(_07801_));
 sky130_fd_sc_hd__nor2_2 _14631_ (.A(_07800_),
    .B(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__xnor2_4 _14632_ (.A(_07790_),
    .B(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__xnor2_4 _14633_ (.A(_07789_),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__nor2_1 _14634_ (.A(_07796_),
    .B(_07798_),
    .Y(_07805_));
 sky130_fd_sc_hd__a21oi_1 _14635_ (.A1(_06839_),
    .A2(_07251_),
    .B1(_07305_),
    .Y(_07806_));
 sky130_fd_sc_hd__nor2_1 _14636_ (.A(_07240_),
    .B(_07360_),
    .Y(_07807_));
 sky130_fd_sc_hd__and2_1 _14637_ (.A(_07440_),
    .B(_07794_),
    .X(_07808_));
 sky130_fd_sc_hd__o31a_1 _14638_ (.A1(net8355),
    .A2(_07806_),
    .A3(_07807_),
    .B1(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__xor2_2 _14639_ (.A(_07795_),
    .B(_07809_),
    .X(_07810_));
 sky130_fd_sc_hd__xor2_1 _14640_ (.A(_07805_),
    .B(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__nand2_1 _14641_ (.A(_07800_),
    .B(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__or2_1 _14642_ (.A(_07800_),
    .B(_07811_),
    .X(_07813_));
 sky130_fd_sc_hd__and2_1 _14643_ (.A(_07812_),
    .B(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__o21ai_1 _14644_ (.A1(_07790_),
    .A2(_07788_),
    .B1(_07802_),
    .Y(_07815_));
 sky130_fd_sc_hd__o31a_1 _14645_ (.A1(_07511_),
    .A2(_07787_),
    .A3(_07803_),
    .B1(_07815_),
    .X(_07816_));
 sky130_fd_sc_hd__xnor2_1 _14646_ (.A(_07814_),
    .B(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__buf_2 _14647_ (.A(net7807),
    .X(_07818_));
 sky130_fd_sc_hd__mux2_1 _14648_ (.A0(_07804_),
    .A1(_07817_),
    .S(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__or2_1 _14649_ (.A(net7811),
    .B(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__buf_2 _14650_ (.A(net7795),
    .X(_07821_));
 sky130_fd_sc_hd__nand2_2 _14651_ (.A(_07805_),
    .B(_07810_),
    .Y(_07822_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(_06699_),
    .A1(_07807_),
    .S(_07305_),
    .X(_07823_));
 sky130_fd_sc_hd__o21ai_1 _14653_ (.A1(net8355),
    .A2(_07823_),
    .B1(_07439_),
    .Y(_07824_));
 sky130_fd_sc_hd__a2bb2o_1 _14654_ (.A1_N(_07808_),
    .A2_N(_07824_),
    .B1(_07809_),
    .B2(_07795_),
    .X(_07825_));
 sky130_fd_sc_hd__a21o_2 _14655_ (.A1(_07808_),
    .A2(_07824_),
    .B1(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__xor2_4 _14656_ (.A(_07822_),
    .B(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__inv_2 _14657_ (.A(_07814_),
    .Y(_07828_));
 sky130_fd_sc_hd__o21a_1 _14658_ (.A1(_07828_),
    .A2(_07816_),
    .B1(_07812_),
    .X(_07829_));
 sky130_fd_sc_hd__xnor2_4 _14659_ (.A(_07827_),
    .B(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__nand2_1 _14660_ (.A(_07814_),
    .B(_07827_),
    .Y(_07831_));
 sky130_fd_sc_hd__or4_4 _14661_ (.A(_07511_),
    .B(_07787_),
    .C(_07803_),
    .D(_07831_),
    .X(_07832_));
 sky130_fd_sc_hd__a21o_1 _14662_ (.A1(_07822_),
    .A2(_07812_),
    .B1(_07826_),
    .X(_07833_));
 sky130_fd_sc_hd__o21a_1 _14663_ (.A1(_07815_),
    .A2(_07831_),
    .B1(_07833_),
    .X(_07834_));
 sky130_fd_sc_hd__o211a_1 _14664_ (.A1(_06696_),
    .A2(_07360_),
    .B1(_07442_),
    .C1(net8491),
    .X(_07835_));
 sky130_fd_sc_hd__and3b_1 _14665_ (.A_N(_07825_),
    .B(_07835_),
    .C(_07439_),
    .X(_07836_));
 sky130_fd_sc_hd__a21o_1 _14666_ (.A1(_07832_),
    .A2(_07834_),
    .B1(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__nand3_1 _14667_ (.A(net564),
    .B(_07834_),
    .C(_07836_),
    .Y(_07838_));
 sky130_fd_sc_hd__and3_4 _14668_ (.A(net7807),
    .B(_07837_),
    .C(_07838_),
    .X(_07839_));
 sky130_fd_sc_hd__clkbuf_1 _14669_ (.A(net7842),
    .X(_07840_));
 sky130_fd_sc_hd__buf_2 _14670_ (.A(net7843),
    .X(_07841_));
 sky130_fd_sc_hd__a211o_1 _14671_ (.A1(_07821_),
    .A2(_07830_),
    .B1(_07839_),
    .C1(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__buf_2 _14672_ (.A(net7850),
    .X(_07843_));
 sky130_fd_sc_hd__a21o_1 _14673_ (.A1(_07820_),
    .A2(_07842_),
    .B1(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__o21ai_1 _14674_ (.A1(_07818_),
    .A2(_07837_),
    .B1(net8491),
    .Y(_07845_));
 sky130_fd_sc_hd__nand2_1 _14675_ (.A(_07841_),
    .B(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__nand2_1 _14676_ (.A(_07843_),
    .B(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__a21o_1 _14677_ (.A1(_07844_),
    .A2(_07847_),
    .B1(net8354),
    .X(_07848_));
 sky130_fd_sc_hd__xnor2_2 _14678_ (.A(_07779_),
    .B(_07655_),
    .Y(_07849_));
 sky130_fd_sc_hd__xnor2_1 _14679_ (.A(_07780_),
    .B(_07783_),
    .Y(_07850_));
 sky130_fd_sc_hd__nor2_1 _14680_ (.A(net7795),
    .B(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__o21ba_1 _14681_ (.A1(_07818_),
    .A2(_07849_),
    .B1_N(_07851_),
    .X(_07852_));
 sky130_fd_sc_hd__xnor2_1 _14682_ (.A(_07510_),
    .B(_07787_),
    .Y(_07853_));
 sky130_fd_sc_hd__xnor2_1 _14683_ (.A(_07784_),
    .B(_07786_),
    .Y(_07854_));
 sky130_fd_sc_hd__nor2_1 _14684_ (.A(net8442),
    .B(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__a21oi_1 _14685_ (.A1(_07818_),
    .A2(_07853_),
    .B1(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__and2_1 _14686_ (.A(net7811),
    .B(_07856_),
    .X(_07857_));
 sky130_fd_sc_hd__a21oi_1 _14687_ (.A1(_07841_),
    .A2(_07852_),
    .B1(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__clkbuf_1 _14688_ (.A(net7812),
    .X(_07859_));
 sky130_fd_sc_hd__clkbuf_4 _14689_ (.A(_07818_),
    .X(_07860_));
 sky130_fd_sc_hd__xor2_4 _14690_ (.A(_07776_),
    .B(_07778_),
    .X(_07861_));
 sky130_fd_sc_hd__nor2_1 _14691_ (.A(_07695_),
    .B(_07774_),
    .Y(_07862_));
 sky130_fd_sc_hd__xnor2_2 _14692_ (.A(_07732_),
    .B(_07862_),
    .Y(_07863_));
 sky130_fd_sc_hd__and2_1 _14693_ (.A(_07821_),
    .B(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__a21o_1 _14694_ (.A1(_07860_),
    .A2(_07861_),
    .B1(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__and3_1 _14695_ (.A(net7813),
    .B(net7811),
    .C(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__a211o_1 _14696_ (.A1(_07843_),
    .A2(_07858_),
    .B1(_07866_),
    .C1(net7839),
    .X(_07867_));
 sky130_fd_sc_hd__clkbuf_2 _14697_ (.A(net4703),
    .X(_07868_));
 sky130_fd_sc_hd__clkbuf_4 _14698_ (.A(net4704),
    .X(_07869_));
 sky130_fd_sc_hd__a31o_2 _14699_ (.A1(net7833),
    .A2(_07848_),
    .A3(_07867_),
    .B1(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__and4_1 _14700_ (.A(net3774),
    .B(_04485_),
    .C(_04479_),
    .D(_06117_),
    .X(_07871_));
 sky130_fd_sc_hd__buf_4 _14701_ (.A(net3775),
    .X(_07872_));
 sky130_fd_sc_hd__mux2_1 _14702_ (.A0(net4381),
    .A1(_07870_),
    .S(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__clkbuf_1 _14703_ (.A(_07873_),
    .X(_00391_));
 sky130_fd_sc_hd__xnor2_1 _14704_ (.A(_07828_),
    .B(_07816_),
    .Y(_07874_));
 sky130_fd_sc_hd__nor2_1 _14705_ (.A(_07818_),
    .B(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__a211o_1 _14706_ (.A1(_07860_),
    .A2(_07830_),
    .B1(_07875_),
    .C1(net7811),
    .X(_07876_));
 sky130_fd_sc_hd__nor2_2 _14707_ (.A(net7795),
    .B(_07837_),
    .Y(_07877_));
 sky130_fd_sc_hd__and3_4 _14708_ (.A(net7795),
    .B(_07837_),
    .C(_07838_),
    .X(_07878_));
 sky130_fd_sc_hd__or3_4 _14709_ (.A(net7843),
    .B(_07877_),
    .C(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__a31o_1 _14710_ (.A1(net7813),
    .A2(_07876_),
    .A3(_07879_),
    .B1(net8354),
    .X(_07880_));
 sky130_fd_sc_hd__nor2_1 _14711_ (.A(net7795),
    .B(_07854_),
    .Y(_07881_));
 sky130_fd_sc_hd__nor2_1 _14712_ (.A(net8442),
    .B(_07850_),
    .Y(_07882_));
 sky130_fd_sc_hd__or3_1 _14713_ (.A(net7811),
    .B(_07881_),
    .C(_07882_),
    .X(_07883_));
 sky130_fd_sc_hd__and2_1 _14714_ (.A(net7795),
    .B(_07853_),
    .X(_07884_));
 sky130_fd_sc_hd__a211o_1 _14715_ (.A1(_07860_),
    .A2(_07804_),
    .B1(_07884_),
    .C1(net7843),
    .X(_07885_));
 sky130_fd_sc_hd__nor2_1 _14716_ (.A(net8444),
    .B(_07849_),
    .Y(_07886_));
 sky130_fd_sc_hd__a21oi_1 _14717_ (.A1(_07821_),
    .A2(_07861_),
    .B1(_07886_),
    .Y(_07887_));
 sky130_fd_sc_hd__nand2_1 _14718_ (.A(_07818_),
    .B(_07863_),
    .Y(_07888_));
 sky130_fd_sc_hd__a21o_1 _14719_ (.A1(_07841_),
    .A2(_07888_),
    .B1(_07843_),
    .X(_07889_));
 sky130_fd_sc_hd__a21oi_1 _14720_ (.A1(net7811),
    .A2(_07887_),
    .B1(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__a311o_1 _14721_ (.A1(_07843_),
    .A2(_07883_),
    .A3(_07885_),
    .B1(_07890_),
    .C1(net7839),
    .X(_07891_));
 sky130_fd_sc_hd__a31o_2 _14722_ (.A1(net7833),
    .A2(_07880_),
    .A3(_07891_),
    .B1(_07869_),
    .X(_07892_));
 sky130_fd_sc_hd__mux2_1 _14723_ (.A0(net4351),
    .A1(_07892_),
    .S(_07872_),
    .X(_07893_));
 sky130_fd_sc_hd__clkbuf_1 _14724_ (.A(_07893_),
    .X(_00392_));
 sky130_fd_sc_hd__nand2_1 _14725_ (.A(_07841_),
    .B(_07856_),
    .Y(_07894_));
 sky130_fd_sc_hd__o21ai_1 _14726_ (.A1(_07841_),
    .A2(_07819_),
    .B1(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand2_1 _14727_ (.A(_07841_),
    .B(_07865_),
    .Y(_07896_));
 sky130_fd_sc_hd__o211a_1 _14728_ (.A1(_07841_),
    .A2(_07852_),
    .B1(_07896_),
    .C1(net7813),
    .X(_07897_));
 sky130_fd_sc_hd__a21oi_1 _14729_ (.A1(_07843_),
    .A2(_07895_),
    .B1(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__a211o_1 _14730_ (.A1(_07821_),
    .A2(_07830_),
    .B1(_07839_),
    .C1(net7811),
    .X(_07899_));
 sky130_fd_sc_hd__or2_1 _14731_ (.A(net7843),
    .B(_07845_),
    .X(_07900_));
 sky130_fd_sc_hd__a31o_1 _14732_ (.A1(net7813),
    .A2(_07899_),
    .A3(_07900_),
    .B1(net8354),
    .X(_07901_));
 sky130_fd_sc_hd__o211ai_1 _14733_ (.A1(net7839),
    .A2(_07898_),
    .B1(_07901_),
    .C1(net7833),
    .Y(_07902_));
 sky130_fd_sc_hd__or2b_2 _14734_ (.A(_07869_),
    .B_N(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__mux2_1 _14735_ (.A0(net4399),
    .A1(_07903_),
    .S(_07872_),
    .X(_07904_));
 sky130_fd_sc_hd__clkbuf_1 _14736_ (.A(_07904_),
    .X(_00393_));
 sky130_fd_sc_hd__a211o_1 _14737_ (.A1(_07860_),
    .A2(_07804_),
    .B1(_07884_),
    .C1(net7811),
    .X(_07905_));
 sky130_fd_sc_hd__a211o_1 _14738_ (.A1(_07860_),
    .A2(_07830_),
    .B1(_07875_),
    .C1(net7843),
    .X(_07906_));
 sky130_fd_sc_hd__nand2_1 _14739_ (.A(net7843),
    .B(_07887_),
    .Y(_07907_));
 sky130_fd_sc_hd__o311a_1 _14740_ (.A1(net7843),
    .A2(_07881_),
    .A3(_07882_),
    .B1(_07907_),
    .C1(net7812),
    .X(_07908_));
 sky130_fd_sc_hd__a311o_1 _14741_ (.A1(net7850),
    .A2(_07905_),
    .A3(_07906_),
    .B1(_07908_),
    .C1(net7839),
    .X(_07909_));
 sky130_fd_sc_hd__o211a_1 _14742_ (.A1(_07877_),
    .A2(_07878_),
    .B1(net7813),
    .C1(net7843),
    .X(_07910_));
 sky130_fd_sc_hd__o21a_1 _14743_ (.A1(net8354),
    .A2(_07910_),
    .B1(net7833),
    .X(_07911_));
 sky130_fd_sc_hd__clkbuf_1 _14744_ (.A(net7784),
    .X(_07912_));
 sky130_fd_sc_hd__clkbuf_4 _14745_ (.A(net7787),
    .X(_07913_));
 sky130_fd_sc_hd__a21bo_1 _14746_ (.A1(_07821_),
    .A2(_07861_),
    .B1_N(_07888_),
    .X(_07914_));
 sky130_fd_sc_hd__and3_1 _14747_ (.A(net7785),
    .B(_07913_),
    .C(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__clkbuf_1 _14748_ (.A(net7823),
    .X(_07916_));
 sky130_fd_sc_hd__a221o_2 _14749_ (.A1(_07909_),
    .A2(_07911_),
    .B1(_07915_),
    .B2(net7824),
    .C1(net7806),
    .X(_07917_));
 sky130_fd_sc_hd__mux2_1 _14750_ (.A0(net4539),
    .A1(_07917_),
    .S(_07872_),
    .X(_07918_));
 sky130_fd_sc_hd__clkbuf_1 _14751_ (.A(_07918_),
    .X(_00394_));
 sky130_fd_sc_hd__a211oi_1 _14752_ (.A1(_07841_),
    .A2(_07852_),
    .B1(_07857_),
    .C1(net7850),
    .Y(_07919_));
 sky130_fd_sc_hd__a31o_1 _14753_ (.A1(_07843_),
    .A2(_07820_),
    .A3(_07842_),
    .B1(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__nor2_1 _14754_ (.A(net7850),
    .B(_07846_),
    .Y(_07921_));
 sky130_fd_sc_hd__mux2_1 _14755_ (.A0(_07920_),
    .A1(_07921_),
    .S(net7839),
    .X(_07922_));
 sky130_fd_sc_hd__nor2_1 _14756_ (.A(net7843),
    .B(_07821_),
    .Y(_07923_));
 sky130_fd_sc_hd__nor2_1 _14757_ (.A(net7845),
    .B(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__nand2_1 _14758_ (.A(_07818_),
    .B(_07861_),
    .Y(_07925_));
 sky130_fd_sc_hd__o21ai_2 _14759_ (.A1(_07860_),
    .A2(_07849_),
    .B1(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__or2_1 _14760_ (.A(net7787),
    .B(_07864_),
    .X(_07927_));
 sky130_fd_sc_hd__o211a_1 _14761_ (.A1(net7846),
    .A2(_07926_),
    .B1(_07927_),
    .C1(net7785),
    .X(_07928_));
 sky130_fd_sc_hd__a221o_2 _14762_ (.A1(net7833),
    .A2(_07922_),
    .B1(_07928_),
    .B2(net7824),
    .C1(net4704),
    .X(_07929_));
 sky130_fd_sc_hd__mux2_1 _14763_ (.A0(net4403),
    .A1(_07929_),
    .S(_07872_),
    .X(_07930_));
 sky130_fd_sc_hd__clkbuf_1 _14764_ (.A(_07930_),
    .X(_00395_));
 sky130_fd_sc_hd__nor2_1 _14765_ (.A(_06505_),
    .B(net7839),
    .Y(_07931_));
 sky130_fd_sc_hd__and3_1 _14766_ (.A(net7813),
    .B(_07883_),
    .C(_07885_),
    .X(_07932_));
 sky130_fd_sc_hd__a31o_1 _14767_ (.A1(_07843_),
    .A2(_07876_),
    .A3(_07879_),
    .B1(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__clkbuf_4 _14768_ (.A(net7785),
    .X(_07934_));
 sky130_fd_sc_hd__or2_1 _14769_ (.A(_07882_),
    .B(_07886_),
    .X(_07935_));
 sky130_fd_sc_hd__mux2_1 _14770_ (.A0(_07914_),
    .A1(_07935_),
    .S(_07913_),
    .X(_07936_));
 sky130_fd_sc_hd__and2_2 _14771_ (.A(_07934_),
    .B(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__a221o_2 _14772_ (.A1(_07931_),
    .A2(_07933_),
    .B1(_07937_),
    .B2(net7824),
    .C1(net4704),
    .X(_07938_));
 sky130_fd_sc_hd__mux2_1 _14773_ (.A0(net4415),
    .A1(_07938_),
    .S(_07872_),
    .X(_07939_));
 sky130_fd_sc_hd__clkbuf_1 _14774_ (.A(_07939_),
    .X(_00396_));
 sky130_fd_sc_hd__a21o_1 _14775_ (.A1(_07899_),
    .A2(_07900_),
    .B1(net7813),
    .X(_07940_));
 sky130_fd_sc_hd__nand2_1 _14776_ (.A(net7833),
    .B(net8354),
    .Y(_07941_));
 sky130_fd_sc_hd__a21oi_1 _14777_ (.A1(net7813),
    .A2(_07895_),
    .B1(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__and3_1 _14778_ (.A(net7843),
    .B(_07821_),
    .C(_07863_),
    .X(_07943_));
 sky130_fd_sc_hd__or2_1 _14779_ (.A(_07851_),
    .B(_07855_),
    .X(_07944_));
 sky130_fd_sc_hd__mux2_1 _14780_ (.A0(_07926_),
    .A1(_07944_),
    .S(_07913_),
    .X(_07945_));
 sky130_fd_sc_hd__mux2_1 _14781_ (.A0(_07943_),
    .A1(_07945_),
    .S(_07934_),
    .X(_07946_));
 sky130_fd_sc_hd__a221o_2 _14782_ (.A1(_07940_),
    .A2(_07942_),
    .B1(_07946_),
    .B2(net7824),
    .C1(net4704),
    .X(_07947_));
 sky130_fd_sc_hd__mux2_1 _14783_ (.A0(net4379),
    .A1(_07947_),
    .S(_07872_),
    .X(_07948_));
 sky130_fd_sc_hd__clkbuf_1 _14784_ (.A(_07948_),
    .X(_00397_));
 sky130_fd_sc_hd__a21o_1 _14785_ (.A1(_07905_),
    .A2(_07906_),
    .B1(_07843_),
    .X(_07949_));
 sky130_fd_sc_hd__o21ai_1 _14786_ (.A1(_07877_),
    .A2(_07878_),
    .B1(_07841_),
    .Y(_07950_));
 sky130_fd_sc_hd__a21oi_1 _14787_ (.A1(_07843_),
    .A2(_07950_),
    .B1(_07941_),
    .Y(_07951_));
 sky130_fd_sc_hd__nor2_1 _14788_ (.A(_07881_),
    .B(_07884_),
    .Y(_07952_));
 sky130_fd_sc_hd__nand2_1 _14789_ (.A(net7846),
    .B(_07935_),
    .Y(_07953_));
 sky130_fd_sc_hd__o211a_1 _14790_ (.A1(net7846),
    .A2(_07952_),
    .B1(_07953_),
    .C1(net7785),
    .X(_07954_));
 sky130_fd_sc_hd__a21oi_1 _14791_ (.A1(_07913_),
    .A2(_07914_),
    .B1(_07934_),
    .Y(_07955_));
 sky130_fd_sc_hd__nor2_1 _14792_ (.A(_07954_),
    .B(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__a221o_1 _14793_ (.A1(_07949_),
    .A2(_07951_),
    .B1(_07956_),
    .B2(net7824),
    .C1(net4704),
    .X(_07957_));
 sky130_fd_sc_hd__mux2_1 _14794_ (.A0(net4392),
    .A1(net7825),
    .S(_07872_),
    .X(_07958_));
 sky130_fd_sc_hd__clkbuf_1 _14795_ (.A(_07958_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _14796_ (.A0(_07804_),
    .A1(_07853_),
    .S(_07818_),
    .X(_07959_));
 sky130_fd_sc_hd__mux4_1 _14797_ (.A0(_07864_),
    .A1(_07926_),
    .A2(_07944_),
    .A3(_07959_),
    .S0(net532),
    .S1(net7785),
    .X(_07960_));
 sky130_fd_sc_hd__a21o_1 _14798_ (.A1(net7824),
    .A2(_07960_),
    .B1(net7806),
    .X(_07961_));
 sky130_fd_sc_hd__a31o_2 _14799_ (.A1(_07844_),
    .A2(_07847_),
    .A3(_07931_),
    .B1(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__mux2_1 _14800_ (.A0(net4390),
    .A1(_07962_),
    .S(_07872_),
    .X(_07963_));
 sky130_fd_sc_hd__clkbuf_1 _14801_ (.A(_07963_),
    .X(_00399_));
 sky130_fd_sc_hd__and3_1 _14802_ (.A(net7813),
    .B(_07876_),
    .C(_07879_),
    .X(_07964_));
 sky130_fd_sc_hd__or2_1 _14803_ (.A(_07881_),
    .B(_07884_),
    .X(_07965_));
 sky130_fd_sc_hd__a21o_1 _14804_ (.A1(_07818_),
    .A2(_07804_),
    .B1(_07875_),
    .X(_07966_));
 sky130_fd_sc_hd__mux4_2 _14805_ (.A0(_07914_),
    .A1(_07935_),
    .A2(_07965_),
    .A3(_07966_),
    .S0(net531),
    .S1(net7785),
    .X(_07967_));
 sky130_fd_sc_hd__a221o_4 _14806_ (.A1(_07964_),
    .A2(_07931_),
    .B1(_07967_),
    .B2(net7823),
    .C1(net3638),
    .X(_07968_));
 sky130_fd_sc_hd__mux2_1 _14807_ (.A0(net4461),
    .A1(_07968_),
    .S(_07872_),
    .X(_07969_));
 sky130_fd_sc_hd__clkbuf_1 _14808_ (.A(_07969_),
    .X(_00400_));
 sky130_fd_sc_hd__and3_1 _14809_ (.A(net7813),
    .B(_07899_),
    .C(_07900_),
    .X(_07970_));
 sky130_fd_sc_hd__nor2_1 _14810_ (.A(_07821_),
    .B(_07874_),
    .Y(_07971_));
 sky130_fd_sc_hd__a21o_1 _14811_ (.A1(_07821_),
    .A2(_07830_),
    .B1(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__mux4_2 _14812_ (.A0(_07926_),
    .A1(_07944_),
    .A2(_07959_),
    .A3(_07972_),
    .S0(net7787),
    .S1(net7785),
    .X(_07973_));
 sky130_fd_sc_hd__a21o_1 _14813_ (.A1(net7793),
    .A2(_07943_),
    .B1(net3638),
    .X(_07974_));
 sky130_fd_sc_hd__a221o_4 _14814_ (.A1(net8354),
    .A2(_07970_),
    .B1(_07973_),
    .B2(net7824),
    .C1(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__buf_4 _14815_ (.A(net3775),
    .X(_07976_));
 sky130_fd_sc_hd__mux2_1 _14816_ (.A0(net3777),
    .A1(_07975_),
    .S(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__clkbuf_1 _14817_ (.A(_07977_),
    .X(_00401_));
 sky130_fd_sc_hd__a21o_1 _14818_ (.A1(_07860_),
    .A2(_07830_),
    .B1(_07878_),
    .X(_07978_));
 sky130_fd_sc_hd__mux4_2 _14819_ (.A0(_07935_),
    .A1(_07965_),
    .A2(_07966_),
    .A3(_07978_),
    .S0(_07913_),
    .S1(net7785),
    .X(_07979_));
 sky130_fd_sc_hd__a221o_1 _14820_ (.A1(net8354),
    .A2(_07910_),
    .B1(_07915_),
    .B2(net7793),
    .C1(net3638),
    .X(_07980_));
 sky130_fd_sc_hd__a21o_2 _14821_ (.A1(net7824),
    .A2(_07979_),
    .B1(_07980_),
    .X(_07981_));
 sky130_fd_sc_hd__mux2_1 _14822_ (.A0(net4496),
    .A1(_07981_),
    .S(_07976_),
    .X(_07982_));
 sky130_fd_sc_hd__clkbuf_1 _14823_ (.A(_07982_),
    .X(_00402_));
 sky130_fd_sc_hd__inv_2 _14824_ (.A(_07944_),
    .Y(_07983_));
 sky130_fd_sc_hd__inv_2 _14825_ (.A(_07959_),
    .Y(_07984_));
 sky130_fd_sc_hd__a21oi_1 _14826_ (.A1(_07821_),
    .A2(_07830_),
    .B1(_07971_),
    .Y(_07985_));
 sky130_fd_sc_hd__nor2_1 _14827_ (.A(_07860_),
    .B(_07837_),
    .Y(_07986_));
 sky130_fd_sc_hd__nor2_1 _14828_ (.A(_07839_),
    .B(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__mux4_2 _14829_ (.A0(_07983_),
    .A1(_07984_),
    .A2(_07985_),
    .A3(_07987_),
    .S0(_07913_),
    .S1(net7785),
    .X(_07988_));
 sky130_fd_sc_hd__clkbuf_2 _14830_ (.A(net7793),
    .X(_07989_));
 sky130_fd_sc_hd__a221o_1 _14831_ (.A1(net8354),
    .A2(_07921_),
    .B1(_07928_),
    .B2(net7794),
    .C1(net7806),
    .X(_07990_));
 sky130_fd_sc_hd__o21bai_4 _14832_ (.A1(net8362),
    .A2(_07988_),
    .B1_N(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__mux2_1 _14833_ (.A0(net4435),
    .A1(_07991_),
    .S(_07976_),
    .X(_07992_));
 sky130_fd_sc_hd__clkbuf_1 _14834_ (.A(_07992_),
    .X(_00403_));
 sky130_fd_sc_hd__a21oi_1 _14835_ (.A1(_07860_),
    .A2(_07804_),
    .B1(_07875_),
    .Y(_07993_));
 sky130_fd_sc_hd__a21oi_1 _14836_ (.A1(_07860_),
    .A2(_07830_),
    .B1(_07878_),
    .Y(_07994_));
 sky130_fd_sc_hd__inv_2 _14837_ (.A(_07877_),
    .Y(_07995_));
 sky130_fd_sc_hd__mux4_1 _14838_ (.A0(_07952_),
    .A1(_07993_),
    .A2(_07994_),
    .A3(_07995_),
    .S0(_07913_),
    .S1(net7785),
    .X(_07996_));
 sky130_fd_sc_hd__nor2_1 _14839_ (.A(net8362),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__a211o_2 _14840_ (.A1(net7794),
    .A2(_07937_),
    .B1(_07997_),
    .C1(net4704),
    .X(_07998_));
 sky130_fd_sc_hd__mux2_1 _14841_ (.A0(net4481),
    .A1(_07998_),
    .S(_07976_),
    .X(_07999_));
 sky130_fd_sc_hd__clkbuf_1 _14842_ (.A(_07999_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(_07959_),
    .A1(_07972_),
    .S(_07913_),
    .X(_08000_));
 sky130_fd_sc_hd__o21ai_2 _14844_ (.A1(_07839_),
    .A2(_07986_),
    .B1(net7846),
    .Y(_08001_));
 sky130_fd_sc_hd__nand2_1 _14845_ (.A(_07934_),
    .B(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__o211a_1 _14846_ (.A1(_07934_),
    .A2(_08000_),
    .B1(_08002_),
    .C1(net7824),
    .X(_08003_));
 sky130_fd_sc_hd__a211o_2 _14847_ (.A1(net7794),
    .A2(_07946_),
    .B1(_08003_),
    .C1(net4704),
    .X(_08004_));
 sky130_fd_sc_hd__mux2_1 _14848_ (.A0(net4430),
    .A1(_08004_),
    .S(_07976_),
    .X(_08005_));
 sky130_fd_sc_hd__clkbuf_1 _14849_ (.A(_08005_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _14850_ (.A0(_07966_),
    .A1(_07978_),
    .S(_07913_),
    .X(_08006_));
 sky130_fd_sc_hd__o21ai_1 _14851_ (.A1(net7811),
    .A2(_07995_),
    .B1(_07934_),
    .Y(_08007_));
 sky130_fd_sc_hd__o211ai_2 _14852_ (.A1(_07934_),
    .A2(_08006_),
    .B1(_08007_),
    .C1(net7824),
    .Y(_08008_));
 sky130_fd_sc_hd__a21oi_1 _14853_ (.A1(net7794),
    .A2(_07956_),
    .B1(net4704),
    .Y(_08009_));
 sky130_fd_sc_hd__nand2_2 _14854_ (.A(_08008_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(net4459),
    .A1(_08010_),
    .S(_07976_),
    .X(_08011_));
 sky130_fd_sc_hd__clkbuf_1 _14856_ (.A(_08011_),
    .X(_00406_));
 sky130_fd_sc_hd__nor2_1 _14857_ (.A(net7846),
    .B(_07987_),
    .Y(_08012_));
 sky130_fd_sc_hd__nor2_1 _14858_ (.A(_07913_),
    .B(_07985_),
    .Y(_08013_));
 sky130_fd_sc_hd__nand2_1 _14859_ (.A(net8491),
    .B(_07934_),
    .Y(_08014_));
 sky130_fd_sc_hd__o311a_1 _14860_ (.A1(_07934_),
    .A2(_08012_),
    .A3(_08013_),
    .B1(_08014_),
    .C1(_06543_),
    .X(_08015_));
 sky130_fd_sc_hd__a21o_1 _14861_ (.A1(_06545_),
    .A2(_07960_),
    .B1(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__a21o_2 _14862_ (.A1(_06505_),
    .A2(_08016_),
    .B1(_07869_),
    .X(_08017_));
 sky130_fd_sc_hd__mux2_1 _14863_ (.A0(net4440),
    .A1(_08017_),
    .S(_07976_),
    .X(_08018_));
 sky130_fd_sc_hd__clkbuf_1 _14864_ (.A(_08018_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _14865_ (.A0(_07877_),
    .A1(_07978_),
    .S(net7846),
    .X(_08019_));
 sky130_fd_sc_hd__nor2_2 _14866_ (.A(_07934_),
    .B(net8362),
    .Y(_08020_));
 sky130_fd_sc_hd__a221o_2 _14867_ (.A1(net7794),
    .A2(_07967_),
    .B1(_08019_),
    .B2(_08020_),
    .C1(_07869_),
    .X(_08021_));
 sky130_fd_sc_hd__mux2_1 _14868_ (.A0(net4428),
    .A1(_08021_),
    .S(_07976_),
    .X(_08022_));
 sky130_fd_sc_hd__clkbuf_1 _14869_ (.A(_08022_),
    .X(_00408_));
 sky130_fd_sc_hd__inv_2 _14870_ (.A(_08001_),
    .Y(_08023_));
 sky130_fd_sc_hd__a221oi_4 _14871_ (.A1(net7794),
    .A2(_07973_),
    .B1(_08023_),
    .B2(_08020_),
    .C1(_07869_),
    .Y(_08024_));
 sky130_fd_sc_hd__inv_2 _14872_ (.A(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__mux2_1 _14873_ (.A0(net4537),
    .A1(_08025_),
    .S(_07976_),
    .X(_08026_));
 sky130_fd_sc_hd__clkbuf_1 _14874_ (.A(_08026_),
    .X(_00409_));
 sky130_fd_sc_hd__nor2_1 _14875_ (.A(net7811),
    .B(_07995_),
    .Y(_08027_));
 sky130_fd_sc_hd__a221o_1 _14876_ (.A1(net7794),
    .A2(_07979_),
    .B1(_08027_),
    .B2(_08020_),
    .C1(_07869_),
    .X(_08028_));
 sky130_fd_sc_hd__mux2_1 _14877_ (.A0(net4524),
    .A1(_08028_),
    .S(_07976_),
    .X(_08029_));
 sky130_fd_sc_hd__clkbuf_1 _14878_ (.A(_08029_),
    .X(_00410_));
 sky130_fd_sc_hd__o21bai_2 _14879_ (.A1(net8370),
    .A2(_07988_),
    .B1_N(_07869_),
    .Y(_08030_));
 sky130_fd_sc_hd__mux2_1 _14880_ (.A0(net4608),
    .A1(_08030_),
    .S(net3775),
    .X(_08031_));
 sky130_fd_sc_hd__clkbuf_1 _14881_ (.A(_08031_),
    .X(_00411_));
 sky130_fd_sc_hd__nor3_1 _14882_ (.A(_07869_),
    .B(net8370),
    .C(_07996_),
    .Y(_08032_));
 sky130_fd_sc_hd__mux2_1 _14883_ (.A0(net4413),
    .A1(_08032_),
    .S(net3775),
    .X(_08033_));
 sky130_fd_sc_hd__clkbuf_1 _14884_ (.A(_08033_),
    .X(_00412_));
 sky130_fd_sc_hd__clkbuf_4 _14885_ (.A(_06239_),
    .X(_08034_));
 sky130_fd_sc_hd__o21ai_2 _14886_ (.A1(_06163_),
    .A2(_06235_),
    .B1(_06237_),
    .Y(_08035_));
 sky130_fd_sc_hd__clkbuf_4 _14887_ (.A(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__clkbuf_4 _14888_ (.A(_06237_),
    .X(_08037_));
 sky130_fd_sc_hd__clkbuf_8 _14889_ (.A(_04481_),
    .X(_08038_));
 sky130_fd_sc_hd__o21a_1 _14890_ (.A1(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A2(_08037_),
    .B1(_08038_),
    .X(_08039_));
 sky130_fd_sc_hd__o221a_1 _14891_ (.A1(net4667),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net3749),
    .C1(net4543),
    .X(_00413_));
 sky130_fd_sc_hd__o21a_1 _14892_ (.A1(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A2(_08037_),
    .B1(_08038_),
    .X(_08040_));
 sky130_fd_sc_hd__o221a_1 _14893_ (.A1(net4506),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net4518),
    .C1(net4679),
    .X(_00414_));
 sky130_fd_sc_hd__o21a_1 _14894_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08037_),
    .B1(_08038_),
    .X(_08041_));
 sky130_fd_sc_hd__o221a_1 _14895_ (.A1(net3945),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net3932),
    .C1(net4671),
    .X(_00415_));
 sky130_fd_sc_hd__o21a_1 _14896_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(_08037_),
    .B1(_08038_),
    .X(_08042_));
 sky130_fd_sc_hd__o221a_1 _14897_ (.A1(net4569),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net3787),
    .C1(net4744),
    .X(_00416_));
 sky130_fd_sc_hd__clkbuf_4 _14898_ (.A(_04481_),
    .X(_08043_));
 sky130_fd_sc_hd__o21a_1 _14899_ (.A1(net4277),
    .A2(_08037_),
    .B1(_08043_),
    .X(_08044_));
 sky130_fd_sc_hd__o221a_1 _14900_ (.A1(net4541),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net4565),
    .C1(net4571),
    .X(_00417_));
 sky130_fd_sc_hd__o21a_1 _14901_ (.A1(net4268),
    .A2(_08037_),
    .B1(_08043_),
    .X(_08045_));
 sky130_fd_sc_hd__o221a_1 _14902_ (.A1(net4547),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net3847),
    .C1(net8238),
    .X(_00418_));
 sky130_fd_sc_hd__o21a_1 _14903_ (.A1(net4236),
    .A2(_08037_),
    .B1(_08043_),
    .X(_08046_));
 sky130_fd_sc_hd__o221a_1 _14904_ (.A1(net4508),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net3757),
    .C1(net8240),
    .X(_00419_));
 sky130_fd_sc_hd__clkbuf_4 _14905_ (.A(_06237_),
    .X(_08047_));
 sky130_fd_sc_hd__o21a_1 _14906_ (.A1(net4280),
    .A2(_08047_),
    .B1(_08043_),
    .X(_08048_));
 sky130_fd_sc_hd__o221a_1 _14907_ (.A1(net4500),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net3768),
    .C1(net4683),
    .X(_00420_));
 sky130_fd_sc_hd__o21a_1 _14908_ (.A1(net4293),
    .A2(_08047_),
    .B1(_08043_),
    .X(_08049_));
 sky130_fd_sc_hd__o221a_1 _14909_ (.A1(net3888),
    .A2(_08034_),
    .B1(_08036_),
    .B2(net3785),
    .C1(net4730),
    .X(_00421_));
 sky130_fd_sc_hd__clkbuf_4 _14910_ (.A(_06239_),
    .X(_08050_));
 sky130_fd_sc_hd__o21a_1 _14911_ (.A1(net8018),
    .A2(_08047_),
    .B1(_08043_),
    .X(_08051_));
 sky130_fd_sc_hd__o221a_1 _14912_ (.A1(net4665),
    .A2(_08050_),
    .B1(_08036_),
    .B2(net4567),
    .C1(net4551),
    .X(_00422_));
 sky130_fd_sc_hd__clkbuf_4 _14913_ (.A(_08035_),
    .X(_08052_));
 sky130_fd_sc_hd__o21a_1 _14914_ (.A1(net8021),
    .A2(_08047_),
    .B1(_08043_),
    .X(_08053_));
 sky130_fd_sc_hd__o221a_1 _14915_ (.A1(net3796),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net3790),
    .C1(net4577),
    .X(_00423_));
 sky130_fd_sc_hd__o21a_1 _14916_ (.A1(net8029),
    .A2(_08047_),
    .B1(_08043_),
    .X(_08054_));
 sky130_fd_sc_hd__o221a_1 _14917_ (.A1(net4669),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net4526),
    .C1(net4585),
    .X(_00424_));
 sky130_fd_sc_hd__o21a_1 _14918_ (.A1(net4917),
    .A2(_08047_),
    .B1(_08043_),
    .X(_08055_));
 sky130_fd_sc_hd__o221a_1 _14919_ (.A1(net4589),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net3751),
    .C1(net4695),
    .X(_00425_));
 sky130_fd_sc_hd__o21a_1 _14920_ (.A1(net8071),
    .A2(_08047_),
    .B1(_08043_),
    .X(_08056_));
 sky130_fd_sc_hd__o221a_1 _14921_ (.A1(net4657),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net3766),
    .C1(net4691),
    .X(_00426_));
 sky130_fd_sc_hd__o21a_1 _14922_ (.A1(net8012),
    .A2(_08047_),
    .B1(_04482_),
    .X(_08057_));
 sky130_fd_sc_hd__o221a_1 _14923_ (.A1(net4610),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net3811),
    .C1(net4738),
    .X(_00427_));
 sky130_fd_sc_hd__o21a_1 _14924_ (.A1(net8009),
    .A2(_08047_),
    .B1(_04482_),
    .X(_08058_));
 sky130_fd_sc_hd__o221a_1 _14925_ (.A1(net4651),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net3669),
    .C1(net4758),
    .X(_00428_));
 sky130_fd_sc_hd__o21a_1 _14926_ (.A1(net8270),
    .A2(_08047_),
    .B1(_04482_),
    .X(_08059_));
 sky130_fd_sc_hd__o221a_1 _14927_ (.A1(net4659),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net3803),
    .C1(net4752),
    .X(_00429_));
 sky130_fd_sc_hd__o21a_1 _14928_ (.A1(net8264),
    .A2(_06237_),
    .B1(_04482_),
    .X(_08060_));
 sky130_fd_sc_hd__o221a_1 _14929_ (.A1(net3875),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net4575),
    .C1(net4719),
    .X(_00430_));
 sky130_fd_sc_hd__o21a_1 _14930_ (.A1(net8467),
    .A2(_06237_),
    .B1(_04482_),
    .X(_08061_));
 sky130_fd_sc_hd__o221a_1 _14931_ (.A1(net3913),
    .A2(_08050_),
    .B1(_08052_),
    .B2(net3820),
    .C1(net4706),
    .X(_00431_));
 sky130_fd_sc_hd__o21a_1 _14932_ (.A1(net8088),
    .A2(_06237_),
    .B1(_04482_),
    .X(_08062_));
 sky130_fd_sc_hd__o221a_1 _14933_ (.A1(net4655),
    .A2(_06239_),
    .B1(_08052_),
    .B2(net3835),
    .C1(net4675),
    .X(_00432_));
 sky130_fd_sc_hd__o21a_1 _14934_ (.A1(net7821),
    .A2(_06237_),
    .B1(_04482_),
    .X(_08063_));
 sky130_fd_sc_hd__o221a_1 _14935_ (.A1(net3943),
    .A2(_06239_),
    .B1(_08035_),
    .B2(net3926),
    .C1(net4661),
    .X(_00433_));
 sky130_fd_sc_hd__o21ai_1 _14936_ (.A1(net3933),
    .A2(_06235_),
    .B1(net1791),
    .Y(_08064_));
 sky130_fd_sc_hd__clkbuf_4 _14937_ (.A(_04481_),
    .X(_01633_));
 sky130_fd_sc_hd__o21ai_1 _14938_ (.A1(net8034),
    .A2(_08037_),
    .B1(_01633_),
    .Y(_08065_));
 sky130_fd_sc_hd__a21oi_1 _14939_ (.A1(_08037_),
    .A2(net1792),
    .B1(net4332),
    .Y(_00434_));
 sky130_fd_sc_hd__or4_1 _14940_ (.A(net3871),
    .B(net3976),
    .C(net3774),
    .D(_04485_),
    .X(_08066_));
 sky130_fd_sc_hd__nor2_2 _14941_ (.A(_04489_),
    .B(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__buf_4 _14942_ (.A(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__mux2_1 _14943_ (.A0(net3822),
    .A1(_07870_),
    .S(_08068_),
    .X(_08069_));
 sky130_fd_sc_hd__clkbuf_1 _14944_ (.A(_08069_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _14945_ (.A0(net4535),
    .A1(_07892_),
    .S(_08068_),
    .X(_08070_));
 sky130_fd_sc_hd__clkbuf_1 _14946_ (.A(_08070_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _14947_ (.A0(net4353),
    .A1(_07903_),
    .S(_08068_),
    .X(_08071_));
 sky130_fd_sc_hd__clkbuf_1 _14948_ (.A(_08071_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _14949_ (.A0(net4485),
    .A1(_07917_),
    .S(_08068_),
    .X(_08072_));
 sky130_fd_sc_hd__clkbuf_1 _14950_ (.A(_08072_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(net4630),
    .A1(_07929_),
    .S(_08068_),
    .X(_08073_));
 sky130_fd_sc_hd__clkbuf_1 _14952_ (.A(_08073_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _14953_ (.A0(net4583),
    .A1(_07938_),
    .S(_08068_),
    .X(_08074_));
 sky130_fd_sc_hd__clkbuf_1 _14954_ (.A(_08074_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _14955_ (.A0(net4383),
    .A1(_07947_),
    .S(_08068_),
    .X(_08075_));
 sky130_fd_sc_hd__clkbuf_1 _14956_ (.A(_08075_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(net4789),
    .A1(net7825),
    .S(_08068_),
    .X(_08076_));
 sky130_fd_sc_hd__clkbuf_1 _14958_ (.A(_08076_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _14959_ (.A0(net4776),
    .A1(_07962_),
    .S(_08068_),
    .X(_08077_));
 sky130_fd_sc_hd__clkbuf_1 _14960_ (.A(_08077_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _14961_ (.A0(net4471),
    .A1(_07968_),
    .S(_08068_),
    .X(_08078_));
 sky130_fd_sc_hd__clkbuf_1 _14962_ (.A(_08078_),
    .X(_00444_));
 sky130_fd_sc_hd__buf_4 _14963_ (.A(_08067_),
    .X(_08079_));
 sky130_fd_sc_hd__mux2_1 _14964_ (.A0(net4397),
    .A1(_07975_),
    .S(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__clkbuf_1 _14965_ (.A(_08080_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _14966_ (.A0(net4373),
    .A1(_07981_),
    .S(_08079_),
    .X(_08081_));
 sky130_fd_sc_hd__clkbuf_1 _14967_ (.A(_08081_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _14968_ (.A0(net4483),
    .A1(_07991_),
    .S(_08079_),
    .X(_08082_));
 sky130_fd_sc_hd__clkbuf_1 _14969_ (.A(_08082_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _14970_ (.A0(net4401),
    .A1(_07998_),
    .S(_08079_),
    .X(_08083_));
 sky130_fd_sc_hd__clkbuf_1 _14971_ (.A(_08083_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _14972_ (.A0(net4405),
    .A1(_08004_),
    .S(_08079_),
    .X(_08084_));
 sky130_fd_sc_hd__clkbuf_1 _14973_ (.A(_08084_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14974_ (.A0(net4522),
    .A1(_08010_),
    .S(_08079_),
    .X(_08085_));
 sky130_fd_sc_hd__clkbuf_1 _14975_ (.A(_08085_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _14976_ (.A0(net4653),
    .A1(_08017_),
    .S(_08079_),
    .X(_08086_));
 sky130_fd_sc_hd__clkbuf_1 _14977_ (.A(_08086_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _14978_ (.A0(net4624),
    .A1(_08021_),
    .S(_08079_),
    .X(_08087_));
 sky130_fd_sc_hd__clkbuf_1 _14979_ (.A(_08087_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _14980_ (.A0(net4520),
    .A1(_08025_),
    .S(_08079_),
    .X(_08088_));
 sky130_fd_sc_hd__clkbuf_1 _14981_ (.A(_08088_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _14982_ (.A0(net4756),
    .A1(_08028_),
    .S(_08079_),
    .X(_08089_));
 sky130_fd_sc_hd__clkbuf_1 _14983_ (.A(_08089_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _14984_ (.A0(net4388),
    .A1(_08030_),
    .S(_08067_),
    .X(_08090_));
 sky130_fd_sc_hd__clkbuf_1 _14985_ (.A(_08090_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _14986_ (.A0(net4622),
    .A1(_08032_),
    .S(_08067_),
    .X(_08091_));
 sky130_fd_sc_hd__clkbuf_1 _14987_ (.A(_08091_),
    .X(_00456_));
 sky130_fd_sc_hd__buf_4 _14988_ (.A(net92),
    .X(_08092_));
 sky130_fd_sc_hd__buf_4 _14989_ (.A(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__and2_1 _14990_ (.A(_08093_),
    .B(net4156),
    .X(_08094_));
 sky130_fd_sc_hd__clkbuf_1 _14991_ (.A(net4157),
    .X(_00457_));
 sky130_fd_sc_hd__nor2_1 _14992_ (.A(net63),
    .B(net7571),
    .Y(_00458_));
 sky130_fd_sc_hd__and2_1 _14993_ (.A(_08093_),
    .B(net4149),
    .X(_08095_));
 sky130_fd_sc_hd__clkbuf_1 _14994_ (.A(net4150),
    .X(_00459_));
 sky130_fd_sc_hd__and2_1 _14995_ (.A(_08093_),
    .B(net4141),
    .X(_08096_));
 sky130_fd_sc_hd__clkbuf_1 _14996_ (.A(net4142),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _14997_ (.A(_08093_),
    .B(net4164),
    .X(_08097_));
 sky130_fd_sc_hd__clkbuf_1 _14998_ (.A(net4165),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _14999_ (.A(_08093_),
    .B(net7727),
    .X(_08098_));
 sky130_fd_sc_hd__clkbuf_1 _15000_ (.A(net4174),
    .X(_00462_));
 sky130_fd_sc_hd__or2_1 _15001_ (.A(_06102_),
    .B(_06158_),
    .X(_08099_));
 sky130_fd_sc_hd__a2bb2o_1 _15002_ (.A1_N(_06145_),
    .A2_N(_08099_),
    .B1(net1013),
    .B2(_06102_),
    .X(_08100_));
 sky130_fd_sc_hd__mux2_1 _15003_ (.A0(net740),
    .A1(_08100_),
    .S(net3985),
    .X(_08101_));
 sky130_fd_sc_hd__inv_2 _15004_ (.A(_06115_),
    .Y(_08102_));
 sky130_fd_sc_hd__buf_6 _15005_ (.A(net4865),
    .X(_08103_));
 sky130_fd_sc_hd__a21oi_1 _15006_ (.A1(_08102_),
    .A2(_06159_),
    .B1(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__mux2_1 _15007_ (.A0(_04567_),
    .A1(net3986),
    .S(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__and2_1 _15008_ (.A(_08038_),
    .B(net3987),
    .X(_08106_));
 sky130_fd_sc_hd__clkbuf_1 _15009_ (.A(net3988),
    .X(_00463_));
 sky130_fd_sc_hd__a2bb2o_1 _15010_ (.A1_N(net4009),
    .A2_N(_08099_),
    .B1(net951),
    .B2(_06102_),
    .X(_08107_));
 sky130_fd_sc_hd__mux2_1 _15011_ (.A0(net1004),
    .A1(net4010),
    .S(net3985),
    .X(_08108_));
 sky130_fd_sc_hd__mux2_1 _15012_ (.A0(_04566_),
    .A1(net4011),
    .S(_08104_),
    .X(_08109_));
 sky130_fd_sc_hd__and2_1 _15013_ (.A(_08038_),
    .B(net4012),
    .X(_08110_));
 sky130_fd_sc_hd__clkbuf_1 _15014_ (.A(net4013),
    .X(_00464_));
 sky130_fd_sc_hd__buf_4 _15015_ (.A(net4182),
    .X(_08111_));
 sky130_fd_sc_hd__o211a_1 _15016_ (.A1(net4183),
    .A2(_08037_),
    .B1(_08034_),
    .C1(_01633_),
    .X(_00465_));
 sky130_fd_sc_hd__nor2_1 _15017_ (.A(_04476_),
    .B(net3452),
    .Y(_08112_));
 sky130_fd_sc_hd__buf_4 _15018_ (.A(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__buf_4 _15019_ (.A(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__buf_4 _15020_ (.A(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__or2b_1 _15021_ (.A(net3628),
    .B_N(_06117_),
    .X(_08116_));
 sky130_fd_sc_hd__buf_4 _15022_ (.A(_08116_),
    .X(_08117_));
 sky130_fd_sc_hd__buf_4 _15023_ (.A(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__buf_4 _15024_ (.A(_08118_),
    .X(_08119_));
 sky130_fd_sc_hd__mux2_1 _15025_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(net4181),
    .X(_08120_));
 sky130_fd_sc_hd__mux2_2 _15026_ (.A0(_07892_),
    .A1(net8403),
    .S(_08114_),
    .X(_08121_));
 sky130_fd_sc_hd__and3_1 _15027_ (.A(net4083),
    .B(net3627),
    .C(_06117_),
    .X(_08122_));
 sky130_fd_sc_hd__buf_4 _15028_ (.A(_08122_),
    .X(_08123_));
 sky130_fd_sc_hd__buf_4 _15029_ (.A(_08123_),
    .X(_08124_));
 sky130_fd_sc_hd__a21o_1 _15030_ (.A1(net4351),
    .A2(_08124_),
    .B1(_06119_),
    .X(_08125_));
 sky130_fd_sc_hd__a21oi_2 _15031_ (.A1(_08119_),
    .A2(_08121_),
    .B1(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__clkbuf_4 _15032_ (.A(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__buf_4 _15033_ (.A(_06121_),
    .X(_08128_));
 sky130_fd_sc_hd__clkbuf_8 _15034_ (.A(_08119_),
    .X(_08129_));
 sky130_fd_sc_hd__nand2_1 _15035_ (.A(net4917),
    .B(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__or2_2 _15036_ (.A(_08128_),
    .B(net4918),
    .X(_08131_));
 sky130_fd_sc_hd__nor2_1 _15037_ (.A(_08127_),
    .B(_08131_),
    .Y(_08132_));
 sky130_fd_sc_hd__buf_4 _15038_ (.A(_08124_),
    .X(_08133_));
 sky130_fd_sc_hd__mux2_1 _15039_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(net4181),
    .X(_08134_));
 sky130_fd_sc_hd__mux2_2 _15040_ (.A0(_07870_),
    .A1(net8365),
    .S(_08114_),
    .X(_08135_));
 sky130_fd_sc_hd__or3b_4 _15041_ (.A(net3774),
    .B(_04485_),
    .C_N(_06117_),
    .X(_08136_));
 sky130_fd_sc_hd__buf_4 _15042_ (.A(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__o21a_1 _15043_ (.A1(net4381),
    .A2(_08119_),
    .B1(_08137_),
    .X(_08138_));
 sky130_fd_sc_hd__o21ai_4 _15044_ (.A1(_08133_),
    .A2(_08135_),
    .B1(_08138_),
    .Y(_08139_));
 sky130_fd_sc_hd__nand2_2 _15045_ (.A(net8261),
    .B(_08119_),
    .Y(_08140_));
 sky130_fd_sc_hd__or2_1 _15046_ (.A(_06120_),
    .B(net8072),
    .X(_08141_));
 sky130_fd_sc_hd__clkbuf_4 _15047_ (.A(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__nor2_1 _15048_ (.A(_08139_),
    .B(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand2_1 _15049_ (.A(_08132_),
    .B(_08143_),
    .Y(_08144_));
 sky130_fd_sc_hd__xnor2_2 _15050_ (.A(net3489),
    .B(net3417),
    .Y(_08145_));
 sky130_fd_sc_hd__nand2_1 _15051_ (.A(_06033_),
    .B(_08145_),
    .Y(_08146_));
 sky130_fd_sc_hd__o211a_1 _15052_ (.A1(net3489),
    .A2(_06033_),
    .B1(_08123_),
    .C1(_08146_),
    .X(_08147_));
 sky130_fd_sc_hd__clkbuf_4 _15053_ (.A(_06118_),
    .X(_08148_));
 sky130_fd_sc_hd__a21o_1 _15054_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(_08117_),
    .B1(_08148_),
    .X(_08149_));
 sky130_fd_sc_hd__and2_1 _15055_ (.A(_06374_),
    .B(_06375_),
    .X(_08150_));
 sky130_fd_sc_hd__or4_1 _15056_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .C(_06349_),
    .D(_06340_),
    .X(_08151_));
 sky130_fd_sc_hd__or4_1 _15057_ (.A(_06334_),
    .B(_06331_),
    .C(_06324_),
    .D(net8409),
    .X(_08152_));
 sky130_fd_sc_hd__or4_1 _15058_ (.A(_06364_),
    .B(_06321_),
    .C(_06317_),
    .D(net8410),
    .X(_08153_));
 sky130_fd_sc_hd__nor3_1 _15059_ (.A(_06361_),
    .B(_06314_),
    .C(net8411),
    .Y(_08154_));
 sky130_fd_sc_hd__inv_2 _15060_ (.A(_06416_),
    .Y(_08155_));
 sky130_fd_sc_hd__a31o_4 _15061_ (.A1(_06370_),
    .A2(_08150_),
    .A3(net8412),
    .B1(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__nand2_1 _15062_ (.A(net3536),
    .B(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__xnor2_2 _15063_ (.A(net3536),
    .B(net4168),
    .Y(_08158_));
 sky130_fd_sc_hd__o21a_1 _15064_ (.A1(_08156_),
    .A2(_08158_),
    .B1(_08148_),
    .X(_08159_));
 sky130_fd_sc_hd__a2bb2o_2 _15065_ (.A1_N(_08147_),
    .A2_N(net7835),
    .B1(_08157_),
    .B2(_08159_),
    .X(_08160_));
 sky130_fd_sc_hd__buf_2 _15066_ (.A(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__buf_4 _15067_ (.A(_08137_),
    .X(_08162_));
 sky130_fd_sc_hd__mux2_1 _15068_ (.A0(_05997_),
    .A1(_06317_),
    .S(net4180),
    .X(_08163_));
 sky130_fd_sc_hd__mux2_2 _15069_ (.A0(_07962_),
    .A1(net8372),
    .S(_08113_),
    .X(_08164_));
 sky130_fd_sc_hd__a21o_2 _15070_ (.A1(net4390),
    .A2(_08123_),
    .B1(_08148_),
    .X(_08165_));
 sky130_fd_sc_hd__a21o_1 _15071_ (.A1(_08118_),
    .A2(_08164_),
    .B1(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__buf_4 _15072_ (.A(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__o21ai_4 _15073_ (.A1(net4776),
    .A2(_08162_),
    .B1(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__or3_1 _15074_ (.A(net3348),
    .B(net3536),
    .C(net4168),
    .X(_08169_));
 sky130_fd_sc_hd__o21ai_1 _15075_ (.A1(net3536),
    .A2(net4168),
    .B1(net3348),
    .Y(_08170_));
 sky130_fd_sc_hd__nand2_1 _15076_ (.A(_08169_),
    .B(_08170_),
    .Y(_08171_));
 sky130_fd_sc_hd__o21a_1 _15077_ (.A1(_08156_),
    .A2(_08171_),
    .B1(_08148_),
    .X(_08172_));
 sky130_fd_sc_hd__nand2_1 _15078_ (.A(net7765),
    .B(net8413),
    .Y(_08173_));
 sky130_fd_sc_hd__a21o_1 _15079_ (.A1(net4277),
    .A2(_08117_),
    .B1(_08148_),
    .X(_08174_));
 sky130_fd_sc_hd__or3_2 _15080_ (.A(net5859),
    .B(net3489),
    .C(net3417),
    .X(_08175_));
 sky130_fd_sc_hd__o21ai_1 _15081_ (.A1(net3489),
    .A2(net3417),
    .B1(net5859),
    .Y(_08176_));
 sky130_fd_sc_hd__nand2_2 _15082_ (.A(_08175_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__nand2_1 _15083_ (.A(_06033_),
    .B(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__o211a_1 _15084_ (.A1(net3315),
    .A2(_06033_),
    .B1(_08123_),
    .C1(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__o2bb2a_4 _15085_ (.A1_N(_08172_),
    .A2_N(_08173_),
    .B1(net8422),
    .B2(_08179_),
    .X(_08180_));
 sky130_fd_sc_hd__clkbuf_8 _15086_ (.A(_08162_),
    .X(_08181_));
 sky130_fd_sc_hd__mux2_1 _15087_ (.A0(net8377),
    .A1(_06321_),
    .S(net4181),
    .X(_08182_));
 sky130_fd_sc_hd__mux2_1 _15088_ (.A0(_07957_),
    .A1(net8378),
    .S(_08113_),
    .X(_08183_));
 sky130_fd_sc_hd__a21o_1 _15089_ (.A1(net4392),
    .A2(_08123_),
    .B1(_08148_),
    .X(_08184_));
 sky130_fd_sc_hd__a21o_4 _15090_ (.A1(_08118_),
    .A2(_08183_),
    .B1(_08184_),
    .X(_08185_));
 sky130_fd_sc_hd__o21a_1 _15091_ (.A1(net3637),
    .A2(_08181_),
    .B1(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__a2bb2o_1 _15092_ (.A1_N(_08161_),
    .A2_N(_08168_),
    .B1(_08180_),
    .B2(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__or2_1 _15093_ (.A(net3372),
    .B(_08175_),
    .X(_08188_));
 sky130_fd_sc_hd__nand2_1 _15094_ (.A(net3372),
    .B(_08175_),
    .Y(_08189_));
 sky130_fd_sc_hd__and2_1 _15095_ (.A(_08188_),
    .B(_08189_),
    .X(_08190_));
 sky130_fd_sc_hd__or2_1 _15096_ (.A(net3372),
    .B(_06033_),
    .X(_08191_));
 sky130_fd_sc_hd__o211a_1 _15097_ (.A1(net7776),
    .A2(_08190_),
    .B1(_08191_),
    .C1(_08124_),
    .X(_08192_));
 sky130_fd_sc_hd__a21o_1 _15098_ (.A1(net4268),
    .A2(_08118_),
    .B1(_06119_),
    .X(_08193_));
 sky130_fd_sc_hd__buf_4 _15099_ (.A(_08156_),
    .X(_08194_));
 sky130_fd_sc_hd__nand2_1 _15100_ (.A(net5887),
    .B(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__or2_2 _15101_ (.A(net5887),
    .B(_08169_),
    .X(_08196_));
 sky130_fd_sc_hd__nand2_1 _15102_ (.A(net5887),
    .B(_08169_),
    .Y(_08197_));
 sky130_fd_sc_hd__nand2_2 _15103_ (.A(_08196_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__o21a_1 _15104_ (.A1(_08194_),
    .A2(_08198_),
    .B1(_06120_),
    .X(_08199_));
 sky130_fd_sc_hd__a2bb2o_4 _15105_ (.A1_N(_08192_),
    .A2_N(net8425),
    .B1(_08195_),
    .B2(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__mux2_1 _15106_ (.A0(_06002_),
    .A1(_06324_),
    .S(net4180),
    .X(_08201_));
 sky130_fd_sc_hd__mux2_1 _15107_ (.A0(_07947_),
    .A1(net8397),
    .S(_08113_),
    .X(_08202_));
 sky130_fd_sc_hd__a21o_1 _15108_ (.A1(net4379),
    .A2(_08123_),
    .B1(_08148_),
    .X(_08203_));
 sky130_fd_sc_hd__a21o_4 _15109_ (.A1(_08118_),
    .A2(_08202_),
    .B1(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__or2_2 _15110_ (.A(net3459),
    .B(_08136_),
    .X(_08205_));
 sky130_fd_sc_hd__nand2_1 _15111_ (.A(_08204_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__buf_2 _15112_ (.A(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__nor2_1 _15113_ (.A(_08200_),
    .B(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__a2bb2o_1 _15114_ (.A1_N(_08179_),
    .A2_N(_08174_),
    .B1(_08173_),
    .B2(_08172_),
    .X(_08209_));
 sky130_fd_sc_hd__o21ai_1 _15115_ (.A1(net3637),
    .A2(_08162_),
    .B1(_08185_),
    .Y(_08210_));
 sky130_fd_sc_hd__clkbuf_4 _15116_ (.A(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__or4_1 _15117_ (.A(_08160_),
    .B(_08168_),
    .C(net8414),
    .D(_08211_),
    .X(_08212_));
 sky130_fd_sc_hd__a21bo_2 _15118_ (.A1(_08187_),
    .A2(_08208_),
    .B1_N(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__xor2_1 _15119_ (.A(net4344),
    .B(_08188_),
    .X(_08214_));
 sky130_fd_sc_hd__mux2_1 _15120_ (.A0(_08214_),
    .A1(net4344),
    .S(_06027_),
    .X(_08215_));
 sky130_fd_sc_hd__mux2_1 _15121_ (.A0(net4236),
    .A1(_08215_),
    .S(_08123_),
    .X(_08216_));
 sky130_fd_sc_hd__nand2_1 _15122_ (.A(net3419),
    .B(_08156_),
    .Y(_08217_));
 sky130_fd_sc_hd__xnor2_2 _15123_ (.A(net3419),
    .B(_08196_),
    .Y(_08218_));
 sky130_fd_sc_hd__o21a_1 _15124_ (.A1(_08156_),
    .A2(_08218_),
    .B1(_08148_),
    .X(_08219_));
 sky130_fd_sc_hd__a2bb2o_2 _15125_ (.A1_N(_06119_),
    .A2_N(_08216_),
    .B1(_08217_),
    .B2(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__buf_2 _15126_ (.A(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__mux2_1 _15127_ (.A0(_06006_),
    .A1(_06331_),
    .S(net4180),
    .X(_08222_));
 sky130_fd_sc_hd__mux2_2 _15128_ (.A0(_07938_),
    .A1(net8393),
    .S(_08113_),
    .X(_08223_));
 sky130_fd_sc_hd__a21o_1 _15129_ (.A1(net4415),
    .A2(_08123_),
    .B1(_08148_),
    .X(_08224_));
 sky130_fd_sc_hd__a21oi_1 _15130_ (.A1(_08118_),
    .A2(_08223_),
    .B1(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__buf_4 _15131_ (.A(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__nor2_1 _15132_ (.A(net4583),
    .B(_08137_),
    .Y(_08227_));
 sky130_fd_sc_hd__or2_1 _15133_ (.A(_08226_),
    .B(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__buf_2 _15134_ (.A(_08228_),
    .X(_08229_));
 sky130_fd_sc_hd__or3_1 _15135_ (.A(net3317),
    .B(net4344),
    .C(_08188_),
    .X(_08230_));
 sky130_fd_sc_hd__o21ai_1 _15136_ (.A1(net4344),
    .A2(_08188_),
    .B1(net3317),
    .Y(_08231_));
 sky130_fd_sc_hd__and2_1 _15137_ (.A(_08230_),
    .B(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__mux2_1 _15138_ (.A0(_08232_),
    .A1(net3317),
    .S(_06027_),
    .X(_08233_));
 sky130_fd_sc_hd__mux2_1 _15139_ (.A0(net4280),
    .A1(_08233_),
    .S(_08122_),
    .X(_08234_));
 sky130_fd_sc_hd__nand2_1 _15140_ (.A(net3339),
    .B(net8413),
    .Y(_08235_));
 sky130_fd_sc_hd__or3_1 _15141_ (.A(net5768),
    .B(net3419),
    .C(_08196_),
    .X(_08236_));
 sky130_fd_sc_hd__o21ai_1 _15142_ (.A1(net3419),
    .A2(_08196_),
    .B1(net3339),
    .Y(_08237_));
 sky130_fd_sc_hd__nand2_1 _15143_ (.A(_08236_),
    .B(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__o21a_1 _15144_ (.A1(_08156_),
    .A2(_08238_),
    .B1(_06118_),
    .X(_08239_));
 sky130_fd_sc_hd__a2bb2o_2 _15145_ (.A1_N(_08148_),
    .A2_N(_08234_),
    .B1(_08235_),
    .B2(_08239_),
    .X(_08240_));
 sky130_fd_sc_hd__buf_2 _15146_ (.A(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__or4_1 _15147_ (.A(_08206_),
    .B(_08221_),
    .C(_08229_),
    .D(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__and2_1 _15148_ (.A(_08204_),
    .B(_08205_),
    .X(_08243_));
 sky130_fd_sc_hd__inv_2 _15149_ (.A(_08220_),
    .Y(_08244_));
 sky130_fd_sc_hd__nor2_2 _15150_ (.A(_08226_),
    .B(_08227_),
    .Y(_08245_));
 sky130_fd_sc_hd__inv_2 _15151_ (.A(_08240_),
    .Y(_08246_));
 sky130_fd_sc_hd__a22o_1 _15152_ (.A1(_08243_),
    .A2(_08244_),
    .B1(_08245_),
    .B2(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__nand2_2 _15153_ (.A(_08242_),
    .B(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__mux2_1 _15154_ (.A0(_06007_),
    .A1(_06334_),
    .S(_04510_),
    .X(_08249_));
 sky130_fd_sc_hd__mux2_1 _15155_ (.A0(_07929_),
    .A1(net8418),
    .S(_08113_),
    .X(_08250_));
 sky130_fd_sc_hd__a21o_1 _15156_ (.A1(net4403),
    .A2(_08124_),
    .B1(_06119_),
    .X(_08251_));
 sky130_fd_sc_hd__a21o_2 _15157_ (.A1(_08118_),
    .A2(_08250_),
    .B1(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__clkbuf_4 _15158_ (.A(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__or2_2 _15159_ (.A(net4630),
    .B(_08137_),
    .X(_08254_));
 sky130_fd_sc_hd__nand2_2 _15160_ (.A(_08253_),
    .B(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__or2_2 _15161_ (.A(net3433),
    .B(_08230_),
    .X(_08256_));
 sky130_fd_sc_hd__nand2_1 _15162_ (.A(net3433),
    .B(_08230_),
    .Y(_08257_));
 sky130_fd_sc_hd__and2_1 _15163_ (.A(_08256_),
    .B(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__mux2_1 _15164_ (.A0(_08258_),
    .A1(net3433),
    .S(net7776),
    .X(_08259_));
 sky130_fd_sc_hd__mux2_1 _15165_ (.A0(net4293),
    .A1(_08259_),
    .S(_08124_),
    .X(_08260_));
 sky130_fd_sc_hd__or2_1 _15166_ (.A(net3457),
    .B(_08236_),
    .X(_08261_));
 sky130_fd_sc_hd__nand2_1 _15167_ (.A(net3457),
    .B(_08236_),
    .Y(_08262_));
 sky130_fd_sc_hd__nand2_1 _15168_ (.A(_08261_),
    .B(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__nor2_1 _15169_ (.A(_08156_),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__a211o_1 _15170_ (.A1(net3457),
    .A2(_08194_),
    .B1(_08264_),
    .C1(_08137_),
    .X(_08265_));
 sky130_fd_sc_hd__o21ai_4 _15171_ (.A1(_06120_),
    .A2(_08260_),
    .B1(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__nor2_2 _15172_ (.A(_08255_),
    .B(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__xnor2_4 _15173_ (.A(_08248_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__xnor2_4 _15174_ (.A(_08213_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__nand2_1 _15175_ (.A(_08244_),
    .B(_08245_),
    .Y(_08270_));
 sky130_fd_sc_hd__nor2_1 _15176_ (.A(net4630),
    .B(_08137_),
    .Y(_08271_));
 sky130_fd_sc_hd__or3b_2 _15177_ (.A(_08271_),
    .B(_08241_),
    .C_N(_08252_),
    .X(_08272_));
 sky130_fd_sc_hd__xnor2_2 _15178_ (.A(_08270_),
    .B(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__mux2_1 _15179_ (.A0(_06009_),
    .A1(_06340_),
    .S(net4180),
    .X(_08274_));
 sky130_fd_sc_hd__mux2_1 _15180_ (.A0(_07917_),
    .A1(net8055),
    .S(_08112_),
    .X(_08275_));
 sky130_fd_sc_hd__a21o_1 _15181_ (.A1(net4539),
    .A2(_08123_),
    .B1(_06118_),
    .X(_08276_));
 sky130_fd_sc_hd__a21oi_4 _15182_ (.A1(_08117_),
    .A2(_08275_),
    .B1(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__nor2_1 _15183_ (.A(net4485),
    .B(_08136_),
    .Y(_08278_));
 sky130_fd_sc_hd__or2_2 _15184_ (.A(_08277_),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__clkbuf_4 _15185_ (.A(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__or2_2 _15186_ (.A(_08266_),
    .B(_08280_),
    .X(_08281_));
 sky130_fd_sc_hd__or2_1 _15187_ (.A(_08270_),
    .B(_08272_),
    .X(_08282_));
 sky130_fd_sc_hd__o21ai_4 _15188_ (.A1(_08273_),
    .A2(_08281_),
    .B1(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__or2b_1 _15189_ (.A(_08269_),
    .B_N(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__a21bo_2 _15190_ (.A1(_08213_),
    .A2(_08268_),
    .B1_N(_08284_),
    .X(_08285_));
 sky130_fd_sc_hd__or2_1 _15191_ (.A(_08132_),
    .B(_08143_),
    .X(_08286_));
 sky130_fd_sc_hd__and2_2 _15192_ (.A(_08144_),
    .B(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__xor2_2 _15193_ (.A(net3445),
    .B(_08256_),
    .X(_08288_));
 sky130_fd_sc_hd__mux2_2 _15194_ (.A0(_08288_),
    .A1(net3445),
    .S(_06027_),
    .X(_08289_));
 sky130_fd_sc_hd__nand2_1 _15195_ (.A(_08133_),
    .B(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__a21oi_1 _15196_ (.A1(net8263),
    .A2(_08119_),
    .B1(_06120_),
    .Y(_08291_));
 sky130_fd_sc_hd__xnor2_1 _15197_ (.A(net3461),
    .B(_08261_),
    .Y(_08292_));
 sky130_fd_sc_hd__mux2_2 _15198_ (.A0(_08292_),
    .A1(_04695_),
    .S(_08194_),
    .X(_08293_));
 sky130_fd_sc_hd__a22o_4 _15199_ (.A1(_08290_),
    .A2(_08291_),
    .B1(_08293_),
    .B2(_06121_),
    .X(_08294_));
 sky130_fd_sc_hd__or3_4 _15200_ (.A(net2898),
    .B(net3461),
    .C(_08261_),
    .X(_08295_));
 sky130_fd_sc_hd__o21ai_1 _15201_ (.A1(net3461),
    .A2(_08261_),
    .B1(net2898),
    .Y(_08296_));
 sky130_fd_sc_hd__and2_1 _15202_ (.A(_08295_),
    .B(_08296_),
    .X(_08297_));
 sky130_fd_sc_hd__mux2_2 _15203_ (.A0(_08297_),
    .A1(net2898),
    .S(_08194_),
    .X(_08298_));
 sky130_fd_sc_hd__or3_4 _15204_ (.A(net4284),
    .B(net3445),
    .C(_08256_),
    .X(_08299_));
 sky130_fd_sc_hd__o21ai_1 _15205_ (.A1(net3445),
    .A2(_08256_),
    .B1(net4284),
    .Y(_08300_));
 sky130_fd_sc_hd__and2_1 _15206_ (.A(_08299_),
    .B(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__mux2_2 _15207_ (.A0(_08301_),
    .A1(net4188),
    .S(_06027_),
    .X(_08302_));
 sky130_fd_sc_hd__a21o_1 _15208_ (.A1(net8021),
    .A2(_08119_),
    .B1(_06120_),
    .X(_08303_));
 sky130_fd_sc_hd__a21o_1 _15209_ (.A1(_08133_),
    .A2(_08302_),
    .B1(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__o21ai_2 _15210_ (.A1(_08181_),
    .A2(_08298_),
    .B1(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__buf_2 _15211_ (.A(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__or4_1 _15212_ (.A(_08255_),
    .B(_08280_),
    .C(_08294_),
    .D(_08306_),
    .X(_08307_));
 sky130_fd_sc_hd__clkbuf_4 _15213_ (.A(_08294_),
    .X(_08308_));
 sky130_fd_sc_hd__buf_4 _15214_ (.A(_08306_),
    .X(_08309_));
 sky130_fd_sc_hd__o22ai_1 _15215_ (.A1(_08255_),
    .A2(_08308_),
    .B1(_08309_),
    .B2(_08280_),
    .Y(_08310_));
 sky130_fd_sc_hd__nand2_2 _15216_ (.A(_08307_),
    .B(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__a31o_1 _15217_ (.A1(net5902),
    .A2(_06502_),
    .A3(_07902_),
    .B1(_08113_),
    .X(_08312_));
 sky130_fd_sc_hd__mux2_1 _15218_ (.A0(_06010_),
    .A1(_06349_),
    .S(_04510_),
    .X(_08313_));
 sky130_fd_sc_hd__nand2_1 _15219_ (.A(_08114_),
    .B(net8044),
    .Y(_08314_));
 sky130_fd_sc_hd__a21o_1 _15220_ (.A1(_08312_),
    .A2(net8045),
    .B1(_08124_),
    .X(_08315_));
 sky130_fd_sc_hd__a21oi_1 _15221_ (.A1(net4399),
    .A2(_08124_),
    .B1(_06119_),
    .Y(_08316_));
 sky130_fd_sc_hd__a2bb2o_2 _15222_ (.A1_N(net4353),
    .A2_N(_08162_),
    .B1(_08315_),
    .B2(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__clkbuf_4 _15223_ (.A(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__nand2_1 _15224_ (.A(net8269),
    .B(_08129_),
    .Y(_08319_));
 sky130_fd_sc_hd__o31a_1 _15225_ (.A1(net7776),
    .A2(_08129_),
    .A3(_08299_),
    .B1(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__or3_1 _15226_ (.A(_08162_),
    .B(_08194_),
    .C(_08295_),
    .X(_08321_));
 sky130_fd_sc_hd__o21a_2 _15227_ (.A1(_08128_),
    .A2(_08320_),
    .B1(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__buf_2 _15228_ (.A(_08322_),
    .X(_08323_));
 sky130_fd_sc_hd__or2_2 _15229_ (.A(_08318_),
    .B(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__xnor2_4 _15230_ (.A(_08311_),
    .B(_08324_),
    .Y(_08325_));
 sky130_fd_sc_hd__buf_4 _15231_ (.A(_08308_),
    .X(_08326_));
 sky130_fd_sc_hd__or2_1 _15232_ (.A(_08305_),
    .B(_08318_),
    .X(_08327_));
 sky130_fd_sc_hd__o21bai_4 _15233_ (.A1(net4535),
    .A2(_08162_),
    .B1_N(_08126_),
    .Y(_08328_));
 sky130_fd_sc_hd__clkbuf_4 _15234_ (.A(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__nor2_1 _15235_ (.A(_08322_),
    .B(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__nor2_1 _15236_ (.A(_08280_),
    .B(_08294_),
    .Y(_08331_));
 sky130_fd_sc_hd__xnor2_1 _15237_ (.A(_08331_),
    .B(_08327_),
    .Y(_08332_));
 sky130_fd_sc_hd__nand2_1 _15238_ (.A(_08330_),
    .B(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__o31a_2 _15239_ (.A1(_08280_),
    .A2(_08326_),
    .A3(_08327_),
    .B1(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__xor2_4 _15240_ (.A(_08325_),
    .B(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__xor2_4 _15241_ (.A(_08287_),
    .B(_08335_),
    .X(_08336_));
 sky130_fd_sc_hd__xnor2_4 _15242_ (.A(_08285_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__buf_4 _15243_ (.A(_08131_),
    .X(_08338_));
 sky130_fd_sc_hd__nor2_2 _15244_ (.A(_08338_),
    .B(_08139_),
    .Y(_08339_));
 sky130_fd_sc_hd__xnor2_1 _15245_ (.A(_08330_),
    .B(_08332_),
    .Y(_08340_));
 sky130_fd_sc_hd__a21boi_4 _15246_ (.A1(net3822),
    .A2(_08128_),
    .B1_N(_08139_),
    .Y(_08341_));
 sky130_fd_sc_hd__nor2_1 _15247_ (.A(_08322_),
    .B(_08341_),
    .Y(_08342_));
 sky130_fd_sc_hd__or2_1 _15248_ (.A(_08294_),
    .B(_08317_),
    .X(_08343_));
 sky130_fd_sc_hd__nor2_1 _15249_ (.A(_08306_),
    .B(_08328_),
    .Y(_08344_));
 sky130_fd_sc_hd__xnor2_2 _15250_ (.A(_08343_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__or3_1 _15251_ (.A(_08306_),
    .B(_08328_),
    .C(_08343_),
    .X(_08346_));
 sky130_fd_sc_hd__a21boi_1 _15252_ (.A1(_08342_),
    .A2(_08345_),
    .B1_N(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__nand2_1 _15253_ (.A(_08340_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nor2_1 _15254_ (.A(_08340_),
    .B(_08347_),
    .Y(_08349_));
 sky130_fd_sc_hd__a21o_2 _15255_ (.A1(_08339_),
    .A2(_08348_),
    .B1(_08349_),
    .X(_08350_));
 sky130_fd_sc_hd__and2b_1 _15256_ (.A_N(_08337_),
    .B(_08350_),
    .X(_08351_));
 sky130_fd_sc_hd__a21oi_1 _15257_ (.A1(_08285_),
    .A2(_08336_),
    .B1(_08351_),
    .Y(_08352_));
 sky130_fd_sc_hd__or2_1 _15258_ (.A(_08144_),
    .B(_08352_),
    .X(_08353_));
 sky130_fd_sc_hd__inv_2 _15259_ (.A(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__or4_1 _15260_ (.A(_08168_),
    .B(_08211_),
    .C(_08221_),
    .D(_08241_),
    .X(_08355_));
 sky130_fd_sc_hd__a2bb2o_1 _15261_ (.A1_N(_08168_),
    .A2_N(_08221_),
    .B1(_08246_),
    .B2(_08186_),
    .X(_08356_));
 sky130_fd_sc_hd__nand2_1 _15262_ (.A(_08355_),
    .B(_08356_),
    .Y(_08357_));
 sky130_fd_sc_hd__or3_1 _15263_ (.A(_08207_),
    .B(_08266_),
    .C(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__nand2_1 _15264_ (.A(_08355_),
    .B(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__o21ai_1 _15265_ (.A1(_07968_),
    .A2(_07975_),
    .B1(_07981_),
    .Y(_08360_));
 sky130_fd_sc_hd__or3_1 _15266_ (.A(_07968_),
    .B(_07975_),
    .C(_07981_),
    .X(_08361_));
 sky130_fd_sc_hd__a21o_1 _15267_ (.A1(_08360_),
    .A2(_08361_),
    .B1(_08114_),
    .X(_08362_));
 sky130_fd_sc_hd__nand2_1 _15268_ (.A(net4181),
    .B(_06361_),
    .Y(_08363_));
 sky130_fd_sc_hd__o211a_1 _15269_ (.A1(_04511_),
    .A2(_06020_),
    .B1(_08114_),
    .C1(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__nor2_1 _15270_ (.A(_08124_),
    .B(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__a22o_4 _15271_ (.A1(net4496),
    .A2(_08133_),
    .B1(_08362_),
    .B2(_08365_),
    .X(_08366_));
 sky130_fd_sc_hd__nand2_1 _15272_ (.A(net4373),
    .B(_06120_),
    .Y(_08367_));
 sky130_fd_sc_hd__a21boi_1 _15273_ (.A1(_08181_),
    .A2(_08366_),
    .B1_N(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__xor2_1 _15274_ (.A(_07968_),
    .B(_07975_),
    .X(_08369_));
 sky130_fd_sc_hd__mux2_1 _15275_ (.A0(net8497),
    .A1(_06364_),
    .S(net4181),
    .X(_08370_));
 sky130_fd_sc_hd__nand2_1 _15276_ (.A(_08113_),
    .B(net8498),
    .Y(_08371_));
 sky130_fd_sc_hd__o211a_2 _15277_ (.A1(_08113_),
    .A2(_08369_),
    .B1(_08371_),
    .C1(_08118_),
    .X(_08372_));
 sky130_fd_sc_hd__o21ai_2 _15278_ (.A1(net3777),
    .A2(_08118_),
    .B1(_08137_),
    .Y(_08373_));
 sky130_fd_sc_hd__or2_4 _15279_ (.A(_08372_),
    .B(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__nand2_1 _15280_ (.A(net4397),
    .B(_06120_),
    .Y(_08375_));
 sky130_fd_sc_hd__and2_1 _15281_ (.A(_08374_),
    .B(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__or4_2 _15282_ (.A(_08161_),
    .B(net8414),
    .C(_08368_),
    .D(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__or2_1 _15283_ (.A(_04476_),
    .B(net3452),
    .X(_08378_));
 sky130_fd_sc_hd__nand2_1 _15284_ (.A(net4181),
    .B(_06314_),
    .Y(_08379_));
 sky130_fd_sc_hd__o21a_1 _15285_ (.A1(_04510_),
    .A2(_06025_),
    .B1(_08112_),
    .X(_08380_));
 sky130_fd_sc_hd__a22o_2 _15286_ (.A1(_07968_),
    .A2(net3453),
    .B1(_08379_),
    .B2(_08380_),
    .X(_08381_));
 sky130_fd_sc_hd__o21ai_2 _15287_ (.A1(net4461),
    .A2(_08117_),
    .B1(_08136_),
    .Y(_08382_));
 sky130_fd_sc_hd__a21o_4 _15288_ (.A1(_08119_),
    .A2(_08381_),
    .B1(_08382_),
    .X(_08383_));
 sky130_fd_sc_hd__a21boi_4 _15289_ (.A1(net4471),
    .A2(_06121_),
    .B1_N(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__or2_1 _15290_ (.A(_08200_),
    .B(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__nand2_1 _15291_ (.A(_08374_),
    .B(_08375_),
    .Y(_08386_));
 sky130_fd_sc_hd__a2bb2o_1 _15292_ (.A1_N(_08161_),
    .A2_N(_08368_),
    .B1(_08386_),
    .B2(_08180_),
    .X(_08387_));
 sky130_fd_sc_hd__nand3b_1 _15293_ (.A_N(_08385_),
    .B(_08387_),
    .C(_08377_),
    .Y(_08388_));
 sky130_fd_sc_hd__buf_2 _15294_ (.A(_08168_),
    .X(_08389_));
 sky130_fd_sc_hd__or4_1 _15295_ (.A(_08389_),
    .B(_08221_),
    .C(_08241_),
    .D(_08384_),
    .X(_08390_));
 sky130_fd_sc_hd__clkbuf_4 _15296_ (.A(_08241_),
    .X(_08391_));
 sky130_fd_sc_hd__buf_2 _15297_ (.A(_08384_),
    .X(_08392_));
 sky130_fd_sc_hd__o22ai_1 _15298_ (.A1(_08389_),
    .A2(_08391_),
    .B1(_08392_),
    .B2(_08221_),
    .Y(_08393_));
 sky130_fd_sc_hd__nand2_1 _15299_ (.A(_08390_),
    .B(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__nor2_1 _15300_ (.A(_08211_),
    .B(_08266_),
    .Y(_08395_));
 sky130_fd_sc_hd__xor2_1 _15301_ (.A(_08394_),
    .B(_08395_),
    .X(_08396_));
 sky130_fd_sc_hd__a21o_1 _15302_ (.A1(_08377_),
    .A2(_08388_),
    .B1(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__nand3_1 _15303_ (.A(_08377_),
    .B(_08388_),
    .C(_08396_),
    .Y(_08398_));
 sky130_fd_sc_hd__nand2_1 _15304_ (.A(_08397_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__xnor2_2 _15305_ (.A(_08359_),
    .B(_08399_),
    .Y(_08400_));
 sky130_fd_sc_hd__buf_2 _15306_ (.A(_08161_),
    .X(_08401_));
 sky130_fd_sc_hd__clkbuf_4 _15307_ (.A(net8414),
    .X(_08402_));
 sky130_fd_sc_hd__clkbuf_4 _15308_ (.A(_08368_),
    .X(_08403_));
 sky130_fd_sc_hd__o21a_4 _15309_ (.A1(_07968_),
    .A2(_07975_),
    .B1(_07981_),
    .X(_08404_));
 sky130_fd_sc_hd__xnor2_2 _15310_ (.A(_07991_),
    .B(_08404_),
    .Y(_08405_));
 sky130_fd_sc_hd__nand2_1 _15311_ (.A(_04511_),
    .B(_08150_),
    .Y(_08406_));
 sky130_fd_sc_hd__o211a_1 _15312_ (.A1(_04511_),
    .A2(net8500),
    .B1(_08114_),
    .C1(_08406_),
    .X(_08407_));
 sky130_fd_sc_hd__a211o_2 _15313_ (.A1(net3453),
    .A2(_08405_),
    .B1(_08407_),
    .C1(_08133_),
    .X(_08408_));
 sky130_fd_sc_hd__o21a_1 _15314_ (.A1(net3532),
    .A2(_08119_),
    .B1(_08162_),
    .X(_08409_));
 sky130_fd_sc_hd__a22oi_2 _15315_ (.A1(net3600),
    .A2(_06121_),
    .B1(_08408_),
    .B2(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__clkbuf_4 _15316_ (.A(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__or4_1 _15317_ (.A(_08401_),
    .B(_08402_),
    .C(_08403_),
    .D(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__nand2_2 _15318_ (.A(_08181_),
    .B(_08366_),
    .Y(_08413_));
 sky130_fd_sc_hd__nand2_2 _15319_ (.A(_08413_),
    .B(_08367_),
    .Y(_08414_));
 sky130_fd_sc_hd__a2bb2o_1 _15320_ (.A1_N(_08401_),
    .A2_N(_08411_),
    .B1(_08180_),
    .B2(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__nand2_1 _15321_ (.A(_08412_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__clkbuf_4 _15322_ (.A(_08200_),
    .X(_08417_));
 sky130_fd_sc_hd__buf_2 _15323_ (.A(_08376_),
    .X(_08418_));
 sky130_fd_sc_hd__nor2_1 _15324_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__xnor2_2 _15325_ (.A(_08416_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__buf_4 _15326_ (.A(net3453),
    .X(_08421_));
 sky130_fd_sc_hd__a211oi_4 _15327_ (.A1(_07989_),
    .A2(_07937_),
    .B1(_07997_),
    .C1(_07868_),
    .Y(_08422_));
 sky130_fd_sc_hd__nor2_2 _15328_ (.A(_07991_),
    .B(_08404_),
    .Y(_08423_));
 sky130_fd_sc_hd__xnor2_4 _15329_ (.A(_08422_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__nand2_1 _15330_ (.A(_04511_),
    .B(_06370_),
    .Y(_08425_));
 sky130_fd_sc_hd__o211a_2 _15331_ (.A1(_04511_),
    .A2(_05989_),
    .B1(_08114_),
    .C1(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__a211o_2 _15332_ (.A1(_08421_),
    .A2(_08424_),
    .B1(_08426_),
    .C1(_08133_),
    .X(_08427_));
 sky130_fd_sc_hd__o21a_2 _15333_ (.A1(net3599),
    .A2(_08119_),
    .B1(_08137_),
    .X(_08428_));
 sky130_fd_sc_hd__and2_1 _15334_ (.A(net4401),
    .B(_06121_),
    .X(_08429_));
 sky130_fd_sc_hd__a21o_2 _15335_ (.A1(_08427_),
    .A2(_08428_),
    .B1(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__mux2_1 _15336_ (.A0(net3417),
    .A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .S(_08117_),
    .X(_08431_));
 sky130_fd_sc_hd__or2_1 _15337_ (.A(_06119_),
    .B(net8399),
    .X(_08432_));
 sky130_fd_sc_hd__o21a_4 _15338_ (.A1(net4168),
    .A2(_08137_),
    .B1(net8400),
    .X(_08433_));
 sky130_fd_sc_hd__nand2_1 _15339_ (.A(_08430_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__inv_2 _15340_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .Y(_08435_));
 sky130_fd_sc_hd__o21ba_1 _15341_ (.A1(_06632_),
    .A2(_07988_),
    .B1_N(_07990_),
    .X(_08436_));
 sky130_fd_sc_hd__a211oi_1 _15342_ (.A1(_07989_),
    .A2(_07946_),
    .B1(_08003_),
    .C1(_07868_),
    .Y(_08437_));
 sky130_fd_sc_hd__a31o_1 _15343_ (.A1(_08436_),
    .A2(_08422_),
    .A3(_08360_),
    .B1(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__or4_4 _15344_ (.A(_07991_),
    .B(_07998_),
    .C(_08004_),
    .D(_08404_),
    .X(_08439_));
 sky130_fd_sc_hd__mux2_1 _15345_ (.A0(_05985_),
    .A1(_06416_),
    .S(net4180),
    .X(_08440_));
 sky130_fd_sc_hd__a21oi_4 _15346_ (.A1(_08113_),
    .A2(_08440_),
    .B1(_08123_),
    .Y(_08441_));
 sky130_fd_sc_hd__inv_2 _15347_ (.A(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a31o_4 _15348_ (.A1(net3453),
    .A2(_08438_),
    .A3(_08439_),
    .B1(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__or4_4 _15349_ (.A(net8065),
    .B(_06120_),
    .C(_08133_),
    .D(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__inv_2 _15350_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .Y(_08445_));
 sky130_fd_sc_hd__nor2_2 _15351_ (.A(net8041),
    .B(_08124_),
    .Y(_08446_));
 sky130_fd_sc_hd__and4_1 _15352_ (.A(_08436_),
    .B(_08422_),
    .C(_08437_),
    .D(_08360_),
    .X(_08447_));
 sky130_fd_sc_hd__o41a_1 _15353_ (.A1(_07991_),
    .A2(_07998_),
    .A3(_08004_),
    .A4(_08404_),
    .B1(_08010_),
    .X(_08448_));
 sky130_fd_sc_hd__a311o_1 _15354_ (.A1(_08008_),
    .A2(_08009_),
    .A3(_08447_),
    .B1(_08448_),
    .C1(_08114_),
    .X(_08449_));
 sky130_fd_sc_hd__a22o_4 _15355_ (.A1(net3574),
    .A2(_08133_),
    .B1(_08441_),
    .B2(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__and3_1 _15356_ (.A(_08181_),
    .B(_08446_),
    .C(_08450_),
    .X(_08451_));
 sky130_fd_sc_hd__xor2_2 _15357_ (.A(_08444_),
    .B(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__xor2_2 _15358_ (.A(_08434_),
    .B(_08452_),
    .X(_08453_));
 sky130_fd_sc_hd__inv_2 _15359_ (.A(_08428_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand2_1 _15360_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08117_),
    .Y(_08455_));
 sky130_fd_sc_hd__or4b_4 _15361_ (.A(_08454_),
    .B(_08444_),
    .C(net8033),
    .D_N(_08427_),
    .X(_08456_));
 sky130_fd_sc_hd__o21ai_2 _15362_ (.A1(net4168),
    .A2(_08162_),
    .B1(net8400),
    .Y(_08457_));
 sky130_fd_sc_hd__clkbuf_4 _15363_ (.A(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__nor2_1 _15364_ (.A(_08410_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__nand2_1 _15365_ (.A(net3531),
    .B(_08133_),
    .Y(_08460_));
 sky130_fd_sc_hd__a21o_1 _15366_ (.A1(_08460_),
    .A2(_08443_),
    .B1(_06121_),
    .X(_08461_));
 sky130_fd_sc_hd__nand2_1 _15367_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_08117_),
    .Y(_08462_));
 sky130_fd_sc_hd__nor2_1 _15368_ (.A(_06119_),
    .B(net4877),
    .Y(_08463_));
 sky130_fd_sc_hd__buf_2 _15369_ (.A(_08463_),
    .X(_08464_));
 sky130_fd_sc_hd__a21o_1 _15370_ (.A1(_08421_),
    .A2(_08424_),
    .B1(_08426_),
    .X(_08465_));
 sky130_fd_sc_hd__a2bb2o_1 _15371_ (.A1_N(_08461_),
    .A2_N(net8033),
    .B1(_08464_),
    .B2(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__nand3_2 _15372_ (.A(_08456_),
    .B(_08459_),
    .C(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__nand2_1 _15373_ (.A(_08456_),
    .B(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__xor2_2 _15374_ (.A(_08453_),
    .B(_08468_),
    .X(_08469_));
 sky130_fd_sc_hd__xnor2_2 _15375_ (.A(_08420_),
    .B(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__a21o_1 _15376_ (.A1(_08456_),
    .A2(_08466_),
    .B1(_08459_),
    .X(_08471_));
 sky130_fd_sc_hd__a21oi_4 _15377_ (.A1(net3453),
    .A2(_08405_),
    .B1(net8501),
    .Y(_08472_));
 sky130_fd_sc_hd__or2_1 _15378_ (.A(_06119_),
    .B(net4877),
    .X(_08473_));
 sky130_fd_sc_hd__clkbuf_4 _15379_ (.A(_08473_),
    .X(_08474_));
 sky130_fd_sc_hd__nor2_1 _15380_ (.A(_08472_),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__a31o_1 _15381_ (.A1(_08427_),
    .A2(_08428_),
    .A3(net8042),
    .B1(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__and4_1 _15382_ (.A(_08427_),
    .B(_08428_),
    .C(net8042),
    .D(_08475_),
    .X(_08477_));
 sky130_fd_sc_hd__a31o_1 _15383_ (.A1(_08414_),
    .A2(_08433_),
    .A3(_08476_),
    .B1(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__nand3_1 _15384_ (.A(_08467_),
    .B(_08471_),
    .C(_08478_),
    .Y(_08479_));
 sky130_fd_sc_hd__a21bo_1 _15385_ (.A1(_08377_),
    .A2(_08387_),
    .B1_N(_08385_),
    .X(_08480_));
 sky130_fd_sc_hd__and2_1 _15386_ (.A(_08388_),
    .B(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__a21o_1 _15387_ (.A1(_08467_),
    .A2(_08471_),
    .B1(_08478_),
    .X(_08482_));
 sky130_fd_sc_hd__and3_1 _15388_ (.A(_08479_),
    .B(_08481_),
    .C(_08482_),
    .X(_08483_));
 sky130_fd_sc_hd__a31o_1 _15389_ (.A1(_08467_),
    .A2(_08471_),
    .A3(_08478_),
    .B1(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__xnor2_2 _15390_ (.A(_08470_),
    .B(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__xnor2_2 _15391_ (.A(_08400_),
    .B(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__a21oi_1 _15392_ (.A1(_08479_),
    .A2(_08482_),
    .B1(_08481_),
    .Y(_08487_));
 sky130_fd_sc_hd__or4b_1 _15393_ (.A(_08403_),
    .B(_08458_),
    .C(_08477_),
    .D_N(_08476_),
    .X(_08488_));
 sky130_fd_sc_hd__nand4_1 _15394_ (.A(_08427_),
    .B(_08428_),
    .C(net8042),
    .D(_08475_),
    .Y(_08489_));
 sky130_fd_sc_hd__a22o_1 _15395_ (.A1(_08414_),
    .A2(_08433_),
    .B1(_08489_),
    .B2(_08476_),
    .X(_08490_));
 sky130_fd_sc_hd__buf_2 _15396_ (.A(_08133_),
    .X(_08491_));
 sky130_fd_sc_hd__or4b_2 _15397_ (.A(net8041),
    .B(_06120_),
    .C(_08491_),
    .D_N(_08408_),
    .X(_08492_));
 sky130_fd_sc_hd__or3b_1 _15398_ (.A(_06121_),
    .B(net4877),
    .C_N(_08366_),
    .X(_08493_));
 sky130_fd_sc_hd__nand2_4 _15399_ (.A(_08137_),
    .B(net8042),
    .Y(_08494_));
 sky130_fd_sc_hd__and4bb_1 _15400_ (.A_N(_08494_),
    .B_N(_08472_),
    .C(_08366_),
    .D(_08464_),
    .X(_08495_));
 sky130_fd_sc_hd__a21oi_4 _15401_ (.A1(_08492_),
    .A2(_08493_),
    .B1(_08495_),
    .Y(_08496_));
 sky130_fd_sc_hd__nor2_2 _15402_ (.A(_08418_),
    .B(_08458_),
    .Y(_08497_));
 sky130_fd_sc_hd__a21o_1 _15403_ (.A1(_08496_),
    .A2(_08497_),
    .B1(_08495_),
    .X(_08498_));
 sky130_fd_sc_hd__a21o_1 _15404_ (.A1(_08488_),
    .A2(_08490_),
    .B1(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__nor2_1 _15405_ (.A(net8414),
    .B(_08384_),
    .Y(_08500_));
 sky130_fd_sc_hd__nor2_1 _15406_ (.A(_08161_),
    .B(_08418_),
    .Y(_08501_));
 sky130_fd_sc_hd__xor2_1 _15407_ (.A(_08500_),
    .B(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__nor2_1 _15408_ (.A(_08389_),
    .B(_08417_),
    .Y(_08503_));
 sky130_fd_sc_hd__xor2_1 _15409_ (.A(_08502_),
    .B(_08503_),
    .X(_08504_));
 sky130_fd_sc_hd__nand3_1 _15410_ (.A(_08488_),
    .B(_08490_),
    .C(_08498_),
    .Y(_08505_));
 sky130_fd_sc_hd__a21boi_1 _15411_ (.A1(_08499_),
    .A2(_08504_),
    .B1_N(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__o21ai_2 _15412_ (.A1(_08483_),
    .A2(_08487_),
    .B1(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__a22o_1 _15413_ (.A1(_08186_),
    .A2(_08244_),
    .B1(_08246_),
    .B2(_08243_),
    .X(_08508_));
 sky130_fd_sc_hd__clkbuf_4 _15414_ (.A(_08266_),
    .X(_08509_));
 sky130_fd_sc_hd__nor2_1 _15415_ (.A(_08229_),
    .B(_08509_),
    .Y(_08510_));
 sky130_fd_sc_hd__or4_1 _15416_ (.A(_08211_),
    .B(_08207_),
    .C(_08221_),
    .D(_08241_),
    .X(_08511_));
 sky130_fd_sc_hd__a21bo_1 _15417_ (.A1(_08508_),
    .A2(_08510_),
    .B1_N(_08511_),
    .X(_08512_));
 sky130_fd_sc_hd__nand2_1 _15418_ (.A(_08500_),
    .B(_08501_),
    .Y(_08513_));
 sky130_fd_sc_hd__a21bo_1 _15419_ (.A1(_08502_),
    .A2(_08503_),
    .B1_N(_08513_),
    .X(_08514_));
 sky130_fd_sc_hd__o21ai_1 _15420_ (.A1(_08207_),
    .A2(_08509_),
    .B1(_08357_),
    .Y(_08515_));
 sky130_fd_sc_hd__nand2_1 _15421_ (.A(_08358_),
    .B(_08515_),
    .Y(_08516_));
 sky130_fd_sc_hd__xnor2_2 _15422_ (.A(_08514_),
    .B(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__xor2_2 _15423_ (.A(_08512_),
    .B(_08517_),
    .X(_08518_));
 sky130_fd_sc_hd__or3_4 _15424_ (.A(_08483_),
    .B(_08487_),
    .C(_08506_),
    .X(_08519_));
 sky130_fd_sc_hd__a21boi_2 _15425_ (.A1(_08507_),
    .A2(_08518_),
    .B1_N(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__xor2_1 _15426_ (.A(_08486_),
    .B(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__nor2_1 _15427_ (.A(_08229_),
    .B(_08294_),
    .Y(_08522_));
 sky130_fd_sc_hd__nor2_1 _15428_ (.A(_08255_),
    .B(_08306_),
    .Y(_08523_));
 sky130_fd_sc_hd__xnor2_1 _15429_ (.A(_08522_),
    .B(_08523_),
    .Y(_08524_));
 sky130_fd_sc_hd__or2_1 _15430_ (.A(_08280_),
    .B(_08323_),
    .X(_08525_));
 sky130_fd_sc_hd__xnor2_1 _15431_ (.A(_08524_),
    .B(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__o31a_1 _15432_ (.A1(_08311_),
    .A2(_08318_),
    .A3(_08323_),
    .B1(_08307_),
    .X(_08527_));
 sky130_fd_sc_hd__and2_1 _15433_ (.A(_08315_),
    .B(_08316_),
    .X(_08528_));
 sky130_fd_sc_hd__clkbuf_4 _15434_ (.A(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__o22a_1 _15435_ (.A1(_08127_),
    .A2(_08142_),
    .B1(_08529_),
    .B2(_08338_),
    .X(_08530_));
 sky130_fd_sc_hd__or3b_1 _15436_ (.A(_08529_),
    .B(_08142_),
    .C_N(_08132_),
    .X(_08531_));
 sky130_fd_sc_hd__or2b_1 _15437_ (.A(_08530_),
    .B_N(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__nand2_1 _15438_ (.A(net8267),
    .B(_08129_),
    .Y(_08533_));
 sky130_fd_sc_hd__or2_1 _15439_ (.A(_06122_),
    .B(net8008),
    .X(_08534_));
 sky130_fd_sc_hd__buf_2 _15440_ (.A(_08534_),
    .X(_08535_));
 sky130_fd_sc_hd__nor2_1 _15441_ (.A(_08139_),
    .B(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__xnor2_1 _15442_ (.A(_08532_),
    .B(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__xor2_1 _15443_ (.A(_08526_),
    .B(_08527_),
    .X(_08538_));
 sky130_fd_sc_hd__nand2_1 _15444_ (.A(_08537_),
    .B(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__o21ai_1 _15445_ (.A1(_08526_),
    .A2(_08527_),
    .B1(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__a32o_1 _15446_ (.A1(_08358_),
    .A2(_08514_),
    .A3(_08515_),
    .B1(_08517_),
    .B2(_08512_),
    .X(_08541_));
 sky130_fd_sc_hd__clkbuf_4 _15447_ (.A(_08277_),
    .X(_08542_));
 sky130_fd_sc_hd__clkbuf_4 _15448_ (.A(_08529_),
    .X(_08543_));
 sky130_fd_sc_hd__o22ai_2 _15449_ (.A1(_08338_),
    .A2(_08542_),
    .B1(_08543_),
    .B2(_08142_),
    .Y(_08544_));
 sky130_fd_sc_hd__or2_1 _15450_ (.A(_08142_),
    .B(_08277_),
    .X(_08545_));
 sky130_fd_sc_hd__nor3_1 _15451_ (.A(_08338_),
    .B(_08529_),
    .C(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__inv_2 _15452_ (.A(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand2_1 _15453_ (.A(_08544_),
    .B(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__nor2_1 _15454_ (.A(_08127_),
    .B(_08535_),
    .Y(_08549_));
 sky130_fd_sc_hd__xnor2_1 _15455_ (.A(_08548_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__or4_1 _15456_ (.A(_08207_),
    .B(_08229_),
    .C(_08294_),
    .D(_08305_),
    .X(_08551_));
 sky130_fd_sc_hd__o22ai_1 _15457_ (.A1(_08207_),
    .A2(_08294_),
    .B1(_08306_),
    .B2(_08229_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_1 _15458_ (.A(_08551_),
    .B(_08552_),
    .Y(_08553_));
 sky130_fd_sc_hd__or2_1 _15459_ (.A(_08255_),
    .B(_08323_),
    .X(_08554_));
 sky130_fd_sc_hd__xnor2_1 _15460_ (.A(_08553_),
    .B(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__nand2_1 _15461_ (.A(_08522_),
    .B(_08523_),
    .Y(_08556_));
 sky130_fd_sc_hd__o31a_1 _15462_ (.A1(_08280_),
    .A2(_08323_),
    .A3(_08524_),
    .B1(_08556_),
    .X(_08557_));
 sky130_fd_sc_hd__nor2_1 _15463_ (.A(_08555_),
    .B(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__and2_1 _15464_ (.A(_08555_),
    .B(_08557_),
    .X(_08559_));
 sky130_fd_sc_hd__nor2_1 _15465_ (.A(_08558_),
    .B(_08559_),
    .Y(_08560_));
 sky130_fd_sc_hd__xnor2_1 _15466_ (.A(_08550_),
    .B(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__xor2_1 _15467_ (.A(_08541_),
    .B(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__xnor2_1 _15468_ (.A(_08540_),
    .B(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__xnor2_1 _15469_ (.A(_08521_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__and3_1 _15470_ (.A(_08519_),
    .B(_08507_),
    .C(_08518_),
    .X(_08565_));
 sky130_fd_sc_hd__a21oi_1 _15471_ (.A1(_08519_),
    .A2(_08507_),
    .B1(_08518_),
    .Y(_08566_));
 sky130_fd_sc_hd__or2_4 _15472_ (.A(_08565_),
    .B(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__nand3_1 _15473_ (.A(_08505_),
    .B(_08499_),
    .C(_08504_),
    .Y(_08568_));
 sky130_fd_sc_hd__a21o_1 _15474_ (.A1(_08505_),
    .A2(_08499_),
    .B1(_08504_),
    .X(_08569_));
 sky130_fd_sc_hd__xnor2_4 _15475_ (.A(_08496_),
    .B(_08497_),
    .Y(_08570_));
 sky130_fd_sc_hd__or4b_2 _15476_ (.A(_08374_),
    .B(net4877),
    .C(_08494_),
    .D_N(_08366_),
    .X(_08571_));
 sky130_fd_sc_hd__nor2_1 _15477_ (.A(_06119_),
    .B(net8033),
    .Y(_08572_));
 sky130_fd_sc_hd__clkbuf_4 _15478_ (.A(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__a2bb2o_1 _15479_ (.A1_N(_08374_),
    .A2_N(net4877),
    .B1(_08573_),
    .B2(_08366_),
    .X(_08574_));
 sky130_fd_sc_hd__nor2_1 _15480_ (.A(_08384_),
    .B(_08458_),
    .Y(_08575_));
 sky130_fd_sc_hd__nand3_2 _15481_ (.A(_08571_),
    .B(_08574_),
    .C(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand2_2 _15482_ (.A(_08571_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__xnor2_4 _15483_ (.A(_08570_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__or4_1 _15484_ (.A(_08161_),
    .B(_08168_),
    .C(net8414),
    .D(_08384_),
    .X(_08579_));
 sky130_fd_sc_hd__o22ai_2 _15485_ (.A1(_08389_),
    .A2(net8414),
    .B1(_08392_),
    .B2(_08161_),
    .Y(_08580_));
 sky130_fd_sc_hd__nand2_2 _15486_ (.A(_08579_),
    .B(_08580_),
    .Y(_08581_));
 sky130_fd_sc_hd__nor2_2 _15487_ (.A(_08211_),
    .B(_08200_),
    .Y(_08582_));
 sky130_fd_sc_hd__xnor2_4 _15488_ (.A(_08581_),
    .B(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__and2b_1 _15489_ (.A_N(_08570_),
    .B(_08577_),
    .X(_08584_));
 sky130_fd_sc_hd__a21o_1 _15490_ (.A1(_08578_),
    .A2(_08583_),
    .B1(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__a21o_1 _15491_ (.A1(_08568_),
    .A2(_08569_),
    .B1(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__a21bo_2 _15492_ (.A1(_08247_),
    .A2(_08267_),
    .B1_N(_08242_),
    .X(_08587_));
 sky130_fd_sc_hd__a21bo_1 _15493_ (.A1(_08580_),
    .A2(_08582_),
    .B1_N(_08579_),
    .X(_08588_));
 sky130_fd_sc_hd__nand2_1 _15494_ (.A(_08511_),
    .B(_08508_),
    .Y(_08589_));
 sky130_fd_sc_hd__xnor2_2 _15495_ (.A(_08589_),
    .B(_08510_),
    .Y(_08590_));
 sky130_fd_sc_hd__xnor2_2 _15496_ (.A(_08588_),
    .B(_08590_),
    .Y(_08591_));
 sky130_fd_sc_hd__xnor2_4 _15497_ (.A(_08587_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__and3_1 _15498_ (.A(_08568_),
    .B(_08569_),
    .C(_08585_),
    .X(_08593_));
 sky130_fd_sc_hd__a21oi_2 _15499_ (.A1(_08586_),
    .A2(_08592_),
    .B1(_08593_),
    .Y(_08594_));
 sky130_fd_sc_hd__xor2_2 _15500_ (.A(_08567_),
    .B(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__nor2_1 _15501_ (.A(_08325_),
    .B(_08334_),
    .Y(_08596_));
 sky130_fd_sc_hd__a21o_1 _15502_ (.A1(_08287_),
    .A2(_08335_),
    .B1(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__or2b_1 _15503_ (.A(_08591_),
    .B_N(_08587_),
    .X(_08598_));
 sky130_fd_sc_hd__a21bo_1 _15504_ (.A1(_08588_),
    .A2(_08590_),
    .B1_N(_08598_),
    .X(_08599_));
 sky130_fd_sc_hd__or2_1 _15505_ (.A(_08537_),
    .B(_08538_),
    .X(_08600_));
 sky130_fd_sc_hd__nand2_1 _15506_ (.A(_08539_),
    .B(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__xor2_2 _15507_ (.A(_08599_),
    .B(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__xnor2_2 _15508_ (.A(_08597_),
    .B(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__nor2_1 _15509_ (.A(_08567_),
    .B(_08594_),
    .Y(_08604_));
 sky130_fd_sc_hd__a21oi_2 _15510_ (.A1(_08595_),
    .A2(_08603_),
    .B1(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__nor2_2 _15511_ (.A(_08564_),
    .B(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__nand2_2 _15512_ (.A(_08605_),
    .B(_08564_),
    .Y(_08607_));
 sky130_fd_sc_hd__and2b_2 _15513_ (.A_N(_08606_),
    .B(_08607_),
    .X(_08608_));
 sky130_fd_sc_hd__or2b_1 _15514_ (.A(_08601_),
    .B_N(_08599_),
    .X(_08609_));
 sky130_fd_sc_hd__or2b_1 _15515_ (.A(_08602_),
    .B_N(_08597_),
    .X(_08610_));
 sky130_fd_sc_hd__clkbuf_4 _15516_ (.A(_08139_),
    .X(_08611_));
 sky130_fd_sc_hd__nand2_4 _15517_ (.A(net8265),
    .B(_08119_),
    .Y(_08612_));
 sky130_fd_sc_hd__or2_1 _15518_ (.A(_06121_),
    .B(_08612_),
    .X(_08613_));
 sky130_fd_sc_hd__clkbuf_4 _15519_ (.A(_08613_),
    .X(_08614_));
 sky130_fd_sc_hd__or2_1 _15520_ (.A(_08611_),
    .B(_08614_),
    .X(_08615_));
 sky130_fd_sc_hd__clkbuf_4 _15521_ (.A(_08535_),
    .X(_08616_));
 sky130_fd_sc_hd__o31a_1 _15522_ (.A1(_08611_),
    .A2(_08530_),
    .A3(_08616_),
    .B1(_08531_),
    .X(_08617_));
 sky130_fd_sc_hd__nor2_1 _15523_ (.A(_08615_),
    .B(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__and2_1 _15524_ (.A(_08615_),
    .B(_08617_),
    .X(_08619_));
 sky130_fd_sc_hd__or2_1 _15525_ (.A(_08618_),
    .B(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__a21oi_2 _15526_ (.A1(_08609_),
    .A2(_08610_),
    .B1(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__and3_1 _15527_ (.A(_08609_),
    .B(_08610_),
    .C(_08620_),
    .X(_08622_));
 sky130_fd_sc_hd__nor2_2 _15528_ (.A(_08621_),
    .B(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__xnor2_4 _15529_ (.A(_08608_),
    .B(_08623_),
    .Y(_08624_));
 sky130_fd_sc_hd__xnor2_2 _15530_ (.A(_08595_),
    .B(_08603_),
    .Y(_08625_));
 sky130_fd_sc_hd__and2b_1 _15531_ (.A_N(_08593_),
    .B(_08586_),
    .X(_08626_));
 sky130_fd_sc_hd__xnor2_4 _15532_ (.A(_08626_),
    .B(_08592_),
    .Y(_08627_));
 sky130_fd_sc_hd__xnor2_4 _15533_ (.A(_08578_),
    .B(_08583_),
    .Y(_08628_));
 sky130_fd_sc_hd__a21o_1 _15534_ (.A1(_08571_),
    .A2(_08574_),
    .B1(_08575_),
    .X(_08629_));
 sky130_fd_sc_hd__or4_2 _15535_ (.A(net8041),
    .B(_08124_),
    .C(_08381_),
    .D(_08382_),
    .X(_08630_));
 sky130_fd_sc_hd__or4_1 _15536_ (.A(_08372_),
    .B(_08373_),
    .C(net4877),
    .D(_08630_),
    .X(_08631_));
 sky130_fd_sc_hd__o211a_1 _15537_ (.A1(net3626),
    .A2(_08162_),
    .B1(_08167_),
    .C1(_08433_),
    .X(_08632_));
 sky130_fd_sc_hd__o32ai_2 _15538_ (.A1(_08372_),
    .A2(_08373_),
    .A3(net8033),
    .B1(net4877),
    .B2(_08383_),
    .Y(_08633_));
 sky130_fd_sc_hd__nand3_1 _15539_ (.A(_08631_),
    .B(_08632_),
    .C(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand2_1 _15540_ (.A(_08631_),
    .B(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__nand3_2 _15541_ (.A(_08576_),
    .B(_08629_),
    .C(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__a21o_1 _15542_ (.A1(_08576_),
    .A2(_08629_),
    .B1(_08635_),
    .X(_08637_));
 sky130_fd_sc_hd__nand2_1 _15543_ (.A(_08212_),
    .B(_08187_),
    .Y(_08638_));
 sky130_fd_sc_hd__xnor2_1 _15544_ (.A(_08638_),
    .B(_08208_),
    .Y(_08639_));
 sky130_fd_sc_hd__nand3_1 _15545_ (.A(_08636_),
    .B(_08637_),
    .C(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__and2_2 _15546_ (.A(_08636_),
    .B(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__xor2_4 _15547_ (.A(_08628_),
    .B(_08641_),
    .X(_08642_));
 sky130_fd_sc_hd__xnor2_4 _15548_ (.A(_08283_),
    .B(_08269_),
    .Y(_08643_));
 sky130_fd_sc_hd__nor2_1 _15549_ (.A(_08628_),
    .B(_08641_),
    .Y(_08644_));
 sky130_fd_sc_hd__a21oi_4 _15550_ (.A1(_08642_),
    .A2(_08643_),
    .B1(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__xor2_4 _15551_ (.A(_08627_),
    .B(_08645_),
    .X(_08646_));
 sky130_fd_sc_hd__xnor2_4 _15552_ (.A(_08350_),
    .B(_08337_),
    .Y(_08647_));
 sky130_fd_sc_hd__nor2_1 _15553_ (.A(_08627_),
    .B(_08645_),
    .Y(_08648_));
 sky130_fd_sc_hd__a21oi_2 _15554_ (.A1(_08646_),
    .A2(_08647_),
    .B1(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__xor2_1 _15555_ (.A(_08625_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__nand2_1 _15556_ (.A(_08144_),
    .B(_08352_),
    .Y(_08651_));
 sky130_fd_sc_hd__and2_1 _15557_ (.A(_08353_),
    .B(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__nand2_2 _15558_ (.A(_08650_),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__o21ai_4 _15559_ (.A1(_08625_),
    .A2(_08649_),
    .B1(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__xnor2_4 _15560_ (.A(_08624_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__xnor2_4 _15561_ (.A(_08354_),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__xnor2_4 _15562_ (.A(_08646_),
    .B(_08647_),
    .Y(_08657_));
 sky130_fd_sc_hd__xnor2_4 _15563_ (.A(_08642_),
    .B(_08643_),
    .Y(_08658_));
 sky130_fd_sc_hd__a21o_1 _15564_ (.A1(_08636_),
    .A2(_08637_),
    .B1(_08639_),
    .X(_08659_));
 sky130_fd_sc_hd__a21o_1 _15565_ (.A1(_08631_),
    .A2(_08633_),
    .B1(_08632_),
    .X(_08660_));
 sky130_fd_sc_hd__a21oi_4 _15566_ (.A1(_08118_),
    .A2(_08164_),
    .B1(_08165_),
    .Y(_08661_));
 sky130_fd_sc_hd__o21ai_1 _15567_ (.A1(_08661_),
    .A2(_08474_),
    .B1(_08630_),
    .Y(_08662_));
 sky130_fd_sc_hd__and3b_1 _15568_ (.A_N(_08630_),
    .B(_08167_),
    .C(_08464_),
    .X(_08663_));
 sky130_fd_sc_hd__a31o_1 _15569_ (.A1(_08186_),
    .A2(_08433_),
    .A3(_08662_),
    .B1(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__nand3_1 _15570_ (.A(_08634_),
    .B(_08660_),
    .C(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__o2bb2a_4 _15571_ (.A1_N(_08199_),
    .A2_N(_08195_),
    .B1(net8425),
    .B2(_08192_),
    .X(_08666_));
 sky130_fd_sc_hd__nand2_1 _15572_ (.A(_08666_),
    .B(_08245_),
    .Y(_08667_));
 sky130_fd_sc_hd__o2bb2a_1 _15573_ (.A1_N(_08159_),
    .A2_N(_08157_),
    .B1(net7835),
    .B2(_08147_),
    .X(_08668_));
 sky130_fd_sc_hd__o211a_1 _15574_ (.A1(net3637),
    .A2(_08162_),
    .B1(net7836),
    .C1(_08185_),
    .X(_08669_));
 sky130_fd_sc_hd__and3_1 _15575_ (.A(_08180_),
    .B(_08204_),
    .C(_08205_),
    .X(_08670_));
 sky130_fd_sc_hd__xor2_1 _15576_ (.A(_08669_),
    .B(_08670_),
    .X(_08671_));
 sky130_fd_sc_hd__xnor2_1 _15577_ (.A(_08667_),
    .B(_08671_),
    .Y(_08672_));
 sky130_fd_sc_hd__a21o_1 _15578_ (.A1(_08634_),
    .A2(_08660_),
    .B1(_08664_),
    .X(_08673_));
 sky130_fd_sc_hd__nand3_1 _15579_ (.A(_08665_),
    .B(_08672_),
    .C(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand2_1 _15580_ (.A(_08665_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__nand3_1 _15581_ (.A(_08640_),
    .B(_08659_),
    .C(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__a21o_1 _15582_ (.A1(_08640_),
    .A2(_08659_),
    .B1(_08675_),
    .X(_08677_));
 sky130_fd_sc_hd__or3_1 _15583_ (.A(_08240_),
    .B(_08277_),
    .C(_08278_),
    .X(_08678_));
 sky130_fd_sc_hd__or4b_1 _15584_ (.A(_08220_),
    .B(_08678_),
    .C(_08271_),
    .D_N(_08252_),
    .X(_08679_));
 sky130_fd_sc_hd__nor2_1 _15585_ (.A(_08277_),
    .B(_08278_),
    .Y(_08680_));
 sky130_fd_sc_hd__a32o_1 _15586_ (.A1(_08244_),
    .A2(_08252_),
    .A3(_08254_),
    .B1(_08680_),
    .B2(_08246_),
    .X(_08681_));
 sky130_fd_sc_hd__or4bb_2 _15587_ (.A(_08266_),
    .B(_08317_),
    .C_N(_08679_),
    .D_N(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__nand2_1 _15588_ (.A(_08679_),
    .B(_08682_),
    .Y(_08683_));
 sky130_fd_sc_hd__a32o_1 _15589_ (.A1(_08666_),
    .A2(_08245_),
    .A3(_08671_),
    .B1(_08670_),
    .B2(_08669_),
    .X(_08684_));
 sky130_fd_sc_hd__xnor2_1 _15590_ (.A(_08273_),
    .B(_08281_),
    .Y(_08685_));
 sky130_fd_sc_hd__xor2_1 _15591_ (.A(_08684_),
    .B(_08685_),
    .X(_08686_));
 sky130_fd_sc_hd__xnor2_1 _15592_ (.A(_08683_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__nand3_1 _15593_ (.A(_08676_),
    .B(_08677_),
    .C(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__and2_2 _15594_ (.A(_08676_),
    .B(_08688_),
    .X(_08689_));
 sky130_fd_sc_hd__xor2_4 _15595_ (.A(_08658_),
    .B(_08689_),
    .X(_08690_));
 sky130_fd_sc_hd__clkbuf_4 _15596_ (.A(_08341_),
    .X(_08691_));
 sky130_fd_sc_hd__or4_4 _15597_ (.A(_08308_),
    .B(_08309_),
    .C(_08329_),
    .D(_08691_),
    .X(_08692_));
 sky130_fd_sc_hd__xor2_2 _15598_ (.A(_08342_),
    .B(_08345_),
    .X(_08693_));
 sky130_fd_sc_hd__or2b_2 _15599_ (.A(_08692_),
    .B_N(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__or2b_1 _15600_ (.A(_08685_),
    .B_N(_08684_),
    .X(_08695_));
 sky130_fd_sc_hd__or2b_1 _15601_ (.A(_08686_),
    .B_N(_08683_),
    .X(_08696_));
 sky130_fd_sc_hd__nand2_2 _15602_ (.A(_08695_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__and2b_1 _15603_ (.A_N(_08349_),
    .B(_08348_),
    .X(_08698_));
 sky130_fd_sc_hd__xnor2_4 _15604_ (.A(_08339_),
    .B(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__xnor2_4 _15605_ (.A(_08697_),
    .B(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__xnor2_4 _15606_ (.A(_08694_),
    .B(_08700_),
    .Y(_08701_));
 sky130_fd_sc_hd__nor2_1 _15607_ (.A(_08658_),
    .B(_08689_),
    .Y(_08702_));
 sky130_fd_sc_hd__a21oi_4 _15608_ (.A1(_08690_),
    .A2(_08701_),
    .B1(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__xnor2_4 _15609_ (.A(_08657_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__and2b_1 _15610_ (.A_N(_08699_),
    .B(_08697_),
    .X(_08705_));
 sky130_fd_sc_hd__and2b_1 _15611_ (.A_N(_08694_),
    .B(_08700_),
    .X(_08706_));
 sky130_fd_sc_hd__nor2_2 _15612_ (.A(_08705_),
    .B(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__xnor2_4 _15613_ (.A(_08704_),
    .B(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__and3_1 _15614_ (.A(net7836),
    .B(_08204_),
    .C(_08205_),
    .X(_08709_));
 sky130_fd_sc_hd__or3_1 _15615_ (.A(net8414),
    .B(_08225_),
    .C(_08227_),
    .X(_08710_));
 sky130_fd_sc_hd__xnor2_1 _15616_ (.A(_08709_),
    .B(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__and3_1 _15617_ (.A(_08180_),
    .B(_08245_),
    .C(_08709_),
    .X(_08712_));
 sky130_fd_sc_hd__a41o_1 _15618_ (.A1(_08666_),
    .A2(_08253_),
    .A3(_08254_),
    .A4(_08711_),
    .B1(_08712_),
    .X(_08713_));
 sky130_fd_sc_hd__a2bb2o_1 _15619_ (.A1_N(_08266_),
    .A2_N(_08318_),
    .B1(_08679_),
    .B2(_08681_),
    .X(_08714_));
 sky130_fd_sc_hd__nand3_2 _15620_ (.A(_08682_),
    .B(_08713_),
    .C(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__or4_1 _15621_ (.A(_08220_),
    .B(_08240_),
    .C(_08279_),
    .D(_08317_),
    .X(_08716_));
 sky130_fd_sc_hd__nor2_1 _15622_ (.A(_08266_),
    .B(_08328_),
    .Y(_08717_));
 sky130_fd_sc_hd__o22ai_1 _15623_ (.A1(_08221_),
    .A2(_08279_),
    .B1(_08318_),
    .B2(_08241_),
    .Y(_08718_));
 sky130_fd_sc_hd__nand3_1 _15624_ (.A(_08716_),
    .B(_08717_),
    .C(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__nand2_1 _15625_ (.A(_08716_),
    .B(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__a21o_1 _15626_ (.A1(_08682_),
    .A2(_08714_),
    .B1(_08713_),
    .X(_08721_));
 sky130_fd_sc_hd__and2_1 _15627_ (.A(_08715_),
    .B(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__nand2_1 _15628_ (.A(_08720_),
    .B(_08722_),
    .Y(_08723_));
 sky130_fd_sc_hd__xor2_2 _15629_ (.A(_08692_),
    .B(_08693_),
    .X(_08724_));
 sky130_fd_sc_hd__a21oi_4 _15630_ (.A1(_08715_),
    .A2(_08723_),
    .B1(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__xnor2_4 _15631_ (.A(_08690_),
    .B(_08701_),
    .Y(_08726_));
 sky130_fd_sc_hd__a21o_1 _15632_ (.A1(_08676_),
    .A2(_08677_),
    .B1(_08687_),
    .X(_08727_));
 sky130_fd_sc_hd__a21o_1 _15633_ (.A1(_08665_),
    .A2(_08673_),
    .B1(_08672_),
    .X(_08728_));
 sky130_fd_sc_hd__or4b_1 _15634_ (.A(_08210_),
    .B(_08457_),
    .C(_08663_),
    .D_N(_08662_),
    .X(_08729_));
 sky130_fd_sc_hd__or3_1 _15635_ (.A(_08661_),
    .B(_08473_),
    .C(_08630_),
    .X(_08730_));
 sky130_fd_sc_hd__a22o_1 _15636_ (.A1(_08186_),
    .A2(_08433_),
    .B1(_08730_),
    .B2(_08662_),
    .X(_08731_));
 sky130_fd_sc_hd__a22o_1 _15637_ (.A1(_08185_),
    .A2(_08463_),
    .B1(_08572_),
    .B2(_08166_),
    .X(_08732_));
 sky130_fd_sc_hd__and4_1 _15638_ (.A(_08166_),
    .B(_08185_),
    .C(_08463_),
    .D(_08572_),
    .X(_08733_));
 sky130_fd_sc_hd__a31o_1 _15639_ (.A1(_08243_),
    .A2(_08433_),
    .A3(_08732_),
    .B1(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__nand3_2 _15640_ (.A(_08729_),
    .B(_08731_),
    .C(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__or3b_1 _15641_ (.A(_08271_),
    .B(_08200_),
    .C_N(_08252_),
    .X(_08736_));
 sky130_fd_sc_hd__xnor2_1 _15642_ (.A(_08736_),
    .B(_08711_),
    .Y(_08737_));
 sky130_fd_sc_hd__a21o_1 _15643_ (.A1(_08729_),
    .A2(_08731_),
    .B1(_08734_),
    .X(_08738_));
 sky130_fd_sc_hd__nand3_1 _15644_ (.A(_08735_),
    .B(_08737_),
    .C(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__nand2_1 _15645_ (.A(_08735_),
    .B(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__xor2_2 _15646_ (.A(_08720_),
    .B(_08722_),
    .X(_08741_));
 sky130_fd_sc_hd__nand2_1 _15647_ (.A(_08674_),
    .B(_08728_),
    .Y(_08742_));
 sky130_fd_sc_hd__xnor2_2 _15648_ (.A(_08742_),
    .B(_08740_),
    .Y(_08743_));
 sky130_fd_sc_hd__a32o_1 _15649_ (.A1(_08674_),
    .A2(_08728_),
    .A3(_08740_),
    .B1(_08741_),
    .B2(_08743_),
    .X(_08744_));
 sky130_fd_sc_hd__nand3_1 _15650_ (.A(_08688_),
    .B(_08727_),
    .C(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__a21o_1 _15651_ (.A1(_08688_),
    .A2(_08727_),
    .B1(_08744_),
    .X(_08746_));
 sky130_fd_sc_hd__and3_1 _15652_ (.A(_08715_),
    .B(_08723_),
    .C(_08724_),
    .X(_08747_));
 sky130_fd_sc_hd__nor2_1 _15653_ (.A(_08725_),
    .B(_08747_),
    .Y(_08748_));
 sky130_fd_sc_hd__nand3_1 _15654_ (.A(_08745_),
    .B(_08746_),
    .C(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__and2_2 _15655_ (.A(_08745_),
    .B(_08749_),
    .X(_08750_));
 sky130_fd_sc_hd__xor2_4 _15656_ (.A(_08726_),
    .B(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__nor2_1 _15657_ (.A(_08726_),
    .B(_08750_),
    .Y(_08752_));
 sky130_fd_sc_hd__a21oi_2 _15658_ (.A1(_08725_),
    .A2(_08751_),
    .B1(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__nor2_1 _15659_ (.A(_08708_),
    .B(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__or2_1 _15660_ (.A(_08650_),
    .B(_08652_),
    .X(_08755_));
 sky130_fd_sc_hd__nand2_1 _15661_ (.A(_08653_),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__or2_1 _15662_ (.A(_08657_),
    .B(_08703_),
    .X(_08757_));
 sky130_fd_sc_hd__o21a_1 _15663_ (.A1(_08704_),
    .A2(_08707_),
    .B1(_08757_),
    .X(_08758_));
 sky130_fd_sc_hd__nor2_1 _15664_ (.A(_08756_),
    .B(_08758_),
    .Y(_08759_));
 sky130_fd_sc_hd__nand2_1 _15665_ (.A(_08756_),
    .B(_08758_),
    .Y(_08760_));
 sky130_fd_sc_hd__nor2b_2 _15666_ (.A(_08759_),
    .B_N(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__nand2_1 _15667_ (.A(_08754_),
    .B(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__xnor2_4 _15668_ (.A(_08725_),
    .B(_08751_),
    .Y(_08763_));
 sky130_fd_sc_hd__a21o_1 _15669_ (.A1(_08745_),
    .A2(_08746_),
    .B1(_08748_),
    .X(_08764_));
 sky130_fd_sc_hd__xor2_2 _15670_ (.A(_08741_),
    .B(_08743_),
    .X(_08765_));
 sky130_fd_sc_hd__a21o_1 _15671_ (.A1(_08735_),
    .A2(_08738_),
    .B1(_08737_),
    .X(_08766_));
 sky130_fd_sc_hd__or4b_1 _15672_ (.A(_08206_),
    .B(_08457_),
    .C(_08733_),
    .D_N(_08732_),
    .X(_08767_));
 sky130_fd_sc_hd__or4b_1 _15673_ (.A(_08661_),
    .B(_08473_),
    .C(_08494_),
    .D_N(_08185_),
    .X(_08768_));
 sky130_fd_sc_hd__a22o_1 _15674_ (.A1(_08243_),
    .A2(_08433_),
    .B1(_08768_),
    .B2(_08732_),
    .X(_08769_));
 sky130_fd_sc_hd__a22o_1 _15675_ (.A1(_08204_),
    .A2(_08464_),
    .B1(_08573_),
    .B2(_08185_),
    .X(_08770_));
 sky130_fd_sc_hd__and4_1 _15676_ (.A(_08185_),
    .B(_08204_),
    .C(_08464_),
    .D(_08573_),
    .X(_08771_));
 sky130_fd_sc_hd__a31o_1 _15677_ (.A1(_08245_),
    .A2(_08433_),
    .A3(_08770_),
    .B1(_08771_),
    .X(_08772_));
 sky130_fd_sc_hd__nor2_1 _15678_ (.A(_08200_),
    .B(_08280_),
    .Y(_08773_));
 sky130_fd_sc_hd__or3_1 _15679_ (.A(_08160_),
    .B(_08225_),
    .C(_08227_),
    .X(_08774_));
 sky130_fd_sc_hd__or4b_1 _15680_ (.A(net8414),
    .B(_08774_),
    .C(_08271_),
    .D_N(_08252_),
    .X(_08775_));
 sky130_fd_sc_hd__a32o_1 _15681_ (.A1(_08180_),
    .A2(_08252_),
    .A3(_08254_),
    .B1(_08245_),
    .B2(net7836),
    .X(_08776_));
 sky130_fd_sc_hd__nand2_1 _15682_ (.A(_08775_),
    .B(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__xnor2_1 _15683_ (.A(_08773_),
    .B(_08777_),
    .Y(_08778_));
 sky130_fd_sc_hd__nand2_1 _15684_ (.A(_08767_),
    .B(_08769_),
    .Y(_08779_));
 sky130_fd_sc_hd__xnor2_1 _15685_ (.A(_08779_),
    .B(_08772_),
    .Y(_08780_));
 sky130_fd_sc_hd__a32o_1 _15686_ (.A1(_08767_),
    .A2(_08769_),
    .A3(_08772_),
    .B1(_08778_),
    .B2(_08780_),
    .X(_08781_));
 sky130_fd_sc_hd__or2_1 _15687_ (.A(_08266_),
    .B(_08341_),
    .X(_08782_));
 sky130_fd_sc_hd__nor2_1 _15688_ (.A(_08220_),
    .B(_08317_),
    .Y(_08783_));
 sky130_fd_sc_hd__nor2_1 _15689_ (.A(_08241_),
    .B(_08328_),
    .Y(_08784_));
 sky130_fd_sc_hd__xnor2_1 _15690_ (.A(_08783_),
    .B(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__nand2_1 _15691_ (.A(_08783_),
    .B(_08784_),
    .Y(_08786_));
 sky130_fd_sc_hd__o21ai_1 _15692_ (.A1(_08782_),
    .A2(_08785_),
    .B1(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__a21bo_1 _15693_ (.A1(_08773_),
    .A2(_08776_),
    .B1_N(_08775_),
    .X(_08788_));
 sky130_fd_sc_hd__a21o_1 _15694_ (.A1(_08716_),
    .A2(_08718_),
    .B1(_08717_),
    .X(_08789_));
 sky130_fd_sc_hd__nand3_1 _15695_ (.A(_08719_),
    .B(_08788_),
    .C(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__a21o_1 _15696_ (.A1(_08719_),
    .A2(_08789_),
    .B1(_08788_),
    .X(_08791_));
 sky130_fd_sc_hd__nand2_1 _15697_ (.A(_08790_),
    .B(_08791_),
    .Y(_08792_));
 sky130_fd_sc_hd__xnor2_1 _15698_ (.A(_08787_),
    .B(_08792_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand2_1 _15699_ (.A(_08739_),
    .B(_08766_),
    .Y(_08794_));
 sky130_fd_sc_hd__xnor2_1 _15700_ (.A(_08794_),
    .B(_08781_),
    .Y(_08795_));
 sky130_fd_sc_hd__a32o_1 _15701_ (.A1(_08739_),
    .A2(_08766_),
    .A3(_08781_),
    .B1(_08793_),
    .B2(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__xor2_1 _15702_ (.A(_08765_),
    .B(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__a21bo_1 _15703_ (.A1(_08787_),
    .A2(_08791_),
    .B1_N(_08790_),
    .X(_08798_));
 sky130_fd_sc_hd__buf_4 _15704_ (.A(_08309_),
    .X(_08799_));
 sky130_fd_sc_hd__o22ai_2 _15705_ (.A1(_08326_),
    .A2(_08329_),
    .B1(_08691_),
    .B2(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__nand2_1 _15706_ (.A(_08692_),
    .B(_08800_),
    .Y(_08801_));
 sky130_fd_sc_hd__xnor2_1 _15707_ (.A(_08798_),
    .B(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__nand2_1 _15708_ (.A(_08765_),
    .B(_08796_),
    .Y(_08803_));
 sky130_fd_sc_hd__a21bo_1 _15709_ (.A1(_08797_),
    .A2(_08802_),
    .B1_N(_08803_),
    .X(_08804_));
 sky130_fd_sc_hd__nand3_1 _15710_ (.A(_08749_),
    .B(_08764_),
    .C(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__and3_1 _15711_ (.A(_08692_),
    .B(_08798_),
    .C(_08800_),
    .X(_08806_));
 sky130_fd_sc_hd__a21o_1 _15712_ (.A1(_08749_),
    .A2(_08764_),
    .B1(_08804_),
    .X(_08807_));
 sky130_fd_sc_hd__nand3_1 _15713_ (.A(_08806_),
    .B(_08805_),
    .C(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__and2_2 _15714_ (.A(_08805_),
    .B(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__nor2_1 _15715_ (.A(_08763_),
    .B(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__xor2_4 _15716_ (.A(_08708_),
    .B(_08753_),
    .X(_08811_));
 sky130_fd_sc_hd__and2_1 _15717_ (.A(_08810_),
    .B(_08811_),
    .X(_08812_));
 sky130_fd_sc_hd__a21o_1 _15718_ (.A1(_08805_),
    .A2(_08807_),
    .B1(_08806_),
    .X(_08813_));
 sky130_fd_sc_hd__nor2_1 _15719_ (.A(_08200_),
    .B(_08318_),
    .Y(_08814_));
 sky130_fd_sc_hd__and3_1 _15720_ (.A(net7836),
    .B(_08252_),
    .C(_08254_),
    .X(_08815_));
 sky130_fd_sc_hd__nor2_1 _15721_ (.A(net8414),
    .B(_08279_),
    .Y(_08816_));
 sky130_fd_sc_hd__xor2_1 _15722_ (.A(_08815_),
    .B(_08816_),
    .X(_08817_));
 sky130_fd_sc_hd__nand2_1 _15723_ (.A(_08815_),
    .B(_08816_),
    .Y(_08818_));
 sky130_fd_sc_hd__a21boi_1 _15724_ (.A1(_08814_),
    .A2(_08817_),
    .B1_N(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__xnor2_1 _15725_ (.A(_08782_),
    .B(_08785_),
    .Y(_08820_));
 sky130_fd_sc_hd__xor2_1 _15726_ (.A(_08819_),
    .B(_08820_),
    .X(_08821_));
 sky130_fd_sc_hd__and4bb_1 _15727_ (.A_N(_08341_),
    .B_N(_08329_),
    .C(_08246_),
    .D(_08244_),
    .X(_08822_));
 sky130_fd_sc_hd__nor2_1 _15728_ (.A(_08819_),
    .B(_08820_),
    .Y(_08823_));
 sky130_fd_sc_hd__a21oi_1 _15729_ (.A1(_08821_),
    .A2(_08822_),
    .B1(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__nor2_1 _15730_ (.A(_08326_),
    .B(_08691_),
    .Y(_08825_));
 sky130_fd_sc_hd__and2b_1 _15731_ (.A_N(_08824_),
    .B(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__xor2_1 _15732_ (.A(_08797_),
    .B(_08802_),
    .X(_08827_));
 sky130_fd_sc_hd__and2b_1 _15733_ (.A_N(_08825_),
    .B(_08824_),
    .X(_08828_));
 sky130_fd_sc_hd__nor2_1 _15734_ (.A(_08826_),
    .B(_08828_),
    .Y(_08829_));
 sky130_fd_sc_hd__xnor2_1 _15735_ (.A(_08793_),
    .B(_08795_),
    .Y(_08830_));
 sky130_fd_sc_hd__xor2_1 _15736_ (.A(_08821_),
    .B(_08822_),
    .X(_08831_));
 sky130_fd_sc_hd__xnor2_1 _15737_ (.A(_08778_),
    .B(_08780_),
    .Y(_08832_));
 sky130_fd_sc_hd__xor2_1 _15738_ (.A(_08814_),
    .B(_08817_),
    .X(_08833_));
 sky130_fd_sc_hd__nor2_1 _15739_ (.A(_08229_),
    .B(_08458_),
    .Y(_08834_));
 sky130_fd_sc_hd__and2b_1 _15740_ (.A_N(_08771_),
    .B(_08770_),
    .X(_08835_));
 sky130_fd_sc_hd__xnor2_2 _15741_ (.A(_08834_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__nor2_1 _15742_ (.A(_08226_),
    .B(_08474_),
    .Y(_08837_));
 sky130_fd_sc_hd__and3_1 _15743_ (.A(_08253_),
    .B(_08254_),
    .C(_08433_),
    .X(_08838_));
 sky130_fd_sc_hd__nand2_1 _15744_ (.A(_08204_),
    .B(_08573_),
    .Y(_08839_));
 sky130_fd_sc_hd__xnor2_1 _15745_ (.A(_08839_),
    .B(_08837_),
    .Y(_08840_));
 sky130_fd_sc_hd__a32o_1 _15746_ (.A1(_08204_),
    .A2(_08573_),
    .A3(_08837_),
    .B1(_08838_),
    .B2(_08840_),
    .X(_08841_));
 sky130_fd_sc_hd__xnor2_1 _15747_ (.A(_08836_),
    .B(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__or2b_1 _15748_ (.A(_08836_),
    .B_N(_08841_),
    .X(_08843_));
 sky130_fd_sc_hd__a21boi_1 _15749_ (.A1(_08833_),
    .A2(_08842_),
    .B1_N(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__xor2_1 _15750_ (.A(_08832_),
    .B(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _15751_ (.A(_08832_),
    .B(_08844_),
    .Y(_08846_));
 sky130_fd_sc_hd__a21oi_1 _15752_ (.A1(_08831_),
    .A2(_08845_),
    .B1(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__xor2_1 _15753_ (.A(_08830_),
    .B(_08847_),
    .X(_08848_));
 sky130_fd_sc_hd__nor2_1 _15754_ (.A(_08830_),
    .B(_08847_),
    .Y(_08849_));
 sky130_fd_sc_hd__a21o_1 _15755_ (.A1(_08829_),
    .A2(_08848_),
    .B1(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__xor2_1 _15756_ (.A(_08827_),
    .B(_08850_),
    .X(_08851_));
 sky130_fd_sc_hd__nand2_1 _15757_ (.A(_08827_),
    .B(_08850_),
    .Y(_08852_));
 sky130_fd_sc_hd__a21bo_1 _15758_ (.A1(_08826_),
    .A2(_08851_),
    .B1_N(_08852_),
    .X(_08853_));
 sky130_fd_sc_hd__nand3_1 _15759_ (.A(_08808_),
    .B(_08813_),
    .C(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__xnor2_4 _15760_ (.A(_08763_),
    .B(_08809_),
    .Y(_08855_));
 sky130_fd_sc_hd__nor2_1 _15761_ (.A(_08854_),
    .B(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__a21o_1 _15762_ (.A1(_08808_),
    .A2(_08813_),
    .B1(_08853_),
    .X(_08857_));
 sky130_fd_sc_hd__and2_1 _15763_ (.A(_08854_),
    .B(_08857_),
    .X(_08858_));
 sky130_fd_sc_hd__xor2_1 _15764_ (.A(_08826_),
    .B(_08851_),
    .X(_08859_));
 sky130_fd_sc_hd__xnor2_1 _15765_ (.A(_08831_),
    .B(_08845_),
    .Y(_08860_));
 sky130_fd_sc_hd__xnor2_1 _15766_ (.A(_08833_),
    .B(_08842_),
    .Y(_08861_));
 sky130_fd_sc_hd__xor2_1 _15767_ (.A(_08838_),
    .B(_08840_),
    .X(_08862_));
 sky130_fd_sc_hd__nor2_1 _15768_ (.A(_08280_),
    .B(_08458_),
    .Y(_08863_));
 sky130_fd_sc_hd__a21o_4 _15769_ (.A1(_08129_),
    .A2(_08223_),
    .B1(_08224_),
    .X(_08864_));
 sky130_fd_sc_hd__a22o_1 _15770_ (.A1(_08253_),
    .A2(_08464_),
    .B1(_08573_),
    .B2(_08864_),
    .X(_08865_));
 sky130_fd_sc_hd__and4_1 _15771_ (.A(_08864_),
    .B(_08253_),
    .C(_08464_),
    .D(_08573_),
    .X(_08866_));
 sky130_fd_sc_hd__a21o_1 _15772_ (.A1(_08863_),
    .A2(_08865_),
    .B1(_08866_),
    .X(_08867_));
 sky130_fd_sc_hd__xor2_1 _15773_ (.A(_08862_),
    .B(_08867_),
    .X(_08868_));
 sky130_fd_sc_hd__or2_1 _15774_ (.A(_08417_),
    .B(_08329_),
    .X(_08869_));
 sky130_fd_sc_hd__o22a_1 _15775_ (.A1(_08161_),
    .A2(_08280_),
    .B1(_08318_),
    .B2(_08402_),
    .X(_08870_));
 sky130_fd_sc_hd__or4_1 _15776_ (.A(_08161_),
    .B(net8414),
    .C(_08279_),
    .D(_08318_),
    .X(_08871_));
 sky130_fd_sc_hd__or2b_1 _15777_ (.A(_08870_),
    .B_N(_08871_),
    .X(_08872_));
 sky130_fd_sc_hd__xor2_1 _15778_ (.A(_08869_),
    .B(_08872_),
    .X(_08873_));
 sky130_fd_sc_hd__and2_1 _15779_ (.A(_08862_),
    .B(_08867_),
    .X(_08874_));
 sky130_fd_sc_hd__a21oi_1 _15780_ (.A1(_08868_),
    .A2(_08873_),
    .B1(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__nor2_1 _15781_ (.A(_08861_),
    .B(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__and2_1 _15782_ (.A(_08861_),
    .B(_08875_),
    .X(_08877_));
 sky130_fd_sc_hd__nor2_1 _15783_ (.A(_08876_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__o21ai_2 _15784_ (.A1(_08869_),
    .A2(_08870_),
    .B1(_08871_),
    .Y(_08879_));
 sky130_fd_sc_hd__buf_2 _15785_ (.A(_08221_),
    .X(_08880_));
 sky130_fd_sc_hd__o22a_1 _15786_ (.A1(_08880_),
    .A2(_08329_),
    .B1(_08691_),
    .B2(_08391_),
    .X(_08881_));
 sky130_fd_sc_hd__or2_1 _15787_ (.A(_08822_),
    .B(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__xnor2_1 _15788_ (.A(_08879_),
    .B(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__a21oi_1 _15789_ (.A1(_08878_),
    .A2(_08883_),
    .B1(_08876_),
    .Y(_08884_));
 sky130_fd_sc_hd__or2_1 _15790_ (.A(_08860_),
    .B(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__or2b_1 _15791_ (.A(_08882_),
    .B_N(_08879_),
    .X(_08886_));
 sky130_fd_sc_hd__xnor2_1 _15792_ (.A(_08860_),
    .B(_08884_),
    .Y(_08887_));
 sky130_fd_sc_hd__or2_1 _15793_ (.A(_08886_),
    .B(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__xnor2_1 _15794_ (.A(_08829_),
    .B(_08848_),
    .Y(_08889_));
 sky130_fd_sc_hd__a21oi_1 _15795_ (.A1(_08885_),
    .A2(_08888_),
    .B1(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__and2_1 _15796_ (.A(_08859_),
    .B(_08890_),
    .X(_08891_));
 sky130_fd_sc_hd__nand2_1 _15797_ (.A(_08858_),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__and3_1 _15798_ (.A(_08854_),
    .B(_08857_),
    .C(_08891_),
    .X(_08893_));
 sky130_fd_sc_hd__a21oi_1 _15799_ (.A1(_08854_),
    .A2(_08857_),
    .B1(_08891_),
    .Y(_08894_));
 sky130_fd_sc_hd__a21o_1 _15800_ (.A1(_08885_),
    .A2(_08888_),
    .B1(_08889_),
    .X(_08895_));
 sky130_fd_sc_hd__xnor2_1 _15801_ (.A(_08868_),
    .B(_08873_),
    .Y(_08896_));
 sky130_fd_sc_hd__or2_1 _15802_ (.A(_08161_),
    .B(_08318_),
    .X(_08897_));
 sky130_fd_sc_hd__nor2_1 _15803_ (.A(_08402_),
    .B(_08328_),
    .Y(_08898_));
 sky130_fd_sc_hd__xnor2_1 _15804_ (.A(_08897_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__or3b_1 _15805_ (.A(_08417_),
    .B(_08691_),
    .C_N(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__o21bai_1 _15806_ (.A1(_08417_),
    .A2(_08691_),
    .B1_N(_08899_),
    .Y(_08901_));
 sky130_fd_sc_hd__and2_1 _15807_ (.A(_08900_),
    .B(_08901_),
    .X(_08902_));
 sky130_fd_sc_hd__or2b_1 _15808_ (.A(_08866_),
    .B_N(_08865_),
    .X(_08903_));
 sky130_fd_sc_hd__xnor2_1 _15809_ (.A(_08863_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__clkbuf_4 _15810_ (.A(_08458_),
    .X(_08905_));
 sky130_fd_sc_hd__nor2_1 _15811_ (.A(_08318_),
    .B(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__nor2_1 _15812_ (.A(_08277_),
    .B(_08474_),
    .Y(_08907_));
 sky130_fd_sc_hd__a21o_1 _15813_ (.A1(_08253_),
    .A2(_08573_),
    .B1(_08907_),
    .X(_08908_));
 sky130_fd_sc_hd__and4bb_1 _15814_ (.A_N(_08494_),
    .B_N(_08277_),
    .C(_08253_),
    .D(_08464_),
    .X(_08909_));
 sky130_fd_sc_hd__a21o_1 _15815_ (.A1(_08906_),
    .A2(_08908_),
    .B1(_08909_),
    .X(_08910_));
 sky130_fd_sc_hd__xor2_1 _15816_ (.A(_08904_),
    .B(_08910_),
    .X(_08911_));
 sky130_fd_sc_hd__and2_1 _15817_ (.A(_08904_),
    .B(_08910_),
    .X(_08912_));
 sky130_fd_sc_hd__a21oi_1 _15818_ (.A1(_08902_),
    .A2(_08911_),
    .B1(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__or2_1 _15819_ (.A(_08896_),
    .B(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__xor2_1 _15820_ (.A(_08896_),
    .B(_08913_),
    .X(_08915_));
 sky130_fd_sc_hd__clkbuf_4 _15821_ (.A(_08402_),
    .X(_08916_));
 sky130_fd_sc_hd__o31a_1 _15822_ (.A1(_08916_),
    .A2(_08329_),
    .A3(_08897_),
    .B1(_08900_),
    .X(_08917_));
 sky130_fd_sc_hd__buf_4 _15823_ (.A(_08880_),
    .X(_08918_));
 sky130_fd_sc_hd__nor2_1 _15824_ (.A(_08918_),
    .B(_08691_),
    .Y(_08919_));
 sky130_fd_sc_hd__and2b_1 _15825_ (.A_N(_08917_),
    .B(_08919_),
    .X(_08920_));
 sky130_fd_sc_hd__and2b_1 _15826_ (.A_N(_08919_),
    .B(_08917_),
    .X(_08921_));
 sky130_fd_sc_hd__nor2_1 _15827_ (.A(_08920_),
    .B(_08921_),
    .Y(_08922_));
 sky130_fd_sc_hd__nand2_1 _15828_ (.A(_08915_),
    .B(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__xnor2_1 _15829_ (.A(_08878_),
    .B(_08883_),
    .Y(_08924_));
 sky130_fd_sc_hd__a21oi_2 _15830_ (.A1(_08914_),
    .A2(_08923_),
    .B1(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__and3_1 _15831_ (.A(_08924_),
    .B(_08914_),
    .C(_08923_),
    .X(_08926_));
 sky130_fd_sc_hd__nor2_1 _15832_ (.A(_08925_),
    .B(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__and2_1 _15833_ (.A(_08920_),
    .B(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__nand2_1 _15834_ (.A(_08889_),
    .B(_08885_),
    .Y(_08929_));
 sky130_fd_sc_hd__nand2_1 _15835_ (.A(_08886_),
    .B(_08887_),
    .Y(_08930_));
 sky130_fd_sc_hd__and2_1 _15836_ (.A(_08888_),
    .B(_08930_),
    .X(_08931_));
 sky130_fd_sc_hd__o211a_1 _15837_ (.A1(_08925_),
    .A2(_08928_),
    .B1(_08929_),
    .C1(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__and3_1 _15838_ (.A(_08859_),
    .B(_08895_),
    .C(_08932_),
    .X(_08933_));
 sky130_fd_sc_hd__o21bai_1 _15839_ (.A1(_08893_),
    .A2(_08894_),
    .B1_N(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__a21bo_1 _15840_ (.A1(_08925_),
    .A2(_08930_),
    .B1_N(_08929_),
    .X(_08935_));
 sky130_fd_sc_hd__nand2_1 _15841_ (.A(_08888_),
    .B(_08935_),
    .Y(_08936_));
 sky130_fd_sc_hd__or2_1 _15842_ (.A(_08915_),
    .B(_08922_),
    .X(_08937_));
 sky130_fd_sc_hd__and2_1 _15843_ (.A(_08923_),
    .B(_08937_),
    .X(_08938_));
 sky130_fd_sc_hd__xnor2_1 _15844_ (.A(_08902_),
    .B(_08911_),
    .Y(_08939_));
 sky130_fd_sc_hd__and2b_1 _15845_ (.A_N(_08909_),
    .B(_08908_),
    .X(_08940_));
 sky130_fd_sc_hd__xnor2_1 _15846_ (.A(_08906_),
    .B(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__nor2_1 _15847_ (.A(_08529_),
    .B(_08494_),
    .Y(_08942_));
 sky130_fd_sc_hd__or2_1 _15848_ (.A(_08329_),
    .B(_08458_),
    .X(_08943_));
 sky130_fd_sc_hd__o22a_1 _15849_ (.A1(_08529_),
    .A2(_08474_),
    .B1(_08494_),
    .B2(_08277_),
    .X(_08944_));
 sky130_fd_sc_hd__o2bb2a_1 _15850_ (.A1_N(_08907_),
    .A2_N(_08942_),
    .B1(_08943_),
    .B2(_08944_),
    .X(_08945_));
 sky130_fd_sc_hd__xor2_1 _15851_ (.A(_08941_),
    .B(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__and4bb_1 _15852_ (.A_N(_08691_),
    .B_N(_08329_),
    .C(net8423),
    .D(net7836),
    .X(_08947_));
 sky130_fd_sc_hd__clkbuf_4 _15853_ (.A(_08401_),
    .X(_08948_));
 sky130_fd_sc_hd__o22a_1 _15854_ (.A1(_08948_),
    .A2(_08329_),
    .B1(_08691_),
    .B2(_08916_),
    .X(_08949_));
 sky130_fd_sc_hd__nor2_1 _15855_ (.A(_08947_),
    .B(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__nand2_1 _15856_ (.A(_08946_),
    .B(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__o21a_1 _15857_ (.A1(_08941_),
    .A2(_08945_),
    .B1(_08951_),
    .X(_08952_));
 sky130_fd_sc_hd__xor2_1 _15858_ (.A(_08939_),
    .B(_08952_),
    .X(_08953_));
 sky130_fd_sc_hd__nand2_1 _15859_ (.A(_08947_),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__o21ai_1 _15860_ (.A1(_08939_),
    .A2(_08952_),
    .B1(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__or2_1 _15861_ (.A(_08946_),
    .B(_08950_),
    .X(_08956_));
 sky130_fd_sc_hd__or2_1 _15862_ (.A(_08948_),
    .B(_08691_),
    .X(_08957_));
 sky130_fd_sc_hd__nor2_1 _15863_ (.A(_08341_),
    .B(_08905_),
    .Y(_08958_));
 sky130_fd_sc_hd__nor2_1 _15864_ (.A(_08126_),
    .B(_08474_),
    .Y(_08959_));
 sky130_fd_sc_hd__xor2_1 _15865_ (.A(_08942_),
    .B(_08959_),
    .X(_08960_));
 sky130_fd_sc_hd__nand2_1 _15866_ (.A(_08958_),
    .B(_08960_),
    .Y(_08961_));
 sky130_fd_sc_hd__and4b_1 _15867_ (.A_N(_08139_),
    .B(net8042),
    .C(_08959_),
    .D(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__o21ai_1 _15868_ (.A1(_08958_),
    .A2(_08960_),
    .B1(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__a21oi_1 _15869_ (.A1(_08907_),
    .A2(_08942_),
    .B1(_08944_),
    .Y(_08964_));
 sky130_fd_sc_hd__xnor2_1 _15870_ (.A(_08943_),
    .B(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__a21bo_1 _15871_ (.A1(_08942_),
    .A2(_08959_),
    .B1_N(_08961_),
    .X(_08966_));
 sky130_fd_sc_hd__o2bb2a_1 _15872_ (.A1_N(_08957_),
    .A2_N(_08963_),
    .B1(_08965_),
    .B2(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__and2_1 _15873_ (.A(_08965_),
    .B(_08966_),
    .X(_08968_));
 sky130_fd_sc_hd__nor2_1 _15874_ (.A(_08957_),
    .B(_08963_),
    .Y(_08969_));
 sky130_fd_sc_hd__or3_1 _15875_ (.A(_08967_),
    .B(_08968_),
    .C(_08969_),
    .X(_08970_));
 sky130_fd_sc_hd__a32o_1 _15876_ (.A1(_08951_),
    .A2(_08956_),
    .A3(_08970_),
    .B1(_08969_),
    .B2(_08968_),
    .X(_08971_));
 sky130_fd_sc_hd__and2_1 _15877_ (.A(_08954_),
    .B(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__o221a_1 _15878_ (.A1(_08947_),
    .A2(_08953_),
    .B1(_08955_),
    .B2(_08938_),
    .C1(_08972_),
    .X(_08973_));
 sky130_fd_sc_hd__a21o_1 _15879_ (.A1(_08938_),
    .A2(_08955_),
    .B1(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__nor2_1 _15880_ (.A(_08920_),
    .B(_08927_),
    .Y(_08975_));
 sky130_fd_sc_hd__nor2_1 _15881_ (.A(_08928_),
    .B(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__o2111a_1 _15882_ (.A1(_08925_),
    .A2(_08931_),
    .B1(_08974_),
    .C1(_08976_),
    .D1(_08895_),
    .X(_08977_));
 sky130_fd_sc_hd__and3_1 _15883_ (.A(_08859_),
    .B(_08936_),
    .C(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__and4_1 _15884_ (.A(_08858_),
    .B(_08859_),
    .C(_08895_),
    .D(_08932_),
    .X(_08979_));
 sky130_fd_sc_hd__a21oi_2 _15885_ (.A1(_08934_),
    .A2(_08978_),
    .B1(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__a31o_1 _15886_ (.A1(_08808_),
    .A2(_08813_),
    .A3(_08853_),
    .B1(_08893_),
    .X(_08981_));
 sky130_fd_sc_hd__xor2_2 _15887_ (.A(_08855_),
    .B(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__o22ai_4 _15888_ (.A1(_08855_),
    .A2(_08892_),
    .B1(_08980_),
    .B2(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__nor2_2 _15889_ (.A(_08810_),
    .B(_08856_),
    .Y(_08984_));
 sky130_fd_sc_hd__xnor2_4 _15890_ (.A(_08811_),
    .B(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__a22o_2 _15891_ (.A1(_08811_),
    .A2(_08856_),
    .B1(_08983_),
    .B2(_08985_),
    .X(_08986_));
 sky130_fd_sc_hd__nor2_2 _15892_ (.A(_08754_),
    .B(_08812_),
    .Y(_08987_));
 sky130_fd_sc_hd__xnor2_4 _15893_ (.A(_08761_),
    .B(_08987_),
    .Y(_08988_));
 sky130_fd_sc_hd__a22o_4 _15894_ (.A1(_08761_),
    .A2(_08812_),
    .B1(_08986_),
    .B2(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__a21o_1 _15895_ (.A1(_08754_),
    .A2(_08760_),
    .B1(_08759_),
    .X(_08990_));
 sky130_fd_sc_hd__xnor2_4 _15896_ (.A(_08656_),
    .B(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__a2bb2o_4 _15897_ (.A1_N(_08656_),
    .A2_N(_08762_),
    .B1(_08989_),
    .B2(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__a21o_1 _15898_ (.A1(_08550_),
    .A2(_08560_),
    .B1(_08558_),
    .X(_08993_));
 sky130_fd_sc_hd__or2b_1 _15899_ (.A(_08399_),
    .B_N(_08359_),
    .X(_08994_));
 sky130_fd_sc_hd__or4b_1 _15900_ (.A(_08131_),
    .B(_08277_),
    .C(_08142_),
    .D_N(_08253_),
    .X(_08995_));
 sky130_fd_sc_hd__nor2_2 _15901_ (.A(_06122_),
    .B(net4918),
    .Y(_08996_));
 sky130_fd_sc_hd__a21bo_1 _15902_ (.A1(_08996_),
    .A2(_08253_),
    .B1_N(_08545_),
    .X(_08997_));
 sky130_fd_sc_hd__nand2_1 _15903_ (.A(_08995_),
    .B(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__or3_1 _15904_ (.A(_08529_),
    .B(_08535_),
    .C(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__o21ai_1 _15905_ (.A1(_08543_),
    .A2(_08535_),
    .B1(_08998_),
    .Y(_09000_));
 sky130_fd_sc_hd__and2_1 _15906_ (.A(_08999_),
    .B(_09000_),
    .X(_09001_));
 sky130_fd_sc_hd__or4_1 _15907_ (.A(_08211_),
    .B(_08207_),
    .C(_08294_),
    .D(_08305_),
    .X(_09002_));
 sky130_fd_sc_hd__o22ai_1 _15908_ (.A1(_08211_),
    .A2(_08294_),
    .B1(_08306_),
    .B2(_08207_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand2_1 _15909_ (.A(_09002_),
    .B(_09003_),
    .Y(_09004_));
 sky130_fd_sc_hd__or2_1 _15910_ (.A(_08229_),
    .B(_08322_),
    .X(_09005_));
 sky130_fd_sc_hd__xnor2_1 _15911_ (.A(_09004_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__o31a_1 _15912_ (.A1(_08255_),
    .A2(_08323_),
    .A3(_08553_),
    .B1(_08551_),
    .X(_09007_));
 sky130_fd_sc_hd__nor2_1 _15913_ (.A(_09006_),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__and2_1 _15914_ (.A(_09006_),
    .B(_09007_),
    .X(_09009_));
 sky130_fd_sc_hd__nor2_1 _15915_ (.A(_09008_),
    .B(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__xnor2_1 _15916_ (.A(_09001_),
    .B(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__a21o_1 _15917_ (.A1(_08397_),
    .A2(_08994_),
    .B1(_09011_),
    .X(_09012_));
 sky130_fd_sc_hd__nand3_1 _15918_ (.A(_08397_),
    .B(_08994_),
    .C(_09011_),
    .Y(_09013_));
 sky130_fd_sc_hd__nand2_1 _15919_ (.A(_09012_),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__xnor2_1 _15920_ (.A(_08993_),
    .B(_09014_),
    .Y(_09015_));
 sky130_fd_sc_hd__a21bo_1 _15921_ (.A1(_08393_),
    .A2(_08395_),
    .B1_N(_08390_),
    .X(_09016_));
 sky130_fd_sc_hd__a21bo_1 _15922_ (.A1(_08415_),
    .A2(_08419_),
    .B1_N(_08412_),
    .X(_09017_));
 sky130_fd_sc_hd__or4_1 _15923_ (.A(_08221_),
    .B(_08241_),
    .C(_08418_),
    .D(_08392_),
    .X(_09018_));
 sky130_fd_sc_hd__a2bb2o_1 _15924_ (.A1_N(_08392_),
    .A2_N(_08391_),
    .B1(_08244_),
    .B2(_08386_),
    .X(_09019_));
 sky130_fd_sc_hd__nand2_1 _15925_ (.A(_09018_),
    .B(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__nor2_1 _15926_ (.A(_08389_),
    .B(_08509_),
    .Y(_09021_));
 sky130_fd_sc_hd__xnor2_2 _15927_ (.A(_09020_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__xnor2_2 _15928_ (.A(_09017_),
    .B(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__xnor2_2 _15929_ (.A(_09016_),
    .B(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__a21oi_4 _15930_ (.A1(_08427_),
    .A2(_08428_),
    .B1(_08429_),
    .Y(_09025_));
 sky130_fd_sc_hd__or4_1 _15931_ (.A(_08401_),
    .B(_08402_),
    .C(_08410_),
    .D(_09025_),
    .X(_09026_));
 sky130_fd_sc_hd__a2bb2o_1 _15932_ (.A1_N(_08402_),
    .A2_N(_08411_),
    .B1(_08430_),
    .B2(net7836),
    .X(_09027_));
 sky130_fd_sc_hd__nand2_1 _15933_ (.A(_09026_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__nor2_1 _15934_ (.A(_08417_),
    .B(_08403_),
    .Y(_09029_));
 sky130_fd_sc_hd__xnor2_2 _15935_ (.A(_09028_),
    .B(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__a21boi_2 _15936_ (.A1(net4405),
    .A2(_08128_),
    .B1_N(_08461_),
    .Y(_09031_));
 sky130_fd_sc_hd__nor2_1 _15937_ (.A(_08458_),
    .B(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__o21ai_1 _15938_ (.A1(_08010_),
    .A2(net553),
    .B1(_08017_),
    .Y(_09033_));
 sky130_fd_sc_hd__or3_1 _15939_ (.A(_08010_),
    .B(_08017_),
    .C(_08439_),
    .X(_09034_));
 sky130_fd_sc_hd__a31o_1 _15940_ (.A1(net3453),
    .A2(_09033_),
    .A3(_09034_),
    .B1(_08442_),
    .X(_09035_));
 sky130_fd_sc_hd__or4_4 _15941_ (.A(net8041),
    .B(_06121_),
    .C(_08491_),
    .D(_09035_),
    .X(_09036_));
 sky130_fd_sc_hd__nand2_1 _15942_ (.A(_08450_),
    .B(_08464_),
    .Y(_09037_));
 sky130_fd_sc_hd__xor2_2 _15943_ (.A(_09036_),
    .B(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__xnor2_2 _15944_ (.A(_09032_),
    .B(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__nand2_4 _15945_ (.A(_08181_),
    .B(_08450_),
    .Y(_09040_));
 sky130_fd_sc_hd__o32a_1 _15946_ (.A1(_08444_),
    .A2(net8033),
    .A3(_09040_),
    .B1(_08452_),
    .B2(_08434_),
    .X(_09041_));
 sky130_fd_sc_hd__xor2_2 _15947_ (.A(_09039_),
    .B(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__xnor2_2 _15948_ (.A(_09030_),
    .B(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__nand2_1 _15949_ (.A(_08453_),
    .B(_08468_),
    .Y(_09044_));
 sky130_fd_sc_hd__a21bo_1 _15950_ (.A1(_08420_),
    .A2(_08469_),
    .B1_N(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__xnor2_2 _15951_ (.A(_09043_),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__xnor2_2 _15952_ (.A(_09024_),
    .B(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__and2b_1 _15953_ (.A_N(_08470_),
    .B(_08484_),
    .X(_09048_));
 sky130_fd_sc_hd__a21oi_1 _15954_ (.A1(_08400_),
    .A2(_08485_),
    .B1(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__xor2_1 _15955_ (.A(_09047_),
    .B(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__xnor2_1 _15956_ (.A(_09015_),
    .B(_09050_),
    .Y(_09051_));
 sky130_fd_sc_hd__nor2_1 _15957_ (.A(_08486_),
    .B(_08520_),
    .Y(_09052_));
 sky130_fd_sc_hd__a21oi_1 _15958_ (.A1(_08521_),
    .A2(_08563_),
    .B1(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__nor2_1 _15959_ (.A(_09051_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__nand2_1 _15960_ (.A(_09051_),
    .B(_09053_),
    .Y(_09055_));
 sky130_fd_sc_hd__and2b_1 _15961_ (.A_N(_09054_),
    .B(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__or2b_1 _15962_ (.A(_08561_),
    .B_N(_08541_),
    .X(_09057_));
 sky130_fd_sc_hd__or2b_1 _15963_ (.A(_08562_),
    .B_N(_08540_),
    .X(_09058_));
 sky130_fd_sc_hd__a21o_1 _15964_ (.A1(_08544_),
    .A2(_08549_),
    .B1(_08546_),
    .X(_09059_));
 sky130_fd_sc_hd__nand2_4 _15965_ (.A(net8015),
    .B(_08129_),
    .Y(_09060_));
 sky130_fd_sc_hd__or2_1 _15966_ (.A(_08128_),
    .B(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__clkbuf_4 _15967_ (.A(_09061_),
    .X(_09062_));
 sky130_fd_sc_hd__or2_1 _15968_ (.A(_08127_),
    .B(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__o22a_1 _15969_ (.A1(_08127_),
    .A2(_08614_),
    .B1(_09062_),
    .B2(_08611_),
    .X(_09064_));
 sky130_fd_sc_hd__o21ba_1 _15970_ (.A1(_08615_),
    .A2(_09063_),
    .B1_N(_09064_),
    .X(_09065_));
 sky130_fd_sc_hd__xor2_1 _15971_ (.A(_09059_),
    .B(_09065_),
    .X(_09066_));
 sky130_fd_sc_hd__nand2_1 _15972_ (.A(_08618_),
    .B(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__or2_1 _15973_ (.A(_08618_),
    .B(_09066_),
    .X(_09068_));
 sky130_fd_sc_hd__nand2_1 _15974_ (.A(_09067_),
    .B(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__a21oi_4 _15975_ (.A1(_09057_),
    .A2(_09058_),
    .B1(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__and3_1 _15976_ (.A(_09057_),
    .B(_09058_),
    .C(_09069_),
    .X(_09071_));
 sky130_fd_sc_hd__nor2_1 _15977_ (.A(_09070_),
    .B(_09071_),
    .Y(_09072_));
 sky130_fd_sc_hd__xnor2_2 _15978_ (.A(_09056_),
    .B(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__a21oi_2 _15979_ (.A1(_08607_),
    .A2(_08623_),
    .B1(_08606_),
    .Y(_09074_));
 sky130_fd_sc_hd__xor2_2 _15980_ (.A(_09073_),
    .B(_09074_),
    .X(_09075_));
 sky130_fd_sc_hd__xnor2_1 _15981_ (.A(_08621_),
    .B(_09075_),
    .Y(_09076_));
 sky130_fd_sc_hd__or2b_1 _15982_ (.A(_08624_),
    .B_N(_08654_),
    .X(_09077_));
 sky130_fd_sc_hd__a21boi_2 _15983_ (.A1(_08354_),
    .A2(_08655_),
    .B1_N(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__xor2_1 _15984_ (.A(_09076_),
    .B(_09078_),
    .X(_09079_));
 sky130_fd_sc_hd__and2b_1 _15985_ (.A_N(_08759_),
    .B(_08656_),
    .X(_09080_));
 sky130_fd_sc_hd__nand2_1 _15986_ (.A(_09079_),
    .B(_09080_),
    .Y(_09081_));
 sky130_fd_sc_hd__or2_1 _15987_ (.A(_09079_),
    .B(_09080_),
    .X(_09082_));
 sky130_fd_sc_hd__and2_4 _15988_ (.A(_09081_),
    .B(_09082_),
    .X(_09083_));
 sky130_fd_sc_hd__xor2_4 _15989_ (.A(_08992_),
    .B(_09083_),
    .X(_09084_));
 sky130_fd_sc_hd__mux2_1 _15990_ (.A0(net7768),
    .A1(net5887),
    .S(_08111_),
    .X(_09085_));
 sky130_fd_sc_hd__nand2_1 _15991_ (.A(_09084_),
    .B(net7769),
    .Y(_09086_));
 sky130_fd_sc_hd__or2_1 _15992_ (.A(_09084_),
    .B(net7769),
    .X(_09087_));
 sky130_fd_sc_hd__nand2_1 _15993_ (.A(_09086_),
    .B(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__xor2_4 _15994_ (.A(_08989_),
    .B(_08991_),
    .X(_09089_));
 sky130_fd_sc_hd__mux2_1 _15995_ (.A0(net5859),
    .A1(net7765),
    .S(_08111_),
    .X(_09090_));
 sky130_fd_sc_hd__xor2_4 _15996_ (.A(_08986_),
    .B(_08988_),
    .X(_09091_));
 sky130_fd_sc_hd__mux2_1 _15997_ (.A0(net8220),
    .A1(net8227),
    .S(net4182),
    .X(_09092_));
 sky130_fd_sc_hd__and2_1 _15998_ (.A(_09091_),
    .B(net8542),
    .X(_09093_));
 sky130_fd_sc_hd__xor2_4 _15999_ (.A(_08983_),
    .B(_08985_),
    .X(_09094_));
 sky130_fd_sc_hd__mux2_1 _16000_ (.A0(net5929),
    .A1(net4168),
    .S(_04511_),
    .X(_09095_));
 sky130_fd_sc_hd__o211a_1 _16001_ (.A1(_09091_),
    .A2(net8542),
    .B1(_09094_),
    .C1(net3418),
    .X(_09096_));
 sky130_fd_sc_hd__o22a_1 _16002_ (.A1(_09089_),
    .A2(net7766),
    .B1(_09093_),
    .B2(_09096_),
    .X(_09097_));
 sky130_fd_sc_hd__a21oi_1 _16003_ (.A1(_09089_),
    .A2(net7766),
    .B1(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__or2_1 _16004_ (.A(_09088_),
    .B(_09098_),
    .X(_09099_));
 sky130_fd_sc_hd__nand2_1 _16005_ (.A(_09088_),
    .B(_09098_),
    .Y(_09100_));
 sky130_fd_sc_hd__nand2_1 _16006_ (.A(_09099_),
    .B(_09100_),
    .Y(_09101_));
 sky130_fd_sc_hd__buf_4 _16007_ (.A(_08194_),
    .X(_09102_));
 sky130_fd_sc_hd__clkbuf_4 _16008_ (.A(_09102_),
    .X(_09103_));
 sky130_fd_sc_hd__mux2_1 _16009_ (.A0(_09103_),
    .A1(net7777),
    .S(_08111_),
    .X(_09104_));
 sky130_fd_sc_hd__buf_1 _16010_ (.A(net7778),
    .X(_09105_));
 sky130_fd_sc_hd__nor2_1 _16011_ (.A(_09101_),
    .B(net7779),
    .Y(_09106_));
 sky130_fd_sc_hd__a21o_1 _16012_ (.A1(_09101_),
    .A2(net7779),
    .B1(net3454),
    .X(_09107_));
 sky130_fd_sc_hd__o221a_1 _16013_ (.A1(net4559),
    .A2(_08115_),
    .B1(_09106_),
    .B2(_09107_),
    .C1(_01633_),
    .X(_00466_));
 sky130_fd_sc_hd__a21bo_1 _16014_ (.A1(_08992_),
    .A2(_09083_),
    .B1_N(_09081_),
    .X(_09108_));
 sky130_fd_sc_hd__or2_4 _16015_ (.A(_09076_),
    .B(_09078_),
    .X(_09109_));
 sky130_fd_sc_hd__or2b_1 _16016_ (.A(_09014_),
    .B_N(_08993_),
    .X(_09110_));
 sky130_fd_sc_hd__or3_1 _16017_ (.A(_08529_),
    .B(_08614_),
    .C(_09063_),
    .X(_09111_));
 sky130_fd_sc_hd__o21ai_1 _16018_ (.A1(_08543_),
    .A2(_08614_),
    .B1(_09063_),
    .Y(_09112_));
 sky130_fd_sc_hd__and2_1 _16019_ (.A(_09111_),
    .B(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__nand2_2 _16020_ (.A(net8002),
    .B(_08129_),
    .Y(_09114_));
 sky130_fd_sc_hd__or2_1 _16021_ (.A(_06122_),
    .B(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__clkbuf_4 _16022_ (.A(_09115_),
    .X(_09116_));
 sky130_fd_sc_hd__nor2_1 _16023_ (.A(_08611_),
    .B(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__xnor2_1 _16024_ (.A(_09113_),
    .B(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__and3_1 _16025_ (.A(_08995_),
    .B(_08999_),
    .C(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__a21o_1 _16026_ (.A1(_08995_),
    .A2(_08999_),
    .B1(_09118_),
    .X(_09120_));
 sky130_fd_sc_hd__or2b_2 _16027_ (.A(_09119_),
    .B_N(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__or2_1 _16028_ (.A(_08615_),
    .B(_09063_),
    .X(_09122_));
 sky130_fd_sc_hd__nand2_2 _16029_ (.A(_09059_),
    .B(_09065_),
    .Y(_09123_));
 sky130_fd_sc_hd__nand2_1 _16030_ (.A(_09122_),
    .B(_09123_),
    .Y(_09124_));
 sky130_fd_sc_hd__xor2_1 _16031_ (.A(_09121_),
    .B(_09124_),
    .X(_09125_));
 sky130_fd_sc_hd__a21oi_1 _16032_ (.A1(_09012_),
    .A2(_09110_),
    .B1(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__and3_1 _16033_ (.A(_09012_),
    .B(_09110_),
    .C(_09125_),
    .X(_09127_));
 sky130_fd_sc_hd__nor2_1 _16034_ (.A(_09126_),
    .B(_09127_),
    .Y(_09128_));
 sky130_fd_sc_hd__xnor2_1 _16035_ (.A(_09067_),
    .B(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__a21o_1 _16036_ (.A1(_09001_),
    .A2(_09010_),
    .B1(_09008_),
    .X(_09130_));
 sky130_fd_sc_hd__nand2_1 _16037_ (.A(_09017_),
    .B(_09022_),
    .Y(_09131_));
 sky130_fd_sc_hd__or2b_1 _16038_ (.A(_09023_),
    .B_N(_09016_),
    .X(_09132_));
 sky130_fd_sc_hd__buf_2 _16039_ (.A(_08253_),
    .X(_09133_));
 sky130_fd_sc_hd__or4b_1 _16040_ (.A(_08131_),
    .B(_08142_),
    .C(_08226_),
    .D_N(_09133_),
    .X(_09134_));
 sky130_fd_sc_hd__nor2_2 _16041_ (.A(_06123_),
    .B(net8072),
    .Y(_09135_));
 sky130_fd_sc_hd__a22o_1 _16042_ (.A1(_08996_),
    .A2(_08864_),
    .B1(_09133_),
    .B2(_09135_),
    .X(_09136_));
 sky130_fd_sc_hd__nand2_1 _16043_ (.A(_09134_),
    .B(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__nor2_1 _16044_ (.A(_08542_),
    .B(_08616_),
    .Y(_09138_));
 sky130_fd_sc_hd__xnor2_2 _16045_ (.A(_09137_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__or4_1 _16046_ (.A(_08389_),
    .B(_08211_),
    .C(_08294_),
    .D(_08306_),
    .X(_09140_));
 sky130_fd_sc_hd__o22ai_1 _16047_ (.A1(_08389_),
    .A2(_08308_),
    .B1(_08309_),
    .B2(_08211_),
    .Y(_09141_));
 sky130_fd_sc_hd__nand2_1 _16048_ (.A(_09140_),
    .B(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__or2_1 _16049_ (.A(_08207_),
    .B(_08323_),
    .X(_09143_));
 sky130_fd_sc_hd__xnor2_1 _16050_ (.A(_09142_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__o31a_1 _16051_ (.A1(_08229_),
    .A2(_08323_),
    .A3(_09004_),
    .B1(_09002_),
    .X(_09145_));
 sky130_fd_sc_hd__nor2_1 _16052_ (.A(_09144_),
    .B(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__and2_1 _16053_ (.A(_09144_),
    .B(_09145_),
    .X(_09147_));
 sky130_fd_sc_hd__nor2_1 _16054_ (.A(_09146_),
    .B(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__xnor2_1 _16055_ (.A(_09139_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__a21o_1 _16056_ (.A1(_09131_),
    .A2(_09132_),
    .B1(_09149_),
    .X(_09150_));
 sky130_fd_sc_hd__nand3_1 _16057_ (.A(_09131_),
    .B(_09132_),
    .C(_09149_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_1 _16058_ (.A(_09150_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__xnor2_1 _16059_ (.A(_09130_),
    .B(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__a21bo_1 _16060_ (.A1(_09019_),
    .A2(_09021_),
    .B1_N(_09018_),
    .X(_09154_));
 sky130_fd_sc_hd__a21bo_1 _16061_ (.A1(_09027_),
    .A2(_09029_),
    .B1_N(_09026_),
    .X(_09155_));
 sky130_fd_sc_hd__or4_1 _16062_ (.A(_08880_),
    .B(_08391_),
    .C(_08403_),
    .D(_08418_),
    .X(_09156_));
 sky130_fd_sc_hd__a22o_1 _16063_ (.A1(_08244_),
    .A2(_08414_),
    .B1(_08386_),
    .B2(_08246_),
    .X(_09157_));
 sky130_fd_sc_hd__nand2_1 _16064_ (.A(_09156_),
    .B(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__nor2_1 _16065_ (.A(_08509_),
    .B(_08392_),
    .Y(_09159_));
 sky130_fd_sc_hd__xnor2_1 _16066_ (.A(_09158_),
    .B(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__xnor2_1 _16067_ (.A(_09155_),
    .B(_09160_),
    .Y(_09161_));
 sky130_fd_sc_hd__xnor2_1 _16068_ (.A(_09154_),
    .B(_09161_),
    .Y(_09162_));
 sky130_fd_sc_hd__nor2_1 _16069_ (.A(_08417_),
    .B(_08411_),
    .Y(_09163_));
 sky130_fd_sc_hd__or4_1 _16070_ (.A(_08401_),
    .B(_08402_),
    .C(_09025_),
    .D(_09031_),
    .X(_09164_));
 sky130_fd_sc_hd__buf_2 _16071_ (.A(_09031_),
    .X(_09165_));
 sky130_fd_sc_hd__a2bb2o_1 _16072_ (.A1_N(_08401_),
    .A2_N(_09165_),
    .B1(_08180_),
    .B2(_08430_),
    .X(_09166_));
 sky130_fd_sc_hd__and2_1 _16073_ (.A(_09164_),
    .B(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__xor2_2 _16074_ (.A(_09163_),
    .B(_09167_),
    .X(_09168_));
 sky130_fd_sc_hd__and2_1 _16075_ (.A(net3726),
    .B(_08128_),
    .X(_09169_));
 sky130_fd_sc_hd__a21oi_4 _16076_ (.A1(_08181_),
    .A2(_08450_),
    .B1(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__nor2_1 _16077_ (.A(_08458_),
    .B(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__nor4_4 _16078_ (.A(_08010_),
    .B(_08017_),
    .C(_08021_),
    .D(_08439_),
    .Y(_09172_));
 sky130_fd_sc_hd__o31a_1 _16079_ (.A1(_08010_),
    .A2(_08017_),
    .A3(net565),
    .B1(_08021_),
    .X(_09173_));
 sky130_fd_sc_hd__o31ai_4 _16080_ (.A1(_08114_),
    .A2(_09172_),
    .A3(_09173_),
    .B1(_08441_),
    .Y(_09174_));
 sky130_fd_sc_hd__or4_1 _16081_ (.A(net8041),
    .B(_08128_),
    .C(_08491_),
    .D(_09174_),
    .X(_09175_));
 sky130_fd_sc_hd__or4_1 _16082_ (.A(net8065),
    .B(_08128_),
    .C(_08491_),
    .D(_09035_),
    .X(_09176_));
 sky130_fd_sc_hd__or4_4 _16083_ (.A(net8065),
    .B(_08128_),
    .C(_08491_),
    .D(_09174_),
    .X(_09177_));
 sky130_fd_sc_hd__o2bb2a_2 _16084_ (.A1_N(_09175_),
    .A2_N(_09176_),
    .B1(_09036_),
    .B2(_09177_),
    .X(_09178_));
 sky130_fd_sc_hd__xnor2_2 _16085_ (.A(_09171_),
    .B(_09178_),
    .Y(_09179_));
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(net3551),
    .B(_08491_),
    .Y(_09180_));
 sky130_fd_sc_hd__a21o_2 _16087_ (.A1(_09180_),
    .A2(_09035_),
    .B1(_08128_),
    .X(_09181_));
 sky130_fd_sc_hd__nor2_1 _16088_ (.A(net8033),
    .B(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__a32o_1 _16089_ (.A1(_08450_),
    .A2(_08464_),
    .A3(_09182_),
    .B1(_09038_),
    .B2(_09032_),
    .X(_09183_));
 sky130_fd_sc_hd__xnor2_2 _16090_ (.A(_09179_),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__xnor2_2 _16091_ (.A(_09168_),
    .B(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__nor2_1 _16092_ (.A(_09039_),
    .B(_09041_),
    .Y(_09186_));
 sky130_fd_sc_hd__a21oi_2 _16093_ (.A1(_09030_),
    .A2(_09042_),
    .B1(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__xor2_2 _16094_ (.A(_09185_),
    .B(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__xnor2_1 _16095_ (.A(_09162_),
    .B(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__and2b_1 _16096_ (.A_N(_09043_),
    .B(_09045_),
    .X(_09190_));
 sky130_fd_sc_hd__a21oi_1 _16097_ (.A1(_09024_),
    .A2(_09046_),
    .B1(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__nor2_1 _16098_ (.A(_09189_),
    .B(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__nand2_1 _16099_ (.A(_09189_),
    .B(_09191_),
    .Y(_09193_));
 sky130_fd_sc_hd__and2b_1 _16100_ (.A_N(_09192_),
    .B(_09193_),
    .X(_09194_));
 sky130_fd_sc_hd__xnor2_2 _16101_ (.A(_09153_),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__nor2_1 _16102_ (.A(_09047_),
    .B(_09049_),
    .Y(_09196_));
 sky130_fd_sc_hd__a21oi_1 _16103_ (.A1(_09015_),
    .A2(_09050_),
    .B1(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__xor2_1 _16104_ (.A(_09195_),
    .B(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__xnor2_1 _16105_ (.A(_09129_),
    .B(_09198_),
    .Y(_09199_));
 sky130_fd_sc_hd__a21oi_1 _16106_ (.A1(_09055_),
    .A2(_09072_),
    .B1(_09054_),
    .Y(_09200_));
 sky130_fd_sc_hd__nor2_1 _16107_ (.A(_09199_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__nand2_1 _16108_ (.A(_09199_),
    .B(_09200_),
    .Y(_09202_));
 sky130_fd_sc_hd__and2b_1 _16109_ (.A_N(_09201_),
    .B(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__xnor2_4 _16110_ (.A(_09070_),
    .B(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__nor2_1 _16111_ (.A(_09073_),
    .B(_09074_),
    .Y(_09205_));
 sky130_fd_sc_hd__a21oi_2 _16112_ (.A1(_08621_),
    .A2(_09075_),
    .B1(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__xnor2_4 _16113_ (.A(_09204_),
    .B(_09206_),
    .Y(_09207_));
 sky130_fd_sc_hd__xor2_4 _16114_ (.A(_09109_),
    .B(_09207_),
    .X(_09208_));
 sky130_fd_sc_hd__xor2_4 _16115_ (.A(_09108_),
    .B(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__mux2_1 _16116_ (.A0(net8216),
    .A1(net5904),
    .S(_08111_),
    .X(_09210_));
 sky130_fd_sc_hd__xnor2_1 _16117_ (.A(_09209_),
    .B(net3420),
    .Y(_09211_));
 sky130_fd_sc_hd__a21oi_2 _16118_ (.A1(_09086_),
    .A2(_09099_),
    .B1(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__and3_1 _16119_ (.A(_09086_),
    .B(_09099_),
    .C(_09211_),
    .X(_09213_));
 sky130_fd_sc_hd__or3_1 _16120_ (.A(net7779),
    .B(_09212_),
    .C(_09213_),
    .X(_09214_));
 sky130_fd_sc_hd__o21ai_1 _16121_ (.A1(_09212_),
    .A2(_09213_),
    .B1(net7779),
    .Y(_09215_));
 sky130_fd_sc_hd__o21ai_1 _16122_ (.A1(net4612),
    .A2(_08115_),
    .B1(_08038_),
    .Y(_09216_));
 sky130_fd_sc_hd__a31oi_1 _16123_ (.A1(_08115_),
    .A2(_09214_),
    .A3(_09215_),
    .B1(net4613),
    .Y(_00467_));
 sky130_fd_sc_hd__nor2_1 _16124_ (.A(_09204_),
    .B(_09206_),
    .Y(_09217_));
 sky130_fd_sc_hd__a31o_1 _16125_ (.A1(_08618_),
    .A2(_09066_),
    .A3(_09128_),
    .B1(_09126_),
    .X(_09218_));
 sky130_fd_sc_hd__or2_1 _16126_ (.A(_09195_),
    .B(_09197_),
    .X(_09219_));
 sky130_fd_sc_hd__nand2_1 _16127_ (.A(_09129_),
    .B(_09198_),
    .Y(_09220_));
 sky130_fd_sc_hd__or2b_1 _16128_ (.A(_09152_),
    .B_N(_09130_),
    .X(_09221_));
 sky130_fd_sc_hd__nand2_1 _16129_ (.A(_09150_),
    .B(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand2_1 _16130_ (.A(net8068),
    .B(_08129_),
    .Y(_09223_));
 sky130_fd_sc_hd__or2_1 _16131_ (.A(_06124_),
    .B(net4908),
    .X(_09224_));
 sky130_fd_sc_hd__clkbuf_4 _16132_ (.A(_09224_),
    .X(_09225_));
 sky130_fd_sc_hd__or2_2 _16133_ (.A(_08611_),
    .B(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__a21bo_1 _16134_ (.A1(_09112_),
    .A2(_09117_),
    .B1_N(_09111_),
    .X(_09227_));
 sky130_fd_sc_hd__inv_2 _16135_ (.A(_09227_),
    .Y(_09228_));
 sky130_fd_sc_hd__or3_1 _16136_ (.A(_08542_),
    .B(_08616_),
    .C(_09137_),
    .X(_09229_));
 sky130_fd_sc_hd__or2_1 _16137_ (.A(_08277_),
    .B(_08614_),
    .X(_09230_));
 sky130_fd_sc_hd__o21ai_1 _16138_ (.A1(_08529_),
    .A2(_09062_),
    .B1(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__or3_1 _16139_ (.A(_08529_),
    .B(_09062_),
    .C(_09230_),
    .X(_09232_));
 sky130_fd_sc_hd__and2_1 _16140_ (.A(_09231_),
    .B(_09232_),
    .X(_09233_));
 sky130_fd_sc_hd__nor2_1 _16141_ (.A(_08127_),
    .B(_09116_),
    .Y(_09234_));
 sky130_fd_sc_hd__xnor2_1 _16142_ (.A(_09233_),
    .B(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__a21o_1 _16143_ (.A1(_09134_),
    .A2(_09229_),
    .B1(_09235_),
    .X(_09236_));
 sky130_fd_sc_hd__nand3_1 _16144_ (.A(_09134_),
    .B(_09229_),
    .C(_09235_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_1 _16145_ (.A(_09236_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__xnor2_2 _16146_ (.A(_09228_),
    .B(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__a21o_1 _16147_ (.A1(_09122_),
    .A2(_09120_),
    .B1(_09119_),
    .X(_09240_));
 sky130_fd_sc_hd__xor2_2 _16148_ (.A(_09239_),
    .B(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__xor2_2 _16149_ (.A(_09226_),
    .B(_09241_),
    .X(_09242_));
 sky130_fd_sc_hd__xor2_2 _16150_ (.A(_09222_),
    .B(_09242_),
    .X(_09243_));
 sky130_fd_sc_hd__nor2_1 _16151_ (.A(_09123_),
    .B(_09121_),
    .Y(_09244_));
 sky130_fd_sc_hd__xnor2_1 _16152_ (.A(_09243_),
    .B(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__a21o_1 _16153_ (.A1(_09139_),
    .A2(_09148_),
    .B1(_09146_),
    .X(_09246_));
 sky130_fd_sc_hd__or2b_1 _16154_ (.A(_09161_),
    .B_N(_09154_),
    .X(_09247_));
 sky130_fd_sc_hd__a21bo_1 _16155_ (.A1(_09155_),
    .A2(_09160_),
    .B1_N(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__buf_2 _16156_ (.A(_08204_),
    .X(_09249_));
 sky130_fd_sc_hd__and3_1 _16157_ (.A(_08996_),
    .B(_09135_),
    .C(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__nand2_1 _16158_ (.A(_08864_),
    .B(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__a22o_1 _16159_ (.A1(_08996_),
    .A2(_09249_),
    .B1(_08864_),
    .B2(_09135_),
    .X(_09252_));
 sky130_fd_sc_hd__nand2_1 _16160_ (.A(_09251_),
    .B(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__inv_2 _16161_ (.A(_08535_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand2_1 _16162_ (.A(_09133_),
    .B(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__or2_1 _16163_ (.A(_09253_),
    .B(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__nand2_1 _16164_ (.A(_09253_),
    .B(_09255_),
    .Y(_09257_));
 sky130_fd_sc_hd__and2_1 _16165_ (.A(_09256_),
    .B(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__or4_1 _16166_ (.A(_08389_),
    .B(_08308_),
    .C(_08309_),
    .D(_08392_),
    .X(_09259_));
 sky130_fd_sc_hd__o22ai_1 _16167_ (.A1(_08389_),
    .A2(_08309_),
    .B1(_08392_),
    .B2(_08308_),
    .Y(_09260_));
 sky130_fd_sc_hd__nand2_1 _16168_ (.A(_09259_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__clkbuf_4 _16169_ (.A(_08323_),
    .X(_09262_));
 sky130_fd_sc_hd__nor2_1 _16170_ (.A(_08211_),
    .B(_09262_),
    .Y(_09263_));
 sky130_fd_sc_hd__xor2_1 _16171_ (.A(_09261_),
    .B(_09263_),
    .X(_09264_));
 sky130_fd_sc_hd__o31a_1 _16172_ (.A1(_08207_),
    .A2(_09262_),
    .A3(_09142_),
    .B1(_09140_),
    .X(_09265_));
 sky130_fd_sc_hd__nor2_1 _16173_ (.A(_09264_),
    .B(_09265_),
    .Y(_09266_));
 sky130_fd_sc_hd__and2_1 _16174_ (.A(_09264_),
    .B(_09265_),
    .X(_09267_));
 sky130_fd_sc_hd__nor2_1 _16175_ (.A(_09266_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__xor2_2 _16176_ (.A(_09258_),
    .B(_09268_),
    .X(_09269_));
 sky130_fd_sc_hd__xnor2_2 _16177_ (.A(_09248_),
    .B(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__xnor2_2 _16178_ (.A(_09246_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__clkbuf_4 _16179_ (.A(_08509_),
    .X(_09272_));
 sky130_fd_sc_hd__or3_1 _16180_ (.A(_09272_),
    .B(_08392_),
    .C(_09158_),
    .X(_09273_));
 sky130_fd_sc_hd__a21boi_2 _16181_ (.A1(_09163_),
    .A2(_09166_),
    .B1_N(_09164_),
    .Y(_09274_));
 sky130_fd_sc_hd__or2_1 _16182_ (.A(_08241_),
    .B(_08403_),
    .X(_09275_));
 sky130_fd_sc_hd__nor2_1 _16183_ (.A(_08221_),
    .B(_08411_),
    .Y(_09276_));
 sky130_fd_sc_hd__xnor2_1 _16184_ (.A(_09275_),
    .B(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_08509_),
    .B(_08418_),
    .Y(_09278_));
 sky130_fd_sc_hd__and2_1 _16186_ (.A(_09277_),
    .B(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__nor2_1 _16187_ (.A(_09277_),
    .B(_09278_),
    .Y(_09280_));
 sky130_fd_sc_hd__or2_1 _16188_ (.A(_09279_),
    .B(_09280_),
    .X(_09281_));
 sky130_fd_sc_hd__xnor2_1 _16189_ (.A(_09274_),
    .B(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__a21o_1 _16190_ (.A1(_09156_),
    .A2(_09273_),
    .B1(_09282_),
    .X(_09283_));
 sky130_fd_sc_hd__nand3_1 _16191_ (.A(_09156_),
    .B(_09273_),
    .C(_09282_),
    .Y(_09284_));
 sky130_fd_sc_hd__and2_1 _16192_ (.A(_09283_),
    .B(_09284_),
    .X(_09285_));
 sky130_fd_sc_hd__nand2_1 _16193_ (.A(_08666_),
    .B(_08430_),
    .Y(_09286_));
 sky130_fd_sc_hd__or4_1 _16194_ (.A(_08401_),
    .B(_08402_),
    .C(_09165_),
    .D(_09170_),
    .X(_09287_));
 sky130_fd_sc_hd__a21o_1 _16195_ (.A1(_08181_),
    .A2(_08450_),
    .B1(_09169_),
    .X(_09288_));
 sky130_fd_sc_hd__a2bb2o_1 _16196_ (.A1_N(_08402_),
    .A2_N(_09165_),
    .B1(_09288_),
    .B2(net7836),
    .X(_09289_));
 sky130_fd_sc_hd__nand2_1 _16197_ (.A(_09287_),
    .B(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__xor2_2 _16198_ (.A(_09286_),
    .B(_09290_),
    .X(_09291_));
 sky130_fd_sc_hd__a21boi_4 _16199_ (.A1(net3841),
    .A2(_06122_),
    .B1_N(_09181_),
    .Y(_09292_));
 sky130_fd_sc_hd__nor2_1 _16200_ (.A(_08905_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__or2_1 _16201_ (.A(_08024_),
    .B(net75),
    .X(_09294_));
 sky130_fd_sc_hd__nand2_1 _16202_ (.A(_08024_),
    .B(net75),
    .Y(_09295_));
 sky130_fd_sc_hd__a31o_1 _16203_ (.A1(_08421_),
    .A2(_09294_),
    .A3(_09295_),
    .B1(_08442_),
    .X(_09296_));
 sky130_fd_sc_hd__or4_2 _16204_ (.A(net8041),
    .B(_06122_),
    .C(_08491_),
    .D(_09296_),
    .X(_09297_));
 sky130_fd_sc_hd__xor2_2 _16205_ (.A(_09177_),
    .B(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__xor2_2 _16206_ (.A(_09293_),
    .B(_09298_),
    .X(_09299_));
 sky130_fd_sc_hd__nand2_1 _16207_ (.A(_09171_),
    .B(_09178_),
    .Y(_09300_));
 sky130_fd_sc_hd__o21a_1 _16208_ (.A1(_09036_),
    .A2(_09177_),
    .B1(_09300_),
    .X(_09301_));
 sky130_fd_sc_hd__xnor2_2 _16209_ (.A(_09299_),
    .B(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__xnor2_2 _16210_ (.A(_09291_),
    .B(_09302_),
    .Y(_09303_));
 sky130_fd_sc_hd__or2_1 _16211_ (.A(_09171_),
    .B(_09178_),
    .X(_09304_));
 sky130_fd_sc_hd__a32o_1 _16212_ (.A1(_09300_),
    .A2(_09304_),
    .A3(_09183_),
    .B1(_09184_),
    .B2(_09168_),
    .X(_09305_));
 sky130_fd_sc_hd__xnor2_2 _16213_ (.A(_09303_),
    .B(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__xnor2_2 _16214_ (.A(_09285_),
    .B(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__nor2_1 _16215_ (.A(_09185_),
    .B(_09187_),
    .Y(_09308_));
 sky130_fd_sc_hd__a21oi_2 _16216_ (.A1(_09162_),
    .A2(_09188_),
    .B1(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__xor2_2 _16217_ (.A(_09307_),
    .B(_09309_),
    .X(_09310_));
 sky130_fd_sc_hd__xnor2_2 _16218_ (.A(_09271_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__a21oi_2 _16219_ (.A1(_09153_),
    .A2(_09193_),
    .B1(_09192_),
    .Y(_09312_));
 sky130_fd_sc_hd__xor2_1 _16220_ (.A(_09311_),
    .B(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__xnor2_1 _16221_ (.A(_09245_),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__a21oi_2 _16222_ (.A1(_09219_),
    .A2(_09220_),
    .B1(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__and3_1 _16223_ (.A(_09219_),
    .B(_09220_),
    .C(_09314_),
    .X(_09316_));
 sky130_fd_sc_hd__nor2_1 _16224_ (.A(_09315_),
    .B(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__xnor2_1 _16225_ (.A(_09218_),
    .B(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__a21oi_1 _16226_ (.A1(_09070_),
    .A2(_09202_),
    .B1(_09201_),
    .Y(_09319_));
 sky130_fd_sc_hd__xor2_1 _16227_ (.A(_09318_),
    .B(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__nand2_2 _16228_ (.A(_09217_),
    .B(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__or2_1 _16229_ (.A(_09217_),
    .B(_09320_),
    .X(_09322_));
 sky130_fd_sc_hd__nand2_4 _16230_ (.A(_09321_),
    .B(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__a21oi_1 _16231_ (.A1(_09109_),
    .A2(_09081_),
    .B1(_09207_),
    .Y(_09324_));
 sky130_fd_sc_hd__a31oi_4 _16232_ (.A1(_08992_),
    .A2(_09083_),
    .A3(_09208_),
    .B1(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__xor2_4 _16233_ (.A(_09323_),
    .B(_09325_),
    .X(_09326_));
 sky130_fd_sc_hd__mux2_1 _16234_ (.A0(net7781),
    .A1(net5768),
    .S(_08111_),
    .X(_09327_));
 sky130_fd_sc_hd__nand2_1 _16235_ (.A(_09326_),
    .B(net5769),
    .Y(_09328_));
 sky130_fd_sc_hd__or2_1 _16236_ (.A(_09326_),
    .B(net5769),
    .X(_09329_));
 sky130_fd_sc_hd__nand2_1 _16237_ (.A(_09328_),
    .B(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__a21oi_2 _16238_ (.A1(_09209_),
    .A2(net3420),
    .B1(_09212_),
    .Y(_09331_));
 sky130_fd_sc_hd__xnor2_1 _16239_ (.A(_09330_),
    .B(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__nor2_1 _16240_ (.A(net7779),
    .B(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__a21o_1 _16241_ (.A1(net7779),
    .A2(_09332_),
    .B1(net3454),
    .X(_09334_));
 sky130_fd_sc_hd__o221a_1 _16242_ (.A1(net4640),
    .A2(_08115_),
    .B1(_09333_),
    .B2(_09334_),
    .C1(_01633_),
    .X(_00468_));
 sky130_fd_sc_hd__o21ai_4 _16243_ (.A1(_09323_),
    .A2(_09325_),
    .B1(_09321_),
    .Y(_09335_));
 sky130_fd_sc_hd__or2_2 _16244_ (.A(_09318_),
    .B(_09319_),
    .X(_09336_));
 sky130_fd_sc_hd__a21o_1 _16245_ (.A1(_09150_),
    .A2(_09221_),
    .B1(_09242_),
    .X(_09337_));
 sky130_fd_sc_hd__o31ai_4 _16246_ (.A1(_09123_),
    .A2(_09121_),
    .A3(_09243_),
    .B1(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__or2b_1 _16247_ (.A(_09226_),
    .B_N(_09241_),
    .X(_09339_));
 sky130_fd_sc_hd__o21ai_2 _16248_ (.A1(_09239_),
    .A2(_09240_),
    .B1(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__or2b_1 _16249_ (.A(_09270_),
    .B_N(_09246_),
    .X(_09341_));
 sky130_fd_sc_hd__a21bo_1 _16250_ (.A1(_09248_),
    .A2(_09269_),
    .B1_N(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__nand2_1 _16251_ (.A(net8275),
    .B(_08129_),
    .Y(_09343_));
 sky130_fd_sc_hd__or2_1 _16252_ (.A(_06123_),
    .B(net4913),
    .X(_09344_));
 sky130_fd_sc_hd__buf_4 _16253_ (.A(_09344_),
    .X(_09345_));
 sky130_fd_sc_hd__o22a_1 _16254_ (.A1(_08127_),
    .A2(_09225_),
    .B1(_09345_),
    .B2(_08611_),
    .X(_09346_));
 sky130_fd_sc_hd__or2_1 _16255_ (.A(_08127_),
    .B(_09345_),
    .X(_09347_));
 sky130_fd_sc_hd__nor2_1 _16256_ (.A(_09226_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__nor2_1 _16257_ (.A(_09346_),
    .B(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__a21bo_1 _16258_ (.A1(_09231_),
    .A2(_09234_),
    .B1_N(_09232_),
    .X(_09350_));
 sky130_fd_sc_hd__nor2_2 _16259_ (.A(_06122_),
    .B(_08612_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand2_1 _16260_ (.A(_09133_),
    .B(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__or2_1 _16261_ (.A(_08542_),
    .B(_09062_),
    .X(_09353_));
 sky130_fd_sc_hd__nor2_2 _16262_ (.A(_06122_),
    .B(_09060_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_1 _16263_ (.A(_09133_),
    .B(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__nor2_1 _16264_ (.A(_09230_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__a21oi_1 _16265_ (.A1(_09352_),
    .A2(_09353_),
    .B1(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__nor2_1 _16266_ (.A(_08543_),
    .B(_09116_),
    .Y(_09358_));
 sky130_fd_sc_hd__xnor2_1 _16267_ (.A(_09357_),
    .B(_09358_),
    .Y(_09359_));
 sky130_fd_sc_hd__a21oi_1 _16268_ (.A1(_09251_),
    .A2(_09256_),
    .B1(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__and3_1 _16269_ (.A(_09251_),
    .B(_09256_),
    .C(_09359_),
    .X(_09361_));
 sky130_fd_sc_hd__nor2_1 _16270_ (.A(_09360_),
    .B(_09361_),
    .Y(_09362_));
 sky130_fd_sc_hd__xnor2_1 _16271_ (.A(_09350_),
    .B(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__o21a_1 _16272_ (.A1(_09228_),
    .A2(_09238_),
    .B1(_09236_),
    .X(_09364_));
 sky130_fd_sc_hd__nor2_1 _16273_ (.A(_09363_),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__and2_1 _16274_ (.A(_09363_),
    .B(_09364_),
    .X(_09366_));
 sky130_fd_sc_hd__nor2_1 _16275_ (.A(_09365_),
    .B(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__xor2_2 _16276_ (.A(_09349_),
    .B(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__xnor2_2 _16277_ (.A(_09342_),
    .B(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__xnor2_2 _16278_ (.A(_09340_),
    .B(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__a21o_1 _16279_ (.A1(_09258_),
    .A2(_09268_),
    .B1(_09266_),
    .X(_09371_));
 sky130_fd_sc_hd__o21ai_2 _16280_ (.A1(_09274_),
    .A2(_09281_),
    .B1(_09283_),
    .Y(_09372_));
 sky130_fd_sc_hd__buf_2 _16281_ (.A(_08185_),
    .X(_09373_));
 sky130_fd_sc_hd__nand2_1 _16282_ (.A(_08996_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__nand2_1 _16283_ (.A(_09135_),
    .B(_09249_),
    .Y(_09375_));
 sky130_fd_sc_hd__and2_1 _16284_ (.A(_09373_),
    .B(_09250_),
    .X(_09376_));
 sky130_fd_sc_hd__a21o_1 _16285_ (.A1(_09374_),
    .A2(_09375_),
    .B1(_09376_),
    .X(_09377_));
 sky130_fd_sc_hd__nor2_1 _16286_ (.A(_08226_),
    .B(_08535_),
    .Y(_09378_));
 sky130_fd_sc_hd__xnor2_2 _16287_ (.A(_09377_),
    .B(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__or2_1 _16288_ (.A(_08306_),
    .B(_08392_),
    .X(_09380_));
 sky130_fd_sc_hd__or3_1 _16289_ (.A(_08308_),
    .B(_08418_),
    .C(_09380_),
    .X(_09381_));
 sky130_fd_sc_hd__o21ai_1 _16290_ (.A1(_08308_),
    .A2(_08418_),
    .B1(_09380_),
    .Y(_09382_));
 sky130_fd_sc_hd__and2_1 _16291_ (.A(_09381_),
    .B(_09382_),
    .X(_09383_));
 sky130_fd_sc_hd__nor2_1 _16292_ (.A(_08389_),
    .B(_09262_),
    .Y(_09384_));
 sky130_fd_sc_hd__xnor2_2 _16293_ (.A(_09383_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__a21bo_1 _16294_ (.A1(_09260_),
    .A2(_09263_),
    .B1_N(_09259_),
    .X(_09386_));
 sky130_fd_sc_hd__xnor2_2 _16295_ (.A(_09385_),
    .B(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__xor2_2 _16296_ (.A(_09379_),
    .B(_09387_),
    .X(_09388_));
 sky130_fd_sc_hd__xnor2_2 _16297_ (.A(_09372_),
    .B(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__xnor2_2 _16298_ (.A(_09371_),
    .B(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__a31o_1 _16299_ (.A1(_08246_),
    .A2(_08414_),
    .A3(_09276_),
    .B1(_09279_),
    .X(_09391_));
 sky130_fd_sc_hd__nor2_1 _16300_ (.A(_08391_),
    .B(_08411_),
    .Y(_09392_));
 sky130_fd_sc_hd__nand2_1 _16301_ (.A(_08244_),
    .B(_08430_),
    .Y(_09393_));
 sky130_fd_sc_hd__xnor2_1 _16302_ (.A(_09392_),
    .B(_09393_),
    .Y(_09394_));
 sky130_fd_sc_hd__nor2_1 _16303_ (.A(_08509_),
    .B(_08403_),
    .Y(_09395_));
 sky130_fd_sc_hd__xnor2_1 _16304_ (.A(_09394_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__o21ai_1 _16305_ (.A1(_09286_),
    .A2(_09290_),
    .B1(_09287_),
    .Y(_09397_));
 sky130_fd_sc_hd__or2b_1 _16306_ (.A(_09396_),
    .B_N(_09397_),
    .X(_09398_));
 sky130_fd_sc_hd__or2b_1 _16307_ (.A(_09397_),
    .B_N(_09396_),
    .X(_09399_));
 sky130_fd_sc_hd__nand2_1 _16308_ (.A(_09398_),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__xnor2_1 _16309_ (.A(_09391_),
    .B(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__nor2_1 _16310_ (.A(_08417_),
    .B(_09165_),
    .Y(_09402_));
 sky130_fd_sc_hd__clkbuf_4 _16311_ (.A(_09292_),
    .X(_09403_));
 sky130_fd_sc_hd__nand2_1 _16312_ (.A(_08180_),
    .B(_09288_),
    .Y(_09404_));
 sky130_fd_sc_hd__nor3_1 _16313_ (.A(_08948_),
    .B(_09403_),
    .C(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__o21ai_1 _16314_ (.A1(_08948_),
    .A2(_09292_),
    .B1(_09404_),
    .Y(_09406_));
 sky130_fd_sc_hd__and2b_1 _16315_ (.A_N(_09405_),
    .B(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__xor2_1 _16316_ (.A(_09402_),
    .B(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__nand2_1 _16317_ (.A(net3542),
    .B(_08491_),
    .Y(_09409_));
 sky130_fd_sc_hd__a21o_2 _16318_ (.A1(_09409_),
    .A2(_09174_),
    .B1(_06122_),
    .X(_09410_));
 sky130_fd_sc_hd__a21boi_4 _16319_ (.A1(net4624),
    .A2(_06123_),
    .B1_N(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__nor2_1 _16320_ (.A(_08905_),
    .B(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__clkbuf_4 _16321_ (.A(_08491_),
    .X(_09413_));
 sky130_fd_sc_hd__a221oi_2 _16322_ (.A1(_07989_),
    .A2(_07979_),
    .B1(_08027_),
    .B2(_08020_),
    .C1(_07869_),
    .Y(_09414_));
 sky130_fd_sc_hd__a21oi_1 _16323_ (.A1(_08024_),
    .A2(net75),
    .B1(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__a31o_1 _16324_ (.A1(_08024_),
    .A2(_09414_),
    .A3(net75),
    .B1(_08115_),
    .X(_09416_));
 sky130_fd_sc_hd__o21ai_4 _16325_ (.A1(_09415_),
    .A2(_09416_),
    .B1(_08441_),
    .Y(_09417_));
 sky130_fd_sc_hd__or4_1 _16326_ (.A(net8041),
    .B(_06122_),
    .C(_09413_),
    .D(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__nand2_1 _16327_ (.A(net4537),
    .B(_08491_),
    .Y(_09419_));
 sky130_fd_sc_hd__a21oi_1 _16328_ (.A1(_09419_),
    .A2(_09296_),
    .B1(_08474_),
    .Y(_09420_));
 sky130_fd_sc_hd__xnor2_1 _16329_ (.A(_09418_),
    .B(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__xnor2_1 _16330_ (.A(_09412_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__nor2_1 _16331_ (.A(_09177_),
    .B(_09297_),
    .Y(_09423_));
 sky130_fd_sc_hd__a21o_1 _16332_ (.A1(_09293_),
    .A2(_09298_),
    .B1(_09423_),
    .X(_09424_));
 sky130_fd_sc_hd__xnor2_1 _16333_ (.A(_09422_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__xnor2_1 _16334_ (.A(_09408_),
    .B(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__or2b_1 _16335_ (.A(_09301_),
    .B_N(_09299_),
    .X(_09427_));
 sky130_fd_sc_hd__a21bo_1 _16336_ (.A1(_09291_),
    .A2(_09302_),
    .B1_N(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__xnor2_1 _16337_ (.A(_09426_),
    .B(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__xnor2_1 _16338_ (.A(_09401_),
    .B(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__and2b_1 _16339_ (.A_N(_09303_),
    .B(_09305_),
    .X(_09431_));
 sky130_fd_sc_hd__a21oi_1 _16340_ (.A1(_09285_),
    .A2(_09306_),
    .B1(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__nor2_1 _16341_ (.A(_09430_),
    .B(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__nand2_1 _16342_ (.A(_09430_),
    .B(_09432_),
    .Y(_09434_));
 sky130_fd_sc_hd__and2b_1 _16343_ (.A_N(_09433_),
    .B(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__xnor2_2 _16344_ (.A(_09390_),
    .B(_09435_),
    .Y(_09436_));
 sky130_fd_sc_hd__nor2_1 _16345_ (.A(_09307_),
    .B(_09309_),
    .Y(_09437_));
 sky130_fd_sc_hd__a21oi_2 _16346_ (.A1(_09271_),
    .A2(_09310_),
    .B1(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__xor2_2 _16347_ (.A(_09436_),
    .B(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__xnor2_1 _16348_ (.A(_09370_),
    .B(_09439_),
    .Y(_09440_));
 sky130_fd_sc_hd__nor2_1 _16349_ (.A(_09311_),
    .B(_09312_),
    .Y(_09441_));
 sky130_fd_sc_hd__a21oi_1 _16350_ (.A1(_09245_),
    .A2(_09313_),
    .B1(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__nor2_1 _16351_ (.A(_09440_),
    .B(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__nand2_1 _16352_ (.A(_09440_),
    .B(_09442_),
    .Y(_09444_));
 sky130_fd_sc_hd__and2b_1 _16353_ (.A_N(_09443_),
    .B(_09444_),
    .X(_09445_));
 sky130_fd_sc_hd__xnor2_4 _16354_ (.A(_09338_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__a21oi_4 _16355_ (.A1(_09218_),
    .A2(_09317_),
    .B1(_09315_),
    .Y(_09447_));
 sky130_fd_sc_hd__xnor2_4 _16356_ (.A(_09446_),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__xnor2_4 _16357_ (.A(_09336_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__xnor2_4 _16358_ (.A(_09335_),
    .B(_09449_),
    .Y(_09450_));
 sky130_fd_sc_hd__mux2_1 _16359_ (.A0(net8207),
    .A1(net8214),
    .S(_08111_),
    .X(_09451_));
 sky130_fd_sc_hd__and2_1 _16360_ (.A(_09450_),
    .B(net8520),
    .X(_09452_));
 sky130_fd_sc_hd__or2_1 _16361_ (.A(_09450_),
    .B(net8520),
    .X(_09453_));
 sky130_fd_sc_hd__and2b_1 _16362_ (.A_N(_09452_),
    .B(_09453_),
    .X(_09454_));
 sky130_fd_sc_hd__o21ai_2 _16363_ (.A1(_09330_),
    .A2(_09331_),
    .B1(_09328_),
    .Y(_09455_));
 sky130_fd_sc_hd__xnor2_1 _16364_ (.A(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__nor2_1 _16365_ (.A(net7779),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__a21o_1 _16366_ (.A1(net7779),
    .A2(_09456_),
    .B1(net3454),
    .X(_09458_));
 sky130_fd_sc_hd__o221a_1 _16367_ (.A1(net3502),
    .A2(_08115_),
    .B1(_09457_),
    .B2(_09458_),
    .C1(_01633_),
    .X(_00469_));
 sky130_fd_sc_hd__a21o_1 _16368_ (.A1(_09336_),
    .A2(_09321_),
    .B1(_09448_),
    .X(_09459_));
 sky130_fd_sc_hd__o31a_4 _16369_ (.A1(_09323_),
    .A2(_09325_),
    .A3(_09449_),
    .B1(_09459_),
    .X(_09460_));
 sky130_fd_sc_hd__nor2_2 _16370_ (.A(_09446_),
    .B(_09447_),
    .Y(_09461_));
 sky130_fd_sc_hd__a21o_1 _16371_ (.A1(_09338_),
    .A2(_09444_),
    .B1(_09443_),
    .X(_09462_));
 sky130_fd_sc_hd__or2b_1 _16372_ (.A(_09369_),
    .B_N(_09340_),
    .X(_09463_));
 sky130_fd_sc_hd__a21bo_2 _16373_ (.A1(_09342_),
    .A2(_09368_),
    .B1_N(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__a21o_1 _16374_ (.A1(_09349_),
    .A2(_09367_),
    .B1(_09365_),
    .X(_09465_));
 sky130_fd_sc_hd__or2b_1 _16375_ (.A(_09389_),
    .B_N(_09371_),
    .X(_09466_));
 sky130_fd_sc_hd__a21bo_1 _16376_ (.A1(_09372_),
    .A2(_09388_),
    .B1_N(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__or3_1 _16377_ (.A(_08543_),
    .B(_09225_),
    .C(_09347_),
    .X(_09468_));
 sky130_fd_sc_hd__o21ai_1 _16378_ (.A1(_08543_),
    .A2(_09225_),
    .B1(_09347_),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_1 _16379_ (.A(_09468_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__or3b_2 _16380_ (.A(_06124_),
    .B(_09413_),
    .C_N(net7837),
    .X(_09471_));
 sky130_fd_sc_hd__buf_2 _16381_ (.A(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__nor2_1 _16382_ (.A(_08611_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__xnor2_1 _16383_ (.A(_09470_),
    .B(_09473_),
    .Y(_09474_));
 sky130_fd_sc_hd__nand2_1 _16384_ (.A(_09348_),
    .B(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__or2_1 _16385_ (.A(_09348_),
    .B(_09474_),
    .X(_09476_));
 sky130_fd_sc_hd__and2_1 _16386_ (.A(_09475_),
    .B(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__a21o_1 _16387_ (.A1(_09357_),
    .A2(_09358_),
    .B1(_09356_),
    .X(_09478_));
 sky130_fd_sc_hd__nor2_1 _16388_ (.A(_08542_),
    .B(_09115_),
    .Y(_09479_));
 sky130_fd_sc_hd__o21ai_1 _16389_ (.A1(_08226_),
    .A2(_08614_),
    .B1(_09355_),
    .Y(_09480_));
 sky130_fd_sc_hd__nand2_1 _16390_ (.A(_08864_),
    .B(_09354_),
    .Y(_09481_));
 sky130_fd_sc_hd__or2_1 _16391_ (.A(_09352_),
    .B(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__and3_1 _16392_ (.A(_09479_),
    .B(_09480_),
    .C(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__a21oi_1 _16393_ (.A1(_09480_),
    .A2(_09482_),
    .B1(_09479_),
    .Y(_09484_));
 sky130_fd_sc_hd__or2_1 _16394_ (.A(_09483_),
    .B(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__nand2_1 _16395_ (.A(_09374_),
    .B(_09375_),
    .Y(_09486_));
 sky130_fd_sc_hd__a21o_1 _16396_ (.A1(_09486_),
    .A2(_09378_),
    .B1(_09376_),
    .X(_09487_));
 sky130_fd_sc_hd__and2b_1 _16397_ (.A_N(_09485_),
    .B(_09487_),
    .X(_09488_));
 sky130_fd_sc_hd__and2b_1 _16398_ (.A_N(_09487_),
    .B(_09485_),
    .X(_09489_));
 sky130_fd_sc_hd__nor2_1 _16399_ (.A(_09488_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__xnor2_1 _16400_ (.A(_09478_),
    .B(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__a21oi_1 _16401_ (.A1(_09350_),
    .A2(_09362_),
    .B1(_09360_),
    .Y(_09492_));
 sky130_fd_sc_hd__nor2_1 _16402_ (.A(_09491_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__and2_1 _16403_ (.A(_09491_),
    .B(_09492_),
    .X(_09494_));
 sky130_fd_sc_hd__nor2_1 _16404_ (.A(_09493_),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__xor2_2 _16405_ (.A(_09477_),
    .B(_09495_),
    .X(_09496_));
 sky130_fd_sc_hd__xnor2_2 _16406_ (.A(_09467_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__xnor2_4 _16407_ (.A(_09465_),
    .B(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__or2b_1 _16408_ (.A(_09385_),
    .B_N(_09386_),
    .X(_09499_));
 sky130_fd_sc_hd__a21bo_1 _16409_ (.A1(_09379_),
    .A2(_09387_),
    .B1_N(_09499_),
    .X(_09500_));
 sky130_fd_sc_hd__or2b_1 _16410_ (.A(_09400_),
    .B_N(_09391_),
    .X(_09501_));
 sky130_fd_sc_hd__a22o_1 _16411_ (.A1(_08996_),
    .A2(_08167_),
    .B1(_09373_),
    .B2(_09135_),
    .X(_09502_));
 sky130_fd_sc_hd__nand2_1 _16412_ (.A(_09135_),
    .B(_08167_),
    .Y(_09503_));
 sky130_fd_sc_hd__or2_1 _16413_ (.A(_09374_),
    .B(_09503_),
    .X(_09504_));
 sky130_fd_sc_hd__nand2_1 _16414_ (.A(_09502_),
    .B(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__and2_1 _16415_ (.A(_09249_),
    .B(_09254_),
    .X(_09506_));
 sky130_fd_sc_hd__xnor2_2 _16416_ (.A(_09505_),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__or2_1 _16417_ (.A(_08306_),
    .B(_08418_),
    .X(_09508_));
 sky130_fd_sc_hd__or3_1 _16418_ (.A(_08308_),
    .B(_08403_),
    .C(_09508_),
    .X(_09509_));
 sky130_fd_sc_hd__o21ai_1 _16419_ (.A1(_08326_),
    .A2(_08403_),
    .B1(_09508_),
    .Y(_09510_));
 sky130_fd_sc_hd__and2_1 _16420_ (.A(_09509_),
    .B(_09510_),
    .X(_09511_));
 sky130_fd_sc_hd__nor2_1 _16421_ (.A(_09262_),
    .B(_08392_),
    .Y(_09512_));
 sky130_fd_sc_hd__xnor2_1 _16422_ (.A(_09511_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__a21boi_1 _16423_ (.A1(_09383_),
    .A2(_09384_),
    .B1_N(_09381_),
    .Y(_09514_));
 sky130_fd_sc_hd__nor2_1 _16424_ (.A(_09513_),
    .B(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__and2_1 _16425_ (.A(_09513_),
    .B(_09514_),
    .X(_09516_));
 sky130_fd_sc_hd__nor2_1 _16426_ (.A(_09515_),
    .B(_09516_),
    .Y(_09517_));
 sky130_fd_sc_hd__xnor2_1 _16427_ (.A(_09507_),
    .B(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__a21o_1 _16428_ (.A1(_09398_),
    .A2(_09501_),
    .B1(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__nand3_1 _16429_ (.A(_09398_),
    .B(_09501_),
    .C(_09518_),
    .Y(_09520_));
 sky130_fd_sc_hd__nand2_1 _16430_ (.A(_09519_),
    .B(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__xnor2_1 _16431_ (.A(_09500_),
    .B(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__a32o_1 _16432_ (.A1(_08244_),
    .A2(_08430_),
    .A3(_09392_),
    .B1(_09394_),
    .B2(_09395_),
    .X(_09523_));
 sky130_fd_sc_hd__a21oi_1 _16433_ (.A1(_09402_),
    .A2(_09406_),
    .B1(_09405_),
    .Y(_09524_));
 sky130_fd_sc_hd__nand2_1 _16434_ (.A(_08246_),
    .B(_08430_),
    .Y(_09525_));
 sky130_fd_sc_hd__nor2_1 _16435_ (.A(_08880_),
    .B(_09165_),
    .Y(_09526_));
 sky130_fd_sc_hd__xnor2_1 _16436_ (.A(_09525_),
    .B(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__nor2_1 _16437_ (.A(_08509_),
    .B(_08411_),
    .Y(_09528_));
 sky130_fd_sc_hd__xnor2_1 _16438_ (.A(_09527_),
    .B(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__or2_1 _16439_ (.A(_09524_),
    .B(_09529_),
    .X(_09530_));
 sky130_fd_sc_hd__nand2_1 _16440_ (.A(_09524_),
    .B(_09529_),
    .Y(_09531_));
 sky130_fd_sc_hd__nand2_1 _16441_ (.A(_09530_),
    .B(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__xnor2_2 _16442_ (.A(_09523_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__or4_1 _16443_ (.A(_08401_),
    .B(_08916_),
    .C(_09292_),
    .D(_09411_),
    .X(_09534_));
 sky130_fd_sc_hd__o22ai_1 _16444_ (.A1(_08916_),
    .A2(_09403_),
    .B1(_09411_),
    .B2(_08948_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand2_1 _16445_ (.A(_09534_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__clkbuf_4 _16446_ (.A(_08417_),
    .X(_09537_));
 sky130_fd_sc_hd__nor2_1 _16447_ (.A(_09537_),
    .B(_09170_),
    .Y(_09538_));
 sky130_fd_sc_hd__xnor2_2 _16448_ (.A(_09536_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__a21o_2 _16449_ (.A1(_09419_),
    .A2(_09296_),
    .B1(_06123_),
    .X(_09540_));
 sky130_fd_sc_hd__nand2_2 _16450_ (.A(net4520),
    .B(_06123_),
    .Y(_09541_));
 sky130_fd_sc_hd__a21oi_2 _16451_ (.A1(_09540_),
    .A2(_09541_),
    .B1(_08905_),
    .Y(_09542_));
 sky130_fd_sc_hd__inv_2 _16452_ (.A(_08030_),
    .Y(_09543_));
 sky130_fd_sc_hd__a31o_1 _16453_ (.A1(_08024_),
    .A2(_09414_),
    .A3(net75),
    .B1(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__or4b_1 _16454_ (.A(_08025_),
    .B(_08028_),
    .C(_08030_),
    .D_N(net75),
    .X(_09545_));
 sky130_fd_sc_hd__a31o_2 _16455_ (.A1(_08421_),
    .A2(_09544_),
    .A3(_09545_),
    .B1(_08442_),
    .X(_09546_));
 sky130_fd_sc_hd__or4_4 _16456_ (.A(net8041),
    .B(_06123_),
    .C(_09413_),
    .D(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__nand2_1 _16457_ (.A(net3724),
    .B(_09413_),
    .Y(_09548_));
 sky130_fd_sc_hd__a21oi_2 _16458_ (.A1(_09548_),
    .A2(_09417_),
    .B1(_08474_),
    .Y(_09549_));
 sky130_fd_sc_hd__xnor2_2 _16459_ (.A(_09547_),
    .B(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__xor2_2 _16460_ (.A(_09542_),
    .B(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__a21oi_1 _16461_ (.A1(_09548_),
    .A2(_09417_),
    .B1(_06124_),
    .Y(_09552_));
 sky130_fd_sc_hd__a32o_1 _16462_ (.A1(_08446_),
    .A2(_09552_),
    .A3(_09420_),
    .B1(_09421_),
    .B2(_09412_),
    .X(_09553_));
 sky130_fd_sc_hd__xor2_2 _16463_ (.A(_09551_),
    .B(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__xnor2_2 _16464_ (.A(_09539_),
    .B(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__or2b_1 _16465_ (.A(_09422_),
    .B_N(_09424_),
    .X(_09556_));
 sky130_fd_sc_hd__a21bo_1 _16466_ (.A1(_09408_),
    .A2(_09425_),
    .B1_N(_09556_),
    .X(_09557_));
 sky130_fd_sc_hd__xnor2_2 _16467_ (.A(_09555_),
    .B(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__xnor2_1 _16468_ (.A(_09533_),
    .B(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__and2b_1 _16469_ (.A_N(_09426_),
    .B(_09428_),
    .X(_09560_));
 sky130_fd_sc_hd__a21oi_1 _16470_ (.A1(_09401_),
    .A2(_09429_),
    .B1(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__nor2_1 _16471_ (.A(_09559_),
    .B(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__nand2_1 _16472_ (.A(_09559_),
    .B(_09561_),
    .Y(_09563_));
 sky130_fd_sc_hd__and2b_1 _16473_ (.A_N(_09562_),
    .B(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__xnor2_1 _16474_ (.A(_09522_),
    .B(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__a21oi_1 _16475_ (.A1(_09390_),
    .A2(_09434_),
    .B1(_09433_),
    .Y(_09566_));
 sky130_fd_sc_hd__nor2_1 _16476_ (.A(_09565_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand2_1 _16477_ (.A(_09565_),
    .B(_09566_),
    .Y(_09568_));
 sky130_fd_sc_hd__and2b_1 _16478_ (.A_N(_09567_),
    .B(_09568_),
    .X(_09569_));
 sky130_fd_sc_hd__xnor2_4 _16479_ (.A(_09498_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__nor2_1 _16480_ (.A(_09436_),
    .B(_09438_),
    .Y(_09571_));
 sky130_fd_sc_hd__a21oi_4 _16481_ (.A1(_09370_),
    .A2(_09439_),
    .B1(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__xor2_4 _16482_ (.A(_09570_),
    .B(_09572_),
    .X(_09573_));
 sky130_fd_sc_hd__xnor2_4 _16483_ (.A(_09464_),
    .B(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__xnor2_4 _16484_ (.A(_09462_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__xor2_4 _16485_ (.A(_09461_),
    .B(_09575_),
    .X(_09576_));
 sky130_fd_sc_hd__xnor2_4 _16486_ (.A(_09460_),
    .B(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(net8225),
    .A1(net7771),
    .S(_08111_),
    .X(_09578_));
 sky130_fd_sc_hd__nor2_1 _16488_ (.A(_09577_),
    .B(net7772),
    .Y(_09579_));
 sky130_fd_sc_hd__and2_1 _16489_ (.A(_09577_),
    .B(net7772),
    .X(_09580_));
 sky130_fd_sc_hd__nor2_1 _16490_ (.A(_09579_),
    .B(_09580_),
    .Y(_09581_));
 sky130_fd_sc_hd__a21oi_1 _16491_ (.A1(_09453_),
    .A2(_09455_),
    .B1(_09452_),
    .Y(_09582_));
 sky130_fd_sc_hd__xor2_1 _16492_ (.A(net7779),
    .B(_09582_),
    .X(_09583_));
 sky130_fd_sc_hd__nor2_1 _16493_ (.A(_09581_),
    .B(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__a21o_1 _16494_ (.A1(_09581_),
    .A2(_09583_),
    .B1(net3454),
    .X(_09585_));
 sky130_fd_sc_hd__o221a_1 _16495_ (.A1(net4769),
    .A2(_08115_),
    .B1(_09584_),
    .B2(_09585_),
    .C1(_01633_),
    .X(_00470_));
 sky130_fd_sc_hd__o21ba_1 _16496_ (.A1(_09579_),
    .A2(_09582_),
    .B1_N(_09580_),
    .X(_09586_));
 sky130_fd_sc_hd__inv_2 _16497_ (.A(_09576_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand2_1 _16498_ (.A(_09461_),
    .B(_09575_),
    .Y(_09588_));
 sky130_fd_sc_hd__o21ai_4 _16499_ (.A1(_09460_),
    .A2(_09587_),
    .B1(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__or2b_1 _16500_ (.A(_09574_),
    .B_N(_09462_),
    .X(_09590_));
 sky130_fd_sc_hd__or2b_1 _16501_ (.A(_09497_),
    .B_N(_09465_),
    .X(_09591_));
 sky130_fd_sc_hd__a21boi_1 _16502_ (.A1(_09467_),
    .A2(_09496_),
    .B1_N(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__xor2_1 _16503_ (.A(_09475_),
    .B(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__and3_1 _16504_ (.A(net8034),
    .B(_08181_),
    .C(_08129_),
    .X(_09594_));
 sky130_fd_sc_hd__nand2_1 _16505_ (.A(_08611_),
    .B(net7818),
    .Y(_09595_));
 sky130_fd_sc_hd__xnor2_1 _16506_ (.A(_09593_),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__a21o_1 _16507_ (.A1(_09477_),
    .A2(_09495_),
    .B1(_09493_),
    .X(_09597_));
 sky130_fd_sc_hd__or2b_1 _16508_ (.A(_09521_),
    .B_N(_09500_),
    .X(_09598_));
 sky130_fd_sc_hd__nor2_1 _16509_ (.A(_08543_),
    .B(_09345_),
    .Y(_09599_));
 sky130_fd_sc_hd__inv_2 _16510_ (.A(_09116_),
    .Y(_09600_));
 sky130_fd_sc_hd__a2bb2o_1 _16511_ (.A1_N(_09224_),
    .A2_N(_08542_),
    .B1(_09133_),
    .B2(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__nor2_1 _16512_ (.A(_06124_),
    .B(net4908),
    .Y(_09602_));
 sky130_fd_sc_hd__and2_1 _16513_ (.A(_09133_),
    .B(net4909),
    .X(_09603_));
 sky130_fd_sc_hd__nand2_1 _16514_ (.A(_09479_),
    .B(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__and3_1 _16515_ (.A(_09599_),
    .B(_09601_),
    .C(_09604_),
    .X(_09605_));
 sky130_fd_sc_hd__a21oi_1 _16516_ (.A1(_09601_),
    .A2(_09604_),
    .B1(_09599_),
    .Y(_09606_));
 sky130_fd_sc_hd__or2_1 _16517_ (.A(_09605_),
    .B(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__o31a_1 _16518_ (.A1(_08611_),
    .A2(_09470_),
    .A3(_09472_),
    .B1(_09468_),
    .X(_09608_));
 sky130_fd_sc_hd__nor2_1 _16519_ (.A(_09607_),
    .B(_09608_),
    .Y(_09609_));
 sky130_fd_sc_hd__and2_1 _16520_ (.A(_09607_),
    .B(_09608_),
    .X(_09610_));
 sky130_fd_sc_hd__nor2_1 _16521_ (.A(_09609_),
    .B(_09610_),
    .Y(_09611_));
 sky130_fd_sc_hd__buf_4 _16522_ (.A(_09472_),
    .X(_09612_));
 sky130_fd_sc_hd__nor2_1 _16523_ (.A(_08127_),
    .B(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__xor2_1 _16524_ (.A(_09611_),
    .B(_09613_),
    .X(_09614_));
 sky130_fd_sc_hd__a21bo_1 _16525_ (.A1(_09479_),
    .A2(_09480_),
    .B1_N(_09482_),
    .X(_09615_));
 sky130_fd_sc_hd__or2b_1 _16526_ (.A(_09505_),
    .B_N(_09506_),
    .X(_09616_));
 sky130_fd_sc_hd__and2_2 _16527_ (.A(_08185_),
    .B(_09351_),
    .X(_09617_));
 sky130_fd_sc_hd__a22o_1 _16528_ (.A1(_09373_),
    .A2(_09254_),
    .B1(_09351_),
    .B2(_09249_),
    .X(_09618_));
 sky130_fd_sc_hd__a21boi_1 _16529_ (.A1(_09506_),
    .A2(_09617_),
    .B1_N(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__xor2_1 _16530_ (.A(_09481_),
    .B(_09619_),
    .X(_09620_));
 sky130_fd_sc_hd__a21oi_1 _16531_ (.A1(_09504_),
    .A2(_09616_),
    .B1(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__and3_1 _16532_ (.A(_09504_),
    .B(_09616_),
    .C(_09620_),
    .X(_09622_));
 sky130_fd_sc_hd__nor2_1 _16533_ (.A(_09621_),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__xnor2_1 _16534_ (.A(_09615_),
    .B(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__a21oi_1 _16535_ (.A1(_09478_),
    .A2(_09490_),
    .B1(_09488_),
    .Y(_09625_));
 sky130_fd_sc_hd__nor2_1 _16536_ (.A(_09624_),
    .B(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__and2_1 _16537_ (.A(_09624_),
    .B(_09625_),
    .X(_09627_));
 sky130_fd_sc_hd__nor2_1 _16538_ (.A(_09626_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__xnor2_1 _16539_ (.A(_09614_),
    .B(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__a21o_1 _16540_ (.A1(_09519_),
    .A2(_09598_),
    .B1(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__nand3_1 _16541_ (.A(_09519_),
    .B(_09598_),
    .C(_09629_),
    .Y(_09631_));
 sky130_fd_sc_hd__nand2_1 _16542_ (.A(_09630_),
    .B(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__xnor2_1 _16543_ (.A(_09597_),
    .B(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__a21o_1 _16544_ (.A1(_09507_),
    .A2(_09517_),
    .B1(_09515_),
    .X(_09634_));
 sky130_fd_sc_hd__or2b_1 _16545_ (.A(_09532_),
    .B_N(_09523_),
    .X(_09635_));
 sky130_fd_sc_hd__or2_2 _16546_ (.A(_08323_),
    .B(_08418_),
    .X(_09636_));
 sky130_fd_sc_hd__nor2_1 _16547_ (.A(_08338_),
    .B(_08383_),
    .Y(_09637_));
 sky130_fd_sc_hd__xnor2_1 _16548_ (.A(_09636_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__xnor2_1 _16549_ (.A(_09503_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__nor2_1 _16550_ (.A(_08799_),
    .B(_08403_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2_1 _16551_ (.A(_08509_),
    .B(_09025_),
    .Y(_09641_));
 sky130_fd_sc_hd__nor2_1 _16552_ (.A(_08326_),
    .B(_08411_),
    .Y(_09642_));
 sky130_fd_sc_hd__xor2_1 _16553_ (.A(_09641_),
    .B(_09642_),
    .X(_09643_));
 sky130_fd_sc_hd__xnor2_1 _16554_ (.A(_09640_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__a21boi_1 _16555_ (.A1(_09511_),
    .A2(_09512_),
    .B1_N(_09509_),
    .Y(_09645_));
 sky130_fd_sc_hd__nor2_1 _16556_ (.A(_09644_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__nand2_1 _16557_ (.A(_09644_),
    .B(_09645_),
    .Y(_09647_));
 sky130_fd_sc_hd__and2b_1 _16558_ (.A_N(_09646_),
    .B(_09647_),
    .X(_09648_));
 sky130_fd_sc_hd__xnor2_1 _16559_ (.A(_09639_),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21o_1 _16560_ (.A1(_09530_),
    .A2(_09635_),
    .B1(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__nand3_1 _16561_ (.A(_09530_),
    .B(_09635_),
    .C(_09649_),
    .Y(_09651_));
 sky130_fd_sc_hd__nand2_1 _16562_ (.A(_09650_),
    .B(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__xnor2_2 _16563_ (.A(_09634_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__and2_1 _16564_ (.A(_09527_),
    .B(_09528_),
    .X(_09654_));
 sky130_fd_sc_hd__a31o_1 _16565_ (.A1(_08246_),
    .A2(_08430_),
    .A3(_09526_),
    .B1(_09654_),
    .X(_09655_));
 sky130_fd_sc_hd__a21bo_1 _16566_ (.A1(_09535_),
    .A2(_09538_),
    .B1_N(_09534_),
    .X(_09656_));
 sky130_fd_sc_hd__or2_1 _16567_ (.A(_08391_),
    .B(_09165_),
    .X(_09657_));
 sky130_fd_sc_hd__and4b_1 _16568_ (.A_N(_09403_),
    .B(_08244_),
    .C(_08666_),
    .D(_09288_),
    .X(_09658_));
 sky130_fd_sc_hd__o22a_1 _16569_ (.A1(_08880_),
    .A2(_09170_),
    .B1(_09403_),
    .B2(_08417_),
    .X(_09659_));
 sky130_fd_sc_hd__nor2_1 _16570_ (.A(_09658_),
    .B(_09659_),
    .Y(_09660_));
 sky130_fd_sc_hd__xnor2_1 _16571_ (.A(_09657_),
    .B(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__xor2_1 _16572_ (.A(_09656_),
    .B(_09661_),
    .X(_09662_));
 sky130_fd_sc_hd__xor2_1 _16573_ (.A(_09655_),
    .B(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__clkbuf_4 _16574_ (.A(_09411_),
    .X(_09664_));
 sky130_fd_sc_hd__nor2_1 _16575_ (.A(_08916_),
    .B(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__a21o_2 _16576_ (.A1(_09548_),
    .A2(_09417_),
    .B1(_06123_),
    .X(_09666_));
 sky130_fd_sc_hd__nand2_2 _16577_ (.A(net3934),
    .B(_06123_),
    .Y(_09667_));
 sky130_fd_sc_hd__a21o_1 _16578_ (.A1(_09666_),
    .A2(_09667_),
    .B1(_08905_),
    .X(_09668_));
 sky130_fd_sc_hd__a21oi_2 _16579_ (.A1(_09540_),
    .A2(_09541_),
    .B1(_08401_),
    .Y(_09669_));
 sky130_fd_sc_hd__xnor2_2 _16580_ (.A(_09668_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__xor2_2 _16581_ (.A(_09665_),
    .B(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__o21ai_1 _16582_ (.A1(_08032_),
    .A2(_09545_),
    .B1(_08421_),
    .Y(_09672_));
 sky130_fd_sc_hd__a22o_2 _16583_ (.A1(net3507),
    .A2(_09413_),
    .B1(_08441_),
    .B2(_09672_),
    .X(_09673_));
 sky130_fd_sc_hd__a21o_1 _16584_ (.A1(_08573_),
    .A2(_09673_),
    .B1(net4891),
    .X(_09674_));
 sky130_fd_sc_hd__or3b_1 _16585_ (.A(net8035),
    .B(_08494_),
    .C_N(_09673_),
    .X(_09675_));
 sky130_fd_sc_hd__nand2_1 _16586_ (.A(net3587),
    .B(_09413_),
    .Y(_09676_));
 sky130_fd_sc_hd__a21oi_1 _16587_ (.A1(_09676_),
    .A2(_09546_),
    .B1(_08474_),
    .Y(_09677_));
 sky130_fd_sc_hd__nand3_1 _16588_ (.A(_09674_),
    .B(_09675_),
    .C(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__a21o_1 _16589_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09677_),
    .X(_09679_));
 sky130_fd_sc_hd__a21oi_1 _16590_ (.A1(_09676_),
    .A2(_09546_),
    .B1(_06124_),
    .Y(_09680_));
 sky130_fd_sc_hd__a32o_1 _16591_ (.A1(_08446_),
    .A2(_09680_),
    .A3(_09549_),
    .B1(_09550_),
    .B2(_09542_),
    .X(_09681_));
 sky130_fd_sc_hd__nand3_1 _16592_ (.A(_09678_),
    .B(_09679_),
    .C(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__a21o_1 _16593_ (.A1(_09678_),
    .A2(_09679_),
    .B1(_09681_),
    .X(_09683_));
 sky130_fd_sc_hd__nand3_1 _16594_ (.A(_09671_),
    .B(_09682_),
    .C(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__a21o_1 _16595_ (.A1(_09682_),
    .A2(_09683_),
    .B1(_09671_),
    .X(_09685_));
 sky130_fd_sc_hd__nand2_1 _16596_ (.A(_09551_),
    .B(_09553_),
    .Y(_09686_));
 sky130_fd_sc_hd__a21bo_1 _16597_ (.A1(_09539_),
    .A2(_09554_),
    .B1_N(_09686_),
    .X(_09687_));
 sky130_fd_sc_hd__nand3_1 _16598_ (.A(_09684_),
    .B(_09685_),
    .C(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__a21o_1 _16599_ (.A1(_09684_),
    .A2(_09685_),
    .B1(_09687_),
    .X(_09689_));
 sky130_fd_sc_hd__and3_1 _16600_ (.A(_09663_),
    .B(_09688_),
    .C(_09689_),
    .X(_09690_));
 sky130_fd_sc_hd__a21oi_1 _16601_ (.A1(_09688_),
    .A2(_09689_),
    .B1(_09663_),
    .Y(_09691_));
 sky130_fd_sc_hd__or2_2 _16602_ (.A(_09690_),
    .B(_09691_),
    .X(_09692_));
 sky130_fd_sc_hd__and2b_1 _16603_ (.A_N(_09555_),
    .B(_09557_),
    .X(_09693_));
 sky130_fd_sc_hd__a21oi_2 _16604_ (.A1(_09533_),
    .A2(_09558_),
    .B1(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__xor2_2 _16605_ (.A(_09692_),
    .B(_09694_),
    .X(_09695_));
 sky130_fd_sc_hd__xnor2_2 _16606_ (.A(_09653_),
    .B(_09695_),
    .Y(_09696_));
 sky130_fd_sc_hd__a21oi_1 _16607_ (.A1(_09522_),
    .A2(_09563_),
    .B1(_09562_),
    .Y(_09697_));
 sky130_fd_sc_hd__nor2_1 _16608_ (.A(_09696_),
    .B(_09697_),
    .Y(_09698_));
 sky130_fd_sc_hd__and2_1 _16609_ (.A(_09696_),
    .B(_09697_),
    .X(_09699_));
 sky130_fd_sc_hd__nor2_1 _16610_ (.A(_09698_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__xnor2_1 _16611_ (.A(_09633_),
    .B(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__a21oi_1 _16612_ (.A1(_09498_),
    .A2(_09568_),
    .B1(_09567_),
    .Y(_09702_));
 sky130_fd_sc_hd__xor2_1 _16613_ (.A(_09701_),
    .B(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__xnor2_1 _16614_ (.A(_09596_),
    .B(_09703_),
    .Y(_09704_));
 sky130_fd_sc_hd__nor2_1 _16615_ (.A(_09570_),
    .B(_09572_),
    .Y(_09705_));
 sky130_fd_sc_hd__a21oi_1 _16616_ (.A1(_09464_),
    .A2(_09573_),
    .B1(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__nor2_1 _16617_ (.A(_09704_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__and2_1 _16618_ (.A(_09704_),
    .B(_09706_),
    .X(_09708_));
 sky130_fd_sc_hd__or2_1 _16619_ (.A(_09707_),
    .B(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__xnor2_2 _16620_ (.A(_09590_),
    .B(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__xnor2_4 _16621_ (.A(_09589_),
    .B(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__mux2_1 _16622_ (.A0(net4188),
    .A1(net2898),
    .S(_08111_),
    .X(_09712_));
 sky130_fd_sc_hd__xnor2_1 _16623_ (.A(_09105_),
    .B(net4189),
    .Y(_09713_));
 sky130_fd_sc_hd__xnor2_1 _16624_ (.A(_09711_),
    .B(net4190),
    .Y(_09714_));
 sky130_fd_sc_hd__and2_1 _16625_ (.A(_09586_),
    .B(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__o21ai_1 _16626_ (.A1(_09586_),
    .A2(_09714_),
    .B1(_08115_),
    .Y(_09716_));
 sky130_fd_sc_hd__o221a_1 _16627_ (.A1(net7752),
    .A2(_08115_),
    .B1(_09715_),
    .B2(_09716_),
    .C1(_01633_),
    .X(_00471_));
 sky130_fd_sc_hd__and3_1 _16628_ (.A(_04684_),
    .B(_04648_),
    .C(_05057_),
    .X(_09717_));
 sky130_fd_sc_hd__and3_1 _16629_ (.A(_04665_),
    .B(net4121),
    .C(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__or2_1 _16630_ (.A(_04458_),
    .B(net4122),
    .X(_09719_));
 sky130_fd_sc_hd__clkbuf_2 _16631_ (.A(net4123),
    .X(_09720_));
 sky130_fd_sc_hd__nor2_1 _16632_ (.A(_04021_),
    .B(net4124),
    .Y(_00472_));
 sky130_fd_sc_hd__buf_4 _16633_ (.A(_08092_),
    .X(_09721_));
 sky130_fd_sc_hd__or2_1 _16634_ (.A(_04496_),
    .B(_04021_),
    .X(_09722_));
 sky130_fd_sc_hd__and3_1 _16635_ (.A(_09721_),
    .B(net3858),
    .C(_09722_),
    .X(_09723_));
 sky130_fd_sc_hd__clkbuf_1 _16636_ (.A(net3859),
    .X(_00473_));
 sky130_fd_sc_hd__nand2_1 _16637_ (.A(net3955),
    .B(net3858),
    .Y(_09724_));
 sky130_fd_sc_hd__buf_4 _16638_ (.A(_08092_),
    .X(_09725_));
 sky130_fd_sc_hd__and3b_1 _16639_ (.A_N(net7679),
    .B(net3956),
    .C(_09725_),
    .X(_09726_));
 sky130_fd_sc_hd__clkbuf_1 _16640_ (.A(net3957),
    .X(_00474_));
 sky130_fd_sc_hd__nor2_1 _16641_ (.A(net3919),
    .B(net4124),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_4 _16642_ (.A(_04458_),
    .B(net4122),
    .Y(_09727_));
 sky130_fd_sc_hd__and3_1 _16643_ (.A(_04666_),
    .B(net4058),
    .C(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__clkbuf_1 _16644_ (.A(net4059),
    .X(_00476_));
 sky130_fd_sc_hd__nor2_1 _16645_ (.A(net4108),
    .B(net4124),
    .Y(_00477_));
 sky130_fd_sc_hd__nor2_1 _16646_ (.A(net3517),
    .B(net4124),
    .Y(_00478_));
 sky130_fd_sc_hd__nor2_1 _16647_ (.A(net4118),
    .B(net4124),
    .Y(_00479_));
 sky130_fd_sc_hd__and3_1 _16648_ (.A(net4133),
    .B(_04664_),
    .C(net5948),
    .X(_09729_));
 sky130_fd_sc_hd__a31o_1 _16649_ (.A1(_04466_),
    .A2(_04664_),
    .A3(_05184_),
    .B1(net4133),
    .X(_09730_));
 sky130_fd_sc_hd__and3b_1 _16650_ (.A_N(net5949),
    .B(_09727_),
    .C(net4134),
    .X(_09731_));
 sky130_fd_sc_hd__clkbuf_1 _16651_ (.A(net4135),
    .X(_00480_));
 sky130_fd_sc_hd__a21oi_1 _16652_ (.A1(net4089),
    .A2(net5949),
    .B1(_09720_),
    .Y(_09732_));
 sky130_fd_sc_hd__o21a_1 _16653_ (.A1(net4089),
    .A2(net5949),
    .B1(_09732_),
    .X(_00481_));
 sky130_fd_sc_hd__inv_2 _16654_ (.A(net4122),
    .Y(_09733_));
 sky130_fd_sc_hd__or3_4 _16655_ (.A(net3452),
    .B(net3628),
    .C(_09733_),
    .X(_09734_));
 sky130_fd_sc_hd__and2_2 _16656_ (.A(_04479_),
    .B(_09734_),
    .X(_09735_));
 sky130_fd_sc_hd__clkbuf_8 _16657_ (.A(_09735_),
    .X(_09736_));
 sky130_fd_sc_hd__clkbuf_4 _16658_ (.A(_09736_),
    .X(_09737_));
 sky130_fd_sc_hd__nor2_4 _16659_ (.A(_04478_),
    .B(_09734_),
    .Y(_09738_));
 sky130_fd_sc_hd__buf_4 _16660_ (.A(_09738_),
    .X(_09739_));
 sky130_fd_sc_hd__clkbuf_4 _16661_ (.A(_09739_),
    .X(_09740_));
 sky130_fd_sc_hd__a22o_1 _16662_ (.A1(net4080),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_08111_),
    .X(_00482_));
 sky130_fd_sc_hd__a22o_1 _16663_ (.A1(net4246),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07917_),
    .X(_00483_));
 sky130_fd_sc_hd__a22o_1 _16664_ (.A1(net4343),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07929_),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _16665_ (.A1(net4339),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07938_),
    .X(_00485_));
 sky130_fd_sc_hd__a22o_1 _16666_ (.A1(net4303),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07947_),
    .X(_00486_));
 sky130_fd_sc_hd__a22o_1 _16667_ (.A1(net4407),
    .A2(_09737_),
    .B1(_09740_),
    .B2(net7825),
    .X(_00487_));
 sky130_fd_sc_hd__a22o_1 _16668_ (.A1(net4305),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07962_),
    .X(_00488_));
 sky130_fd_sc_hd__a22o_1 _16669_ (.A1(net4512),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07968_),
    .X(_00489_));
 sky130_fd_sc_hd__a22o_1 _16670_ (.A1(net4615),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07975_),
    .X(_00490_));
 sky130_fd_sc_hd__a22o_1 _16671_ (.A1(net4361),
    .A2(_09737_),
    .B1(_09740_),
    .B2(_07981_),
    .X(_00491_));
 sky130_fd_sc_hd__buf_4 _16672_ (.A(_09736_),
    .X(_09741_));
 sky130_fd_sc_hd__buf_4 _16673_ (.A(_09739_),
    .X(_09742_));
 sky130_fd_sc_hd__a22o_1 _16674_ (.A1(net4341),
    .A2(_09741_),
    .B1(_09742_),
    .B2(_07991_),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _16675_ (.A1(net4194),
    .A2(_09741_),
    .B1(_09742_),
    .B2(_07998_),
    .X(_00493_));
 sky130_fd_sc_hd__a22o_1 _16676_ (.A1(net4321),
    .A2(_09741_),
    .B1(_09742_),
    .B2(net672),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _16677_ (.A1(net4259),
    .A2(_09741_),
    .B1(_09742_),
    .B2(net1154),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _16678_ (.A1(net4335),
    .A2(_09741_),
    .B1(_09742_),
    .B2(net744),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_1 _16679_ (.A1(net4271),
    .A2(_09741_),
    .B1(_09742_),
    .B2(net3502),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _16680_ (.A1(net5596),
    .A2(_09741_),
    .B1(_09742_),
    .B2(net4769),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_1 _16681_ (.A1(net777),
    .A2(_09741_),
    .B1(_09742_),
    .B2(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _16682_ (.A1(net756),
    .A2(_09741_),
    .B1(_09742_),
    .B2(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _16683_ (.A1(net967),
    .A2(_09741_),
    .B1(_09742_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00501_));
 sky130_fd_sc_hd__clkbuf_4 _16684_ (.A(_09736_),
    .X(_09743_));
 sky130_fd_sc_hd__clkbuf_4 _16685_ (.A(_09738_),
    .X(_09744_));
 sky130_fd_sc_hd__a22o_1 _16686_ (.A1(net754),
    .A2(_09743_),
    .B1(_09744_),
    .B2(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _16687_ (.A1(net8126),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net4277),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _16688_ (.A1(net8132),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net4268),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _16689_ (.A1(net8138),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net4236),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _16690_ (.A1(net8141),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net4280),
    .X(_00506_));
 sky130_fd_sc_hd__a22o_1 _16691_ (.A1(net8123),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net4293),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _16692_ (.A1(net834),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net8018),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _16693_ (.A1(net822),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net8021),
    .X(_00509_));
 sky130_fd_sc_hd__a22o_1 _16694_ (.A1(net984),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net8029),
    .X(_00510_));
 sky130_fd_sc_hd__a22o_1 _16695_ (.A1(net8120),
    .A2(_09743_),
    .B1(_09744_),
    .B2(net4917),
    .X(_00511_));
 sky130_fd_sc_hd__clkbuf_4 _16696_ (.A(_09736_),
    .X(_09745_));
 sky130_fd_sc_hd__clkbuf_4 _16697_ (.A(_09738_),
    .X(_09746_));
 sky130_fd_sc_hd__a22o_1 _16698_ (.A1(net864),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net7999),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _16699_ (.A1(net1009),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net8012),
    .X(_00513_));
 sky130_fd_sc_hd__a22o_1 _16700_ (.A1(net1038),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net8009),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_1 _16701_ (.A1(net969),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net8015),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _16702_ (.A1(net1015),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net8002),
    .X(_00516_));
 sky130_fd_sc_hd__a22o_1 _16703_ (.A1(net971),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net8068),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _16704_ (.A1(net991),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net8088),
    .X(_00518_));
 sky130_fd_sc_hd__a22o_1 _16705_ (.A1(net8067),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net7837),
    .X(_00519_));
 sky130_fd_sc_hd__a22o_1 _16706_ (.A1(net8079),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net8034),
    .X(_00520_));
 sky130_fd_sc_hd__or2_4 _16707_ (.A(_04489_),
    .B(_09734_),
    .X(_09747_));
 sky130_fd_sc_hd__mux2_1 _16708_ (.A0(_04567_),
    .A1(net7665),
    .S(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__clkbuf_1 _16709_ (.A(net7667),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _16710_ (.A0(_04566_),
    .A1(net7609),
    .S(_09747_),
    .X(_09749_));
 sky130_fd_sc_hd__clkbuf_1 _16711_ (.A(net7611),
    .X(_00522_));
 sky130_fd_sc_hd__xor2_1 _16712_ (.A(net5554),
    .B(_09102_),
    .X(_09750_));
 sky130_fd_sc_hd__xor2_2 _16713_ (.A(net7631),
    .B(_09102_),
    .X(_09751_));
 sky130_fd_sc_hd__xnor2_2 _16714_ (.A(net4007),
    .B(_09102_),
    .Y(_09752_));
 sky130_fd_sc_hd__or2_1 _16715_ (.A(net3999),
    .B(_09102_),
    .X(_09753_));
 sky130_fd_sc_hd__xnor2_1 _16716_ (.A(_06068_),
    .B(_08194_),
    .Y(_09754_));
 sky130_fd_sc_hd__and2_1 _16717_ (.A(_06104_),
    .B(net7713),
    .X(_09755_));
 sky130_fd_sc_hd__a21o_1 _16718_ (.A1(net4034),
    .A2(_09102_),
    .B1(_09755_),
    .X(_09756_));
 sky130_fd_sc_hd__and2_1 _16719_ (.A(net3965),
    .B(_08194_),
    .X(_09757_));
 sky130_fd_sc_hd__nor2_1 _16720_ (.A(net3965),
    .B(_08194_),
    .Y(_09758_));
 sky130_fd_sc_hd__nor2_1 _16721_ (.A(_09757_),
    .B(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__a21o_1 _16722_ (.A1(_09756_),
    .A2(_09759_),
    .B1(_09757_),
    .X(_09760_));
 sky130_fd_sc_hd__nand2_1 _16723_ (.A(net3999),
    .B(_09102_),
    .Y(_09761_));
 sky130_fd_sc_hd__a21bo_1 _16724_ (.A1(_09753_),
    .A2(_09760_),
    .B1_N(_09761_),
    .X(_09762_));
 sky130_fd_sc_hd__o21a_1 _16725_ (.A1(net4049),
    .A2(net3884),
    .B1(_09103_),
    .X(_09763_));
 sky130_fd_sc_hd__a31o_1 _16726_ (.A1(_09751_),
    .A2(_09752_),
    .A3(_09762_),
    .B1(_09763_),
    .X(_09764_));
 sky130_fd_sc_hd__or2_1 _16727_ (.A(_09750_),
    .B(_09764_),
    .X(_09765_));
 sky130_fd_sc_hd__nand2_1 _16728_ (.A(_09750_),
    .B(_09764_),
    .Y(_09766_));
 sky130_fd_sc_hd__nand2_1 _16729_ (.A(net4647),
    .B(_08035_),
    .Y(_09767_));
 sky130_fd_sc_hd__nor2_2 _16730_ (.A(_06058_),
    .B(net4648),
    .Y(_09768_));
 sky130_fd_sc_hd__buf_4 _16731_ (.A(net4648),
    .X(_09769_));
 sky130_fd_sc_hd__a32o_1 _16732_ (.A1(_09765_),
    .A2(_09766_),
    .A3(_09768_),
    .B1(_09769_),
    .B2(net5554),
    .X(_00523_));
 sky130_fd_sc_hd__xor2_1 _16733_ (.A(net5666),
    .B(_09102_),
    .X(_09770_));
 sky130_fd_sc_hd__a21bo_1 _16734_ (.A1(net5554),
    .A2(_09103_),
    .B1_N(_09766_),
    .X(_09771_));
 sky130_fd_sc_hd__xor2_1 _16735_ (.A(_09770_),
    .B(_09771_),
    .X(_09772_));
 sky130_fd_sc_hd__a22o_1 _16736_ (.A1(net5666),
    .A2(_09769_),
    .B1(_09768_),
    .B2(_09772_),
    .X(_00524_));
 sky130_fd_sc_hd__xor2_1 _16737_ (.A(net5472),
    .B(_09102_),
    .X(_09773_));
 sky130_fd_sc_hd__and2_1 _16738_ (.A(_09752_),
    .B(_09762_),
    .X(_09774_));
 sky130_fd_sc_hd__and4_1 _16739_ (.A(_09750_),
    .B(_09751_),
    .C(_09774_),
    .D(_09770_),
    .X(_09775_));
 sky130_fd_sc_hd__o41a_1 _16740_ (.A1(net4049),
    .A2(net3884),
    .A3(net5666),
    .A4(net5554),
    .B1(_09102_),
    .X(_09776_));
 sky130_fd_sc_hd__or3_1 _16741_ (.A(_09773_),
    .B(_09775_),
    .C(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__o21ai_1 _16742_ (.A1(_09775_),
    .A2(_09776_),
    .B1(_09773_),
    .Y(_09778_));
 sky130_fd_sc_hd__a32o_1 _16743_ (.A1(_09768_),
    .A2(_09777_),
    .A3(_09778_),
    .B1(_09769_),
    .B2(net5472),
    .X(_00525_));
 sky130_fd_sc_hd__xnor2_1 _16744_ (.A(net5722),
    .B(_09103_),
    .Y(_09779_));
 sky130_fd_sc_hd__a21bo_1 _16745_ (.A1(net5472),
    .A2(_09103_),
    .B1_N(_09778_),
    .X(_09780_));
 sky130_fd_sc_hd__xnor2_1 _16746_ (.A(_09779_),
    .B(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__a22o_1 _16747_ (.A1(net5722),
    .A2(_09769_),
    .B1(_09768_),
    .B2(_09781_),
    .X(_00526_));
 sky130_fd_sc_hd__o21a_1 _16748_ (.A1(net2968),
    .A2(_09103_),
    .B1(_09780_),
    .X(_09782_));
 sky130_fd_sc_hd__a21oi_1 _16749_ (.A1(net2968),
    .A2(_09103_),
    .B1(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__xnor2_1 _16750_ (.A(net5328),
    .B(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__nand2_1 _16751_ (.A(_09103_),
    .B(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__or2_1 _16752_ (.A(_09103_),
    .B(_09784_),
    .X(_09786_));
 sky130_fd_sc_hd__a32o_1 _16753_ (.A1(_09768_),
    .A2(_09785_),
    .A3(_09786_),
    .B1(_09769_),
    .B2(net5328),
    .X(_00527_));
 sky130_fd_sc_hd__nor3b_2 _16754_ (.A(net3976),
    .B(_04476_),
    .C_N(net3871),
    .Y(_09787_));
 sky130_fd_sc_hd__clkbuf_8 _16755_ (.A(net91),
    .X(_09788_));
 sky130_fd_sc_hd__nand2_1 _16756_ (.A(net4667),
    .B(net3822),
    .Y(_09789_));
 sky130_fd_sc_hd__or2_1 _16757_ (.A(net4667),
    .B(net3822),
    .X(_09790_));
 sky130_fd_sc_hd__and2b_1 _16758_ (.A_N(_08979_),
    .B(_08934_),
    .X(_09791_));
 sky130_fd_sc_hd__a21oi_1 _16759_ (.A1(_09791_),
    .A2(_08978_),
    .B1(net89),
    .Y(_09792_));
 sky130_fd_sc_hd__o21a_2 _16760_ (.A1(_09791_),
    .A2(_08978_),
    .B1(_09792_),
    .X(_09793_));
 sky130_fd_sc_hd__a31o_1 _16761_ (.A1(_09788_),
    .A2(net3805),
    .A3(_09790_),
    .B1(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__mux2_1 _16762_ (.A0(_09794_),
    .A1(net4667),
    .S(_09769_),
    .X(_09795_));
 sky130_fd_sc_hd__clkbuf_1 _16763_ (.A(_09795_),
    .X(_00528_));
 sky130_fd_sc_hd__or2_1 _16764_ (.A(net4506),
    .B(net4535),
    .X(_09796_));
 sky130_fd_sc_hd__nand2_1 _16765_ (.A(net4506),
    .B(net4535),
    .Y(_09797_));
 sky130_fd_sc_hd__nand2_1 _16766_ (.A(_09796_),
    .B(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__xnor2_1 _16767_ (.A(net3805),
    .B(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__o21ai_1 _16768_ (.A1(_08980_),
    .A2(_08982_),
    .B1(_06057_),
    .Y(_09800_));
 sky130_fd_sc_hd__a21o_1 _16769_ (.A1(_08980_),
    .A2(_08982_),
    .B1(_09800_),
    .X(_09801_));
 sky130_fd_sc_hd__o21ai_1 _16770_ (.A1(_06058_),
    .A2(_09799_),
    .B1(_09801_),
    .Y(_09802_));
 sky130_fd_sc_hd__mux2_1 _16771_ (.A0(_09802_),
    .A1(net4506),
    .S(_09769_),
    .X(_09803_));
 sky130_fd_sc_hd__clkbuf_1 _16772_ (.A(_09803_),
    .X(_00529_));
 sky130_fd_sc_hd__o21a_1 _16773_ (.A1(net3805),
    .A2(_09798_),
    .B1(_09797_),
    .X(_09804_));
 sky130_fd_sc_hd__nor2_1 _16774_ (.A(net3945),
    .B(net4353),
    .Y(_09805_));
 sky130_fd_sc_hd__nand2_1 _16775_ (.A(net3945),
    .B(net4353),
    .Y(_09806_));
 sky130_fd_sc_hd__or2b_1 _16776_ (.A(_09805_),
    .B_N(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__xnor2_1 _16777_ (.A(_09804_),
    .B(_09807_),
    .Y(_09808_));
 sky130_fd_sc_hd__buf_4 _16778_ (.A(_08103_),
    .X(_09809_));
 sky130_fd_sc_hd__nand2_1 _16779_ (.A(_09809_),
    .B(_09094_),
    .Y(_09810_));
 sky130_fd_sc_hd__o21ai_1 _16780_ (.A1(_06058_),
    .A2(_09808_),
    .B1(_09810_),
    .Y(_09811_));
 sky130_fd_sc_hd__mux2_1 _16781_ (.A0(_09811_),
    .A1(net3945),
    .S(_09769_),
    .X(_09812_));
 sky130_fd_sc_hd__clkbuf_1 _16782_ (.A(_09812_),
    .X(_00530_));
 sky130_fd_sc_hd__o21a_1 _16783_ (.A1(_09804_),
    .A2(_09805_),
    .B1(_09806_),
    .X(_09813_));
 sky130_fd_sc_hd__nor2_1 _16784_ (.A(net4569),
    .B(net4485),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2_1 _16785_ (.A(net4569),
    .B(net4485),
    .Y(_09815_));
 sky130_fd_sc_hd__or2b_1 _16786_ (.A(_09814_),
    .B_N(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__nor2_1 _16787_ (.A(_09813_),
    .B(_09816_),
    .Y(_09817_));
 sky130_fd_sc_hd__buf_4 _16788_ (.A(net4865),
    .X(_09818_));
 sky130_fd_sc_hd__a21o_1 _16789_ (.A1(_09813_),
    .A2(_09816_),
    .B1(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__nand2_1 _16790_ (.A(_09809_),
    .B(_09091_),
    .Y(_09820_));
 sky130_fd_sc_hd__o21ai_1 _16791_ (.A1(_09817_),
    .A2(_09819_),
    .B1(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__clkbuf_1 _16792_ (.A(net4648),
    .X(_09822_));
 sky130_fd_sc_hd__mux2_1 _16793_ (.A0(_09821_),
    .A1(net4569),
    .S(net4649),
    .X(_09823_));
 sky130_fd_sc_hd__clkbuf_1 _16794_ (.A(_09823_),
    .X(_00531_));
 sky130_fd_sc_hd__or2_1 _16795_ (.A(net4541),
    .B(net4630),
    .X(_09824_));
 sky130_fd_sc_hd__nand2_1 _16796_ (.A(net4541),
    .B(net4630),
    .Y(_09825_));
 sky130_fd_sc_hd__o21ai_2 _16797_ (.A1(_09813_),
    .A2(_09814_),
    .B1(_09815_),
    .Y(_09826_));
 sky130_fd_sc_hd__a21oi_1 _16798_ (.A1(_09824_),
    .A2(net4631),
    .B1(_09826_),
    .Y(_09827_));
 sky130_fd_sc_hd__a31o_1 _16799_ (.A1(_09826_),
    .A2(_09824_),
    .A3(net4631),
    .B1(_06057_),
    .X(_09828_));
 sky130_fd_sc_hd__nand2_1 _16800_ (.A(_09818_),
    .B(_09089_),
    .Y(_09829_));
 sky130_fd_sc_hd__o21ai_1 _16801_ (.A1(_09827_),
    .A2(_09828_),
    .B1(_09829_),
    .Y(_09830_));
 sky130_fd_sc_hd__mux2_1 _16802_ (.A0(_09830_),
    .A1(net4541),
    .S(net4649),
    .X(_09831_));
 sky130_fd_sc_hd__clkbuf_1 _16803_ (.A(_09831_),
    .X(_00532_));
 sky130_fd_sc_hd__a21boi_1 _16804_ (.A1(_09826_),
    .A2(_09824_),
    .B1_N(net4631),
    .Y(_09832_));
 sky130_fd_sc_hd__nor2_1 _16805_ (.A(net4547),
    .B(net4583),
    .Y(_09833_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(net4547),
    .B(net4583),
    .Y(_09834_));
 sky130_fd_sc_hd__or2b_1 _16807_ (.A(_09833_),
    .B_N(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__xnor2_1 _16808_ (.A(net4632),
    .B(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__nand2_1 _16809_ (.A(_09818_),
    .B(_09084_),
    .Y(_09837_));
 sky130_fd_sc_hd__o21ai_1 _16810_ (.A1(_06058_),
    .A2(_09836_),
    .B1(_09837_),
    .Y(_09838_));
 sky130_fd_sc_hd__mux2_1 _16811_ (.A0(_09838_),
    .A1(net4547),
    .S(net4649),
    .X(_09839_));
 sky130_fd_sc_hd__clkbuf_1 _16812_ (.A(_09839_),
    .X(_00533_));
 sky130_fd_sc_hd__o21a_1 _16813_ (.A1(net4632),
    .A2(_09833_),
    .B1(_09834_),
    .X(_09840_));
 sky130_fd_sc_hd__nor2_1 _16814_ (.A(net4508),
    .B(net4383),
    .Y(_09841_));
 sky130_fd_sc_hd__nand2_1 _16815_ (.A(net4508),
    .B(net4383),
    .Y(_09842_));
 sky130_fd_sc_hd__or2b_1 _16816_ (.A(_09841_),
    .B_N(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__nor2_1 _16817_ (.A(net4633),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__buf_4 _16818_ (.A(net4865),
    .X(_09845_));
 sky130_fd_sc_hd__a21o_1 _16819_ (.A1(net4633),
    .A2(_09843_),
    .B1(_09845_),
    .X(_09846_));
 sky130_fd_sc_hd__nand2_1 _16820_ (.A(_09818_),
    .B(_09209_),
    .Y(_09847_));
 sky130_fd_sc_hd__o21ai_1 _16821_ (.A1(net4634),
    .A2(_09846_),
    .B1(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__mux2_1 _16822_ (.A0(_09848_),
    .A1(net4508),
    .S(net4649),
    .X(_09849_));
 sky130_fd_sc_hd__clkbuf_1 _16823_ (.A(_09849_),
    .X(_00534_));
 sky130_fd_sc_hd__o21a_1 _16824_ (.A1(net4633),
    .A2(_09841_),
    .B1(_09842_),
    .X(_09850_));
 sky130_fd_sc_hd__nor2_1 _16825_ (.A(net4500),
    .B(net4789),
    .Y(_09851_));
 sky130_fd_sc_hd__nand2_1 _16826_ (.A(net4500),
    .B(net4789),
    .Y(_09852_));
 sky130_fd_sc_hd__or2b_1 _16827_ (.A(_09851_),
    .B_N(_09852_),
    .X(_09853_));
 sky130_fd_sc_hd__xnor2_1 _16828_ (.A(_09850_),
    .B(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__nand2_1 _16829_ (.A(_09818_),
    .B(_09326_),
    .Y(_09855_));
 sky130_fd_sc_hd__o21ai_1 _16830_ (.A1(_06058_),
    .A2(_09854_),
    .B1(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__mux2_1 _16831_ (.A0(_09856_),
    .A1(net4500),
    .S(net4649),
    .X(_09857_));
 sky130_fd_sc_hd__clkbuf_1 _16832_ (.A(_09857_),
    .X(_00535_));
 sky130_fd_sc_hd__o21a_1 _16833_ (.A1(_09850_),
    .A2(_09851_),
    .B1(_09852_),
    .X(_09858_));
 sky130_fd_sc_hd__nor2_1 _16834_ (.A(net3888),
    .B(net4776),
    .Y(_09859_));
 sky130_fd_sc_hd__nand2_1 _16835_ (.A(net3888),
    .B(net4776),
    .Y(_09860_));
 sky130_fd_sc_hd__or2b_1 _16836_ (.A(_09859_),
    .B_N(net3798),
    .X(_09861_));
 sky130_fd_sc_hd__nor2_1 _16837_ (.A(_09858_),
    .B(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__a21o_1 _16838_ (.A1(_09858_),
    .A2(_09861_),
    .B1(_09845_),
    .X(_09863_));
 sky130_fd_sc_hd__nand2_1 _16839_ (.A(_09818_),
    .B(_09450_),
    .Y(_09864_));
 sky130_fd_sc_hd__o21ai_1 _16840_ (.A1(_09862_),
    .A2(_09863_),
    .B1(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__mux2_1 _16841_ (.A0(_09865_),
    .A1(net3888),
    .S(net4649),
    .X(_09866_));
 sky130_fd_sc_hd__clkbuf_1 _16842_ (.A(_09866_),
    .X(_00536_));
 sky130_fd_sc_hd__or2_1 _16843_ (.A(net4665),
    .B(net4471),
    .X(_09867_));
 sky130_fd_sc_hd__nand2_2 _16844_ (.A(net4665),
    .B(net4471),
    .Y(_09868_));
 sky130_fd_sc_hd__o21ai_1 _16845_ (.A1(_09858_),
    .A2(_09859_),
    .B1(net3798),
    .Y(_09869_));
 sky130_fd_sc_hd__a21oi_1 _16846_ (.A1(_09867_),
    .A2(_09868_),
    .B1(net3799),
    .Y(_09870_));
 sky130_fd_sc_hd__a31o_1 _16847_ (.A1(net3799),
    .A2(_09867_),
    .A3(_09868_),
    .B1(_06057_),
    .X(_09871_));
 sky130_fd_sc_hd__nand2_1 _16848_ (.A(_09818_),
    .B(_09577_),
    .Y(_09872_));
 sky130_fd_sc_hd__o21ai_1 _16849_ (.A1(net3800),
    .A2(_09871_),
    .B1(_09872_),
    .Y(_09873_));
 sky130_fd_sc_hd__mux2_1 _16850_ (.A0(_09873_),
    .A1(net4665),
    .S(net4649),
    .X(_09874_));
 sky130_fd_sc_hd__clkbuf_1 _16851_ (.A(_09874_),
    .X(_00537_));
 sky130_fd_sc_hd__nand2_1 _16852_ (.A(net3799),
    .B(_09867_),
    .Y(_09875_));
 sky130_fd_sc_hd__and2_1 _16853_ (.A(net4581),
    .B(net4397),
    .X(_09876_));
 sky130_fd_sc_hd__nor2_1 _16854_ (.A(net4581),
    .B(net4397),
    .Y(_09877_));
 sky130_fd_sc_hd__a211oi_2 _16855_ (.A1(_09868_),
    .A2(_09875_),
    .B1(_09876_),
    .C1(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__o211a_1 _16856_ (.A1(_09877_),
    .A2(_09876_),
    .B1(_09875_),
    .C1(_09868_),
    .X(_09879_));
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(_09818_),
    .B(_09711_),
    .Y(_09880_));
 sky130_fd_sc_hd__o31ai_1 _16858_ (.A1(_09809_),
    .A2(_09878_),
    .A3(_09879_),
    .B1(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__mux2_1 _16859_ (.A0(_09881_),
    .A1(net4581),
    .S(net4649),
    .X(_09882_));
 sky130_fd_sc_hd__clkbuf_1 _16860_ (.A(_09882_),
    .X(_00538_));
 sky130_fd_sc_hd__or2_1 _16861_ (.A(net4669),
    .B(net4373),
    .X(_09883_));
 sky130_fd_sc_hd__nand2_1 _16862_ (.A(net4669),
    .B(net4373),
    .Y(_09884_));
 sky130_fd_sc_hd__a211o_1 _16863_ (.A1(_09883_),
    .A2(_09884_),
    .B1(_09876_),
    .C1(_09878_),
    .X(_09885_));
 sky130_fd_sc_hd__o211ai_1 _16864_ (.A1(_09876_),
    .A2(_09878_),
    .B1(_09883_),
    .C1(_09884_),
    .Y(_09886_));
 sky130_fd_sc_hd__nor2_1 _16865_ (.A(_09475_),
    .B(_09592_),
    .Y(_09887_));
 sky130_fd_sc_hd__a31o_1 _16866_ (.A1(_08611_),
    .A2(_09593_),
    .A3(net7818),
    .B1(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__or2b_1 _16867_ (.A(_09632_),
    .B_N(_09597_),
    .X(_09889_));
 sky130_fd_sc_hd__a21oi_1 _16868_ (.A1(_09611_),
    .A2(_09613_),
    .B1(_09609_),
    .Y(_09890_));
 sky130_fd_sc_hd__a21oi_2 _16869_ (.A1(_09630_),
    .A2(_09889_),
    .B1(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__and3_1 _16870_ (.A(_09630_),
    .B(_09889_),
    .C(_09890_),
    .X(_09892_));
 sky130_fd_sc_hd__nor2_1 _16871_ (.A(_09891_),
    .B(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__a21o_1 _16872_ (.A1(_09614_),
    .A2(_09628_),
    .B1(_09626_),
    .X(_09894_));
 sky130_fd_sc_hd__or2b_1 _16873_ (.A(_09652_),
    .B_N(_09634_),
    .X(_09895_));
 sky130_fd_sc_hd__nor2_1 _16874_ (.A(_08542_),
    .B(_09345_),
    .Y(_09896_));
 sky130_fd_sc_hd__nand2_1 _16875_ (.A(_09603_),
    .B(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__or2_1 _16876_ (.A(_09603_),
    .B(_09896_),
    .X(_09898_));
 sky130_fd_sc_hd__nand2_1 _16877_ (.A(_09897_),
    .B(_09898_),
    .Y(_09899_));
 sky130_fd_sc_hd__nor2_1 _16878_ (.A(_08543_),
    .B(_09472_),
    .Y(_09900_));
 sky130_fd_sc_hd__xor2_1 _16879_ (.A(_09899_),
    .B(_09900_),
    .X(_09901_));
 sky130_fd_sc_hd__a21oi_1 _16880_ (.A1(_09479_),
    .A2(_09603_),
    .B1(_09605_),
    .Y(_09902_));
 sky130_fd_sc_hd__nor2_1 _16881_ (.A(_09901_),
    .B(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__and2_1 _16882_ (.A(_09901_),
    .B(_09902_),
    .X(_09904_));
 sky130_fd_sc_hd__nor2_1 _16883_ (.A(_09903_),
    .B(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__and2_1 _16884_ (.A(_08127_),
    .B(net7818),
    .X(_09906_));
 sky130_fd_sc_hd__xor2_1 _16885_ (.A(_09905_),
    .B(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__a32o_1 _16886_ (.A1(_08864_),
    .A2(_09354_),
    .A3(_09618_),
    .B1(_09617_),
    .B2(_09506_),
    .X(_09908_));
 sky130_fd_sc_hd__and2_1 _16887_ (.A(_08204_),
    .B(_09354_),
    .X(_09909_));
 sky130_fd_sc_hd__or2_1 _16888_ (.A(_09617_),
    .B(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__nand2_1 _16889_ (.A(_09617_),
    .B(_09909_),
    .Y(_09911_));
 sky130_fd_sc_hd__and2_1 _16890_ (.A(_09910_),
    .B(_09911_),
    .X(_09912_));
 sky130_fd_sc_hd__nor2_1 _16891_ (.A(_08226_),
    .B(_09116_),
    .Y(_09913_));
 sky130_fd_sc_hd__xnor2_1 _16892_ (.A(_09912_),
    .B(_09913_),
    .Y(_09914_));
 sky130_fd_sc_hd__clkbuf_4 _16893_ (.A(_08383_),
    .X(_09915_));
 sky130_fd_sc_hd__or2b_1 _16894_ (.A(_09503_),
    .B_N(_09638_),
    .X(_09916_));
 sky130_fd_sc_hd__o31ai_1 _16895_ (.A1(_08338_),
    .A2(_09915_),
    .A3(_09636_),
    .B1(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__and2b_1 _16896_ (.A_N(_09914_),
    .B(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__and2b_1 _16897_ (.A_N(_09917_),
    .B(_09914_),
    .X(_09919_));
 sky130_fd_sc_hd__nor2_1 _16898_ (.A(_09918_),
    .B(_09919_),
    .Y(_09920_));
 sky130_fd_sc_hd__xnor2_1 _16899_ (.A(_09908_),
    .B(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__a21oi_1 _16900_ (.A1(_09615_),
    .A2(_09623_),
    .B1(_09621_),
    .Y(_09922_));
 sky130_fd_sc_hd__nor2_1 _16901_ (.A(_09921_),
    .B(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__and2_1 _16902_ (.A(_09921_),
    .B(_09922_),
    .X(_09924_));
 sky130_fd_sc_hd__nor2_1 _16903_ (.A(_09923_),
    .B(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__xnor2_1 _16904_ (.A(_09907_),
    .B(_09925_),
    .Y(_09926_));
 sky130_fd_sc_hd__a21o_1 _16905_ (.A1(_09650_),
    .A2(_09895_),
    .B1(_09926_),
    .X(_09927_));
 sky130_fd_sc_hd__nand3_1 _16906_ (.A(_09650_),
    .B(_09895_),
    .C(_09926_),
    .Y(_09928_));
 sky130_fd_sc_hd__nand2_1 _16907_ (.A(_09927_),
    .B(_09928_),
    .Y(_09929_));
 sky130_fd_sc_hd__xnor2_2 _16908_ (.A(_09894_),
    .B(_09929_),
    .Y(_09930_));
 sky130_fd_sc_hd__a21o_1 _16909_ (.A1(_09639_),
    .A2(_09647_),
    .B1(_09646_),
    .X(_09931_));
 sky130_fd_sc_hd__nand2_1 _16910_ (.A(_09656_),
    .B(_09661_),
    .Y(_09932_));
 sky130_fd_sc_hd__a21bo_1 _16911_ (.A1(_09655_),
    .A2(_09662_),
    .B1_N(_09932_),
    .X(_09933_));
 sky130_fd_sc_hd__o22ai_1 _16912_ (.A1(_08338_),
    .A2(_08374_),
    .B1(_08383_),
    .B2(_08142_),
    .Y(_09934_));
 sky130_fd_sc_hd__or2_1 _16913_ (.A(_08142_),
    .B(_08374_),
    .X(_09935_));
 sky130_fd_sc_hd__or3_1 _16914_ (.A(_08338_),
    .B(_08383_),
    .C(_09935_),
    .X(_09936_));
 sky130_fd_sc_hd__nand2_1 _16915_ (.A(_09934_),
    .B(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__or3_1 _16916_ (.A(_08661_),
    .B(_08616_),
    .C(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__o21ai_1 _16917_ (.A1(_08661_),
    .A2(_08616_),
    .B1(_09937_),
    .Y(_09939_));
 sky130_fd_sc_hd__and2_1 _16918_ (.A(_09938_),
    .B(_09939_),
    .X(_09940_));
 sky130_fd_sc_hd__nand2_1 _16919_ (.A(_09641_),
    .B(_09642_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_1 _16920_ (.A(_09640_),
    .B(_09643_),
    .Y(_09942_));
 sky130_fd_sc_hd__nor2_1 _16921_ (.A(_08326_),
    .B(_09025_),
    .Y(_09943_));
 sky130_fd_sc_hd__nor2_1 _16922_ (.A(_08309_),
    .B(_08411_),
    .Y(_09944_));
 sky130_fd_sc_hd__xor2_1 _16923_ (.A(_09943_),
    .B(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__nor2_1 _16924_ (.A(_09262_),
    .B(_08403_),
    .Y(_09946_));
 sky130_fd_sc_hd__xnor2_1 _16925_ (.A(_09945_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__a21oi_1 _16926_ (.A1(_09941_),
    .A2(_09942_),
    .B1(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__and3_1 _16927_ (.A(_09941_),
    .B(_09942_),
    .C(_09947_),
    .X(_09949_));
 sky130_fd_sc_hd__nor2_1 _16928_ (.A(_09948_),
    .B(_09949_),
    .Y(_09950_));
 sky130_fd_sc_hd__xnor2_1 _16929_ (.A(_09940_),
    .B(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__xor2_1 _16930_ (.A(_09933_),
    .B(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__xnor2_1 _16931_ (.A(_09931_),
    .B(_09952_),
    .Y(_09953_));
 sky130_fd_sc_hd__o21bai_2 _16932_ (.A1(_09657_),
    .A2(_09659_),
    .B1_N(_09658_),
    .Y(_09954_));
 sky130_fd_sc_hd__and2b_1 _16933_ (.A_N(_09668_),
    .B(_09669_),
    .X(_09955_));
 sky130_fd_sc_hd__a21o_1 _16934_ (.A1(_09665_),
    .A2(_09670_),
    .B1(_09955_),
    .X(_09956_));
 sky130_fd_sc_hd__or4_1 _16935_ (.A(_08880_),
    .B(_08391_),
    .C(_09170_),
    .D(_09292_),
    .X(_09957_));
 sky130_fd_sc_hd__a2bb2o_1 _16936_ (.A1_N(_08880_),
    .A2_N(_09292_),
    .B1(_08246_),
    .B2(_09288_),
    .X(_09958_));
 sky130_fd_sc_hd__nand2_1 _16937_ (.A(_09957_),
    .B(_09958_),
    .Y(_09959_));
 sky130_fd_sc_hd__nor2_1 _16938_ (.A(_09272_),
    .B(_09165_),
    .Y(_09960_));
 sky130_fd_sc_hd__xnor2_1 _16939_ (.A(_09959_),
    .B(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__xor2_1 _16940_ (.A(_09956_),
    .B(_09961_),
    .X(_09962_));
 sky130_fd_sc_hd__xor2_1 _16941_ (.A(_09954_),
    .B(_09962_),
    .X(_09963_));
 sky130_fd_sc_hd__nor2_1 _16942_ (.A(_09537_),
    .B(_09664_),
    .Y(_09964_));
 sky130_fd_sc_hd__a21oi_1 _16943_ (.A1(_09666_),
    .A2(_09667_),
    .B1(_08401_),
    .Y(_09965_));
 sky130_fd_sc_hd__a21oi_1 _16944_ (.A1(_09540_),
    .A2(_09541_),
    .B1(_08916_),
    .Y(_09966_));
 sky130_fd_sc_hd__xnor2_1 _16945_ (.A(_09965_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__xnor2_1 _16946_ (.A(_09964_),
    .B(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__and2_1 _16947_ (.A(net4622),
    .B(_06123_),
    .X(_09969_));
 sky130_fd_sc_hd__a21oi_4 _16948_ (.A1(_08181_),
    .A2(_09673_),
    .B1(_09969_),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_1 _16949_ (.A(_08474_),
    .B(_08494_),
    .Y(_09971_));
 sky130_fd_sc_hd__o211a_1 _16950_ (.A1(net4877),
    .A2(_08494_),
    .B1(_09673_),
    .C1(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__or3b_1 _16951_ (.A(_08905_),
    .B(_09970_),
    .C_N(_09972_),
    .X(_09973_));
 sky130_fd_sc_hd__a21o_1 _16952_ (.A1(_09676_),
    .A2(_09546_),
    .B1(_06124_),
    .X(_09974_));
 sky130_fd_sc_hd__nand2_1 _16953_ (.A(net4388),
    .B(_06124_),
    .Y(_09975_));
 sky130_fd_sc_hd__and2_2 _16954_ (.A(_09974_),
    .B(_09975_),
    .X(_09976_));
 sky130_fd_sc_hd__o21bai_1 _16955_ (.A1(_08905_),
    .A2(_09976_),
    .B1_N(_09972_),
    .Y(_09977_));
 sky130_fd_sc_hd__a21bo_1 _16956_ (.A1(_09674_),
    .A2(_09677_),
    .B1_N(_09675_),
    .X(_09978_));
 sky130_fd_sc_hd__nand3_2 _16957_ (.A(_09973_),
    .B(_09977_),
    .C(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__a21o_1 _16958_ (.A1(_09973_),
    .A2(_09977_),
    .B1(_09978_),
    .X(_09980_));
 sky130_fd_sc_hd__nand3_1 _16959_ (.A(_09968_),
    .B(_09979_),
    .C(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__a21o_1 _16960_ (.A1(_09979_),
    .A2(_09980_),
    .B1(_09968_),
    .X(_09982_));
 sky130_fd_sc_hd__a21bo_1 _16961_ (.A1(_09671_),
    .A2(_09683_),
    .B1_N(_09682_),
    .X(_09983_));
 sky130_fd_sc_hd__nand3_1 _16962_ (.A(_09981_),
    .B(_09982_),
    .C(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__a21o_1 _16963_ (.A1(_09981_),
    .A2(_09982_),
    .B1(_09983_),
    .X(_09985_));
 sky130_fd_sc_hd__and3_1 _16964_ (.A(_09963_),
    .B(_09984_),
    .C(_09985_),
    .X(_09986_));
 sky130_fd_sc_hd__a21oi_1 _16965_ (.A1(_09984_),
    .A2(_09985_),
    .B1(_09963_),
    .Y(_09987_));
 sky130_fd_sc_hd__or2_2 _16966_ (.A(_09986_),
    .B(_09987_),
    .X(_09988_));
 sky130_fd_sc_hd__a21boi_2 _16967_ (.A1(_09663_),
    .A2(_09689_),
    .B1_N(_09688_),
    .Y(_09989_));
 sky130_fd_sc_hd__xor2_2 _16968_ (.A(_09988_),
    .B(_09989_),
    .X(_09990_));
 sky130_fd_sc_hd__xnor2_1 _16969_ (.A(_09953_),
    .B(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__nor2_1 _16970_ (.A(_09692_),
    .B(_09694_),
    .Y(_09992_));
 sky130_fd_sc_hd__a21oi_2 _16971_ (.A1(_09653_),
    .A2(_09695_),
    .B1(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__nor2_1 _16972_ (.A(_09991_),
    .B(_09993_),
    .Y(_09994_));
 sky130_fd_sc_hd__and2_1 _16973_ (.A(_09991_),
    .B(_09993_),
    .X(_09995_));
 sky130_fd_sc_hd__nor2_2 _16974_ (.A(_09994_),
    .B(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__xnor2_2 _16975_ (.A(_09930_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__a21o_1 _16976_ (.A1(_09633_),
    .A2(_09700_),
    .B1(_09698_),
    .X(_09998_));
 sky130_fd_sc_hd__xnor2_2 _16977_ (.A(_09997_),
    .B(_09998_),
    .Y(_09999_));
 sky130_fd_sc_hd__xnor2_1 _16978_ (.A(_09893_),
    .B(_09999_),
    .Y(_10000_));
 sky130_fd_sc_hd__o2bb2a_1 _16979_ (.A1_N(_09596_),
    .A2_N(_09703_),
    .B1(_09702_),
    .B2(_09701_),
    .X(_10001_));
 sky130_fd_sc_hd__xor2_1 _16980_ (.A(_10000_),
    .B(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__xor2_1 _16981_ (.A(_09888_),
    .B(_10002_),
    .X(_10003_));
 sky130_fd_sc_hd__nand2_2 _16982_ (.A(_09707_),
    .B(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__or2_1 _16983_ (.A(_09707_),
    .B(_10003_),
    .X(_10005_));
 sky130_fd_sc_hd__nand2_4 _16984_ (.A(_10004_),
    .B(_10005_),
    .Y(_10006_));
 sky130_fd_sc_hd__a21o_1 _16985_ (.A1(_09590_),
    .A2(_09588_),
    .B1(_09709_),
    .X(_10007_));
 sky130_fd_sc_hd__o31a_4 _16986_ (.A1(_09460_),
    .A2(_09587_),
    .A3(_09710_),
    .B1(_10007_),
    .X(_10008_));
 sky130_fd_sc_hd__xor2_4 _16987_ (.A(_10006_),
    .B(_10008_),
    .X(_10009_));
 sky130_fd_sc_hd__and2_1 _16988_ (.A(_08103_),
    .B(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__a31o_1 _16989_ (.A1(_09788_),
    .A2(net8375),
    .A3(net8383),
    .B1(_10010_),
    .X(_10011_));
 sky130_fd_sc_hd__mux2_1 _16990_ (.A0(_10011_),
    .A1(net4669),
    .S(net4649),
    .X(_10012_));
 sky130_fd_sc_hd__clkbuf_1 _16991_ (.A(_10012_),
    .X(_00539_));
 sky130_fd_sc_hd__and2_1 _16992_ (.A(net4589),
    .B(net4483),
    .X(_10013_));
 sky130_fd_sc_hd__nor2_1 _16993_ (.A(net4589),
    .B(net4483),
    .Y(_10014_));
 sky130_fd_sc_hd__a211o_1 _16994_ (.A1(_09884_),
    .A2(net8383),
    .B1(_10013_),
    .C1(_10014_),
    .X(_10015_));
 sky130_fd_sc_hd__o211ai_1 _16995_ (.A1(_10013_),
    .A2(_10014_),
    .B1(_09884_),
    .C1(net8383),
    .Y(_10016_));
 sky130_fd_sc_hd__or2_1 _16996_ (.A(_10000_),
    .B(_10001_),
    .X(_10017_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(_09888_),
    .B(_10002_),
    .Y(_10018_));
 sky130_fd_sc_hd__or2b_1 _16998_ (.A(_09929_),
    .B_N(_09894_),
    .X(_10019_));
 sky130_fd_sc_hd__a21oi_2 _16999_ (.A1(_09905_),
    .A2(_09906_),
    .B1(_09903_),
    .Y(_10020_));
 sky130_fd_sc_hd__a21oi_4 _17000_ (.A1(_09927_),
    .A2(_10019_),
    .B1(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__and3_1 _17001_ (.A(_09927_),
    .B(_10019_),
    .C(_10020_),
    .X(_10022_));
 sky130_fd_sc_hd__nor2_2 _17002_ (.A(_10021_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__a21o_1 _17003_ (.A1(_09907_),
    .A2(_09925_),
    .B1(_09923_),
    .X(_10024_));
 sky130_fd_sc_hd__or2b_1 _17004_ (.A(_09951_),
    .B_N(_09933_),
    .X(_10025_));
 sky130_fd_sc_hd__or2b_1 _17005_ (.A(_09952_),
    .B_N(_09931_),
    .X(_10026_));
 sky130_fd_sc_hd__nor2_1 _17006_ (.A(_06124_),
    .B(net4913),
    .Y(_10027_));
 sky130_fd_sc_hd__nor2_1 _17007_ (.A(_08226_),
    .B(_09225_),
    .Y(_10028_));
 sky130_fd_sc_hd__a21o_1 _17008_ (.A1(_09133_),
    .A2(net4914),
    .B1(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__nor2_1 _17009_ (.A(_08226_),
    .B(_09345_),
    .Y(_10030_));
 sky130_fd_sc_hd__nand2_1 _17010_ (.A(_09603_),
    .B(_10030_),
    .Y(_10031_));
 sky130_fd_sc_hd__nand2_1 _17011_ (.A(_10029_),
    .B(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__or2_1 _17012_ (.A(_08542_),
    .B(_09472_),
    .X(_10033_));
 sky130_fd_sc_hd__xnor2_1 _17013_ (.A(_10032_),
    .B(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__o31a_1 _17014_ (.A1(_08543_),
    .A2(_09472_),
    .A3(_09899_),
    .B1(_09897_),
    .X(_10035_));
 sky130_fd_sc_hd__xnor2_1 _17015_ (.A(_10034_),
    .B(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__and2_1 _17016_ (.A(_08543_),
    .B(net7818),
    .X(_10037_));
 sky130_fd_sc_hd__xnor2_1 _17017_ (.A(_10036_),
    .B(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__a21bo_1 _17018_ (.A1(_09912_),
    .A2(_09913_),
    .B1_N(_09911_),
    .X(_10039_));
 sky130_fd_sc_hd__nand2_1 _17019_ (.A(_08167_),
    .B(_09351_),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_1 _17020_ (.A(_09373_),
    .B(_09354_),
    .Y(_10041_));
 sky130_fd_sc_hd__nor2_1 _17021_ (.A(_08661_),
    .B(_09062_),
    .Y(_10042_));
 sky130_fd_sc_hd__a22o_1 _17022_ (.A1(_10040_),
    .A2(_10041_),
    .B1(_10042_),
    .B2(_09617_),
    .X(_10043_));
 sky130_fd_sc_hd__nand2_1 _17023_ (.A(_09249_),
    .B(_09600_),
    .Y(_10044_));
 sky130_fd_sc_hd__xnor2_1 _17024_ (.A(_10043_),
    .B(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__a21oi_1 _17025_ (.A1(_09936_),
    .A2(_09938_),
    .B1(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__and3_1 _17026_ (.A(_09936_),
    .B(_09938_),
    .C(_10045_),
    .X(_10047_));
 sky130_fd_sc_hd__nor2_1 _17027_ (.A(_10046_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__xnor2_1 _17028_ (.A(_10039_),
    .B(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__a21oi_1 _17029_ (.A1(_09908_),
    .A2(_09920_),
    .B1(_09918_),
    .Y(_10050_));
 sky130_fd_sc_hd__nor2_1 _17030_ (.A(_10049_),
    .B(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__and2_1 _17031_ (.A(_10049_),
    .B(_10050_),
    .X(_10052_));
 sky130_fd_sc_hd__nor2_1 _17032_ (.A(_10051_),
    .B(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__xnor2_1 _17033_ (.A(_10038_),
    .B(_10053_),
    .Y(_10054_));
 sky130_fd_sc_hd__a21o_1 _17034_ (.A1(_10025_),
    .A2(_10026_),
    .B1(_10054_),
    .X(_10055_));
 sky130_fd_sc_hd__nand3_1 _17035_ (.A(_10025_),
    .B(_10026_),
    .C(_10054_),
    .Y(_10056_));
 sky130_fd_sc_hd__nand2_1 _17036_ (.A(_10055_),
    .B(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__xnor2_2 _17037_ (.A(_10024_),
    .B(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__a21o_1 _17038_ (.A1(_09940_),
    .A2(_09950_),
    .B1(_09948_),
    .X(_10059_));
 sky130_fd_sc_hd__nand2_1 _17039_ (.A(_09956_),
    .B(_09961_),
    .Y(_10060_));
 sky130_fd_sc_hd__nand2_1 _17040_ (.A(_09954_),
    .B(_09962_),
    .Y(_10061_));
 sky130_fd_sc_hd__buf_2 _17041_ (.A(net4918),
    .X(_10062_));
 sky130_fd_sc_hd__nor2_1 _17042_ (.A(_10062_),
    .B(_08413_),
    .Y(_10063_));
 sky130_fd_sc_hd__xor2_1 _17043_ (.A(_09935_),
    .B(_10063_),
    .X(_10064_));
 sky130_fd_sc_hd__or3_1 _17044_ (.A(_09915_),
    .B(_08616_),
    .C(_10064_),
    .X(_10065_));
 sky130_fd_sc_hd__o21ai_1 _17045_ (.A1(_09915_),
    .A2(_08616_),
    .B1(_10064_),
    .Y(_10066_));
 sky130_fd_sc_hd__and2_1 _17046_ (.A(_10065_),
    .B(_10066_),
    .X(_10067_));
 sky130_fd_sc_hd__nor2_1 _17047_ (.A(_08309_),
    .B(_09025_),
    .Y(_10068_));
 sky130_fd_sc_hd__nor2_1 _17048_ (.A(_08308_),
    .B(_09165_),
    .Y(_10069_));
 sky130_fd_sc_hd__xor2_1 _17049_ (.A(_10068_),
    .B(_10069_),
    .X(_10070_));
 sky130_fd_sc_hd__nor2_1 _17050_ (.A(_09262_),
    .B(_08411_),
    .Y(_10071_));
 sky130_fd_sc_hd__xnor2_1 _17051_ (.A(_10070_),
    .B(_10071_),
    .Y(_10072_));
 sky130_fd_sc_hd__nand2_1 _17052_ (.A(_09943_),
    .B(_09944_),
    .Y(_10073_));
 sky130_fd_sc_hd__a21boi_1 _17053_ (.A1(_09945_),
    .A2(_09946_),
    .B1_N(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__nor2_1 _17054_ (.A(_10072_),
    .B(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__nand2_1 _17055_ (.A(_10072_),
    .B(_10074_),
    .Y(_10076_));
 sky130_fd_sc_hd__and2b_1 _17056_ (.A_N(_10075_),
    .B(_10076_),
    .X(_10077_));
 sky130_fd_sc_hd__xnor2_1 _17057_ (.A(_10067_),
    .B(_10077_),
    .Y(_10078_));
 sky130_fd_sc_hd__a21o_1 _17058_ (.A1(_10060_),
    .A2(_10061_),
    .B1(_10078_),
    .X(_10079_));
 sky130_fd_sc_hd__nand3_1 _17059_ (.A(_10060_),
    .B(_10061_),
    .C(_10078_),
    .Y(_10080_));
 sky130_fd_sc_hd__nand2_1 _17060_ (.A(_10079_),
    .B(_10080_),
    .Y(_10081_));
 sky130_fd_sc_hd__xnor2_1 _17061_ (.A(_10059_),
    .B(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__a21bo_1 _17062_ (.A1(_09958_),
    .A2(_09960_),
    .B1_N(_09957_),
    .X(_10083_));
 sky130_fd_sc_hd__and2_1 _17063_ (.A(_09965_),
    .B(_09966_),
    .X(_10084_));
 sky130_fd_sc_hd__nor3_1 _17064_ (.A(_09537_),
    .B(_09664_),
    .C(_09967_),
    .Y(_10085_));
 sky130_fd_sc_hd__or4_1 _17065_ (.A(_08880_),
    .B(_08391_),
    .C(_09292_),
    .D(_09411_),
    .X(_10086_));
 sky130_fd_sc_hd__o22ai_1 _17066_ (.A1(_08391_),
    .A2(_09292_),
    .B1(_09411_),
    .B2(_08880_),
    .Y(_10087_));
 sky130_fd_sc_hd__nand2_1 _17067_ (.A(_10086_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__or2_1 _17068_ (.A(_08509_),
    .B(_09170_),
    .X(_10089_));
 sky130_fd_sc_hd__xor2_1 _17069_ (.A(_10088_),
    .B(_10089_),
    .X(_10090_));
 sky130_fd_sc_hd__o21a_1 _17070_ (.A1(_10084_),
    .A2(_10085_),
    .B1(_10090_),
    .X(_10091_));
 sky130_fd_sc_hd__or3_1 _17071_ (.A(_10084_),
    .B(_10085_),
    .C(_10090_),
    .X(_10092_));
 sky130_fd_sc_hd__or2b_1 _17072_ (.A(_10091_),
    .B_N(_10092_),
    .X(_10093_));
 sky130_fd_sc_hd__xnor2_2 _17073_ (.A(_10083_),
    .B(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__and2_1 _17074_ (.A(_09540_),
    .B(_09541_),
    .X(_10095_));
 sky130_fd_sc_hd__buf_4 _17075_ (.A(_10095_),
    .X(_10096_));
 sky130_fd_sc_hd__nor2_1 _17076_ (.A(_09537_),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__a21o_1 _17077_ (.A1(_09666_),
    .A2(_09667_),
    .B1(_08402_),
    .X(_10098_));
 sky130_fd_sc_hd__a21oi_1 _17078_ (.A1(_09974_),
    .A2(_09975_),
    .B1(_08948_),
    .Y(_10099_));
 sky130_fd_sc_hd__xnor2_1 _17079_ (.A(_10098_),
    .B(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__xor2_1 _17080_ (.A(_10097_),
    .B(_10100_),
    .X(_10101_));
 sky130_fd_sc_hd__and2_1 _17081_ (.A(_09673_),
    .B(_09971_),
    .X(_10102_));
 sky130_fd_sc_hd__nor2_1 _17082_ (.A(_08905_),
    .B(_09970_),
    .Y(_10103_));
 sky130_fd_sc_hd__nand2_1 _17083_ (.A(_08573_),
    .B(_09673_),
    .Y(_10104_));
 sky130_fd_sc_hd__or4_4 _17084_ (.A(_08905_),
    .B(net4877),
    .C(_10104_),
    .D(_09970_),
    .X(_10105_));
 sky130_fd_sc_hd__o21a_2 _17085_ (.A1(_10102_),
    .A2(_10103_),
    .B1(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__xnor2_1 _17086_ (.A(_10101_),
    .B(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__a21oi_1 _17087_ (.A1(_09979_),
    .A2(_09981_),
    .B1(_10107_),
    .Y(_10108_));
 sky130_fd_sc_hd__and3_1 _17088_ (.A(_09979_),
    .B(_09981_),
    .C(_10107_),
    .X(_10109_));
 sky130_fd_sc_hd__nor2_1 _17089_ (.A(_10108_),
    .B(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__xnor2_2 _17090_ (.A(_10094_),
    .B(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__a21boi_2 _17091_ (.A1(_09963_),
    .A2(_09985_),
    .B1_N(_09984_),
    .Y(_10112_));
 sky130_fd_sc_hd__xor2_2 _17092_ (.A(_10111_),
    .B(_10112_),
    .X(_10113_));
 sky130_fd_sc_hd__xnor2_1 _17093_ (.A(_10082_),
    .B(_10113_),
    .Y(_10114_));
 sky130_fd_sc_hd__nor2_1 _17094_ (.A(_09988_),
    .B(_09989_),
    .Y(_10115_));
 sky130_fd_sc_hd__a21oi_1 _17095_ (.A1(_09953_),
    .A2(_09990_),
    .B1(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__nor2_1 _17096_ (.A(_10114_),
    .B(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__nand2_1 _17097_ (.A(_10114_),
    .B(_10116_),
    .Y(_10118_));
 sky130_fd_sc_hd__and2b_1 _17098_ (.A_N(_10117_),
    .B(_10118_),
    .X(_10119_));
 sky130_fd_sc_hd__xnor2_2 _17099_ (.A(_10058_),
    .B(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__a21oi_2 _17100_ (.A1(_09930_),
    .A2(_09996_),
    .B1(_09994_),
    .Y(_10121_));
 sky130_fd_sc_hd__xor2_2 _17101_ (.A(_10120_),
    .B(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__xnor2_2 _17102_ (.A(_10023_),
    .B(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__or2b_1 _17103_ (.A(_09997_),
    .B_N(_09998_),
    .X(_10124_));
 sky130_fd_sc_hd__a21boi_2 _17104_ (.A1(_09893_),
    .A2(_09999_),
    .B1_N(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__xor2_2 _17105_ (.A(_10123_),
    .B(_10125_),
    .X(_10126_));
 sky130_fd_sc_hd__xnor2_1 _17106_ (.A(_09891_),
    .B(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__a21oi_1 _17107_ (.A1(_10017_),
    .A2(_10018_),
    .B1(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__and3_1 _17108_ (.A(_10017_),
    .B(_10018_),
    .C(_10127_),
    .X(_10129_));
 sky130_fd_sc_hd__or2_2 _17109_ (.A(_10128_),
    .B(_10129_),
    .X(_10130_));
 sky130_fd_sc_hd__o21ai_2 _17110_ (.A1(_10006_),
    .A2(_10008_),
    .B1(_10004_),
    .Y(_10131_));
 sky130_fd_sc_hd__xnor2_4 _17111_ (.A(_10130_),
    .B(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__and2_1 _17112_ (.A(_08103_),
    .B(_10132_),
    .X(_10133_));
 sky130_fd_sc_hd__a31o_1 _17113_ (.A1(_09788_),
    .A2(_10015_),
    .A3(_10016_),
    .B1(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__mux2_1 _17114_ (.A0(_10134_),
    .A1(net4589),
    .S(net4649),
    .X(_10135_));
 sky130_fd_sc_hd__clkbuf_1 _17115_ (.A(_10135_),
    .X(_00540_));
 sky130_fd_sc_hd__nand2_1 _17116_ (.A(net4657),
    .B(net4401),
    .Y(_10136_));
 sky130_fd_sc_hd__or2_1 _17117_ (.A(net4657),
    .B(net4401),
    .X(_10137_));
 sky130_fd_sc_hd__inv_2 _17118_ (.A(_10015_),
    .Y(_10138_));
 sky130_fd_sc_hd__a211o_1 _17119_ (.A1(_10136_),
    .A2(_10137_),
    .B1(_10013_),
    .C1(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__o211ai_2 _17120_ (.A1(_10013_),
    .A2(_10138_),
    .B1(_10136_),
    .C1(_10137_),
    .Y(_10140_));
 sky130_fd_sc_hd__or2b_1 _17121_ (.A(_10057_),
    .B_N(_10024_),
    .X(_10141_));
 sky130_fd_sc_hd__or2b_1 _17122_ (.A(_10036_),
    .B_N(_10037_),
    .X(_10142_));
 sky130_fd_sc_hd__o21a_1 _17123_ (.A1(_10034_),
    .A2(_10035_),
    .B1(_10142_),
    .X(_10143_));
 sky130_fd_sc_hd__a21oi_2 _17124_ (.A1(_10055_),
    .A2(_10141_),
    .B1(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__and3_1 _17125_ (.A(_10055_),
    .B(_10141_),
    .C(_10143_),
    .X(_10145_));
 sky130_fd_sc_hd__nor2_2 _17126_ (.A(_10144_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__a21o_1 _17127_ (.A1(_10038_),
    .A2(_10053_),
    .B1(_10051_),
    .X(_10147_));
 sky130_fd_sc_hd__or2b_1 _17128_ (.A(_10081_),
    .B_N(_10059_),
    .X(_10148_));
 sky130_fd_sc_hd__and2_1 _17129_ (.A(_09249_),
    .B(net4909),
    .X(_10149_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(_09249_),
    .B(net4914),
    .Y(_10150_));
 sky130_fd_sc_hd__inv_2 _17131_ (.A(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__nand2_1 _17132_ (.A(_10028_),
    .B(_10151_),
    .Y(_10152_));
 sky130_fd_sc_hd__o21a_1 _17133_ (.A1(_10030_),
    .A2(_10149_),
    .B1(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__and2b_1 _17134_ (.A_N(_09472_),
    .B(_09133_),
    .X(_10154_));
 sky130_fd_sc_hd__xnor2_1 _17135_ (.A(_10153_),
    .B(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__o31a_1 _17136_ (.A1(_08542_),
    .A2(_09612_),
    .A3(_10032_),
    .B1(_10031_),
    .X(_10156_));
 sky130_fd_sc_hd__nor2_1 _17137_ (.A(_10155_),
    .B(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__and2_1 _17138_ (.A(_10155_),
    .B(_10156_),
    .X(_10158_));
 sky130_fd_sc_hd__nor2_1 _17139_ (.A(_10157_),
    .B(_10158_),
    .Y(_10159_));
 sky130_fd_sc_hd__and2_1 _17140_ (.A(_08542_),
    .B(net7818),
    .X(_10160_));
 sky130_fd_sc_hd__xor2_1 _17141_ (.A(_10159_),
    .B(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__o2bb2ai_1 _17142_ (.A1_N(_09617_),
    .A2_N(_10042_),
    .B1(_10043_),
    .B2(_10044_),
    .Y(_10162_));
 sky130_fd_sc_hd__clkbuf_4 _17143_ (.A(_08413_),
    .X(_10163_));
 sky130_fd_sc_hd__or3_1 _17144_ (.A(_10062_),
    .B(_10163_),
    .C(_09935_),
    .X(_10164_));
 sky130_fd_sc_hd__nor2_1 _17145_ (.A(_08383_),
    .B(_08614_),
    .Y(_10165_));
 sky130_fd_sc_hd__or3_1 _17146_ (.A(_08383_),
    .B(_09062_),
    .C(_10040_),
    .X(_10166_));
 sky130_fd_sc_hd__o21a_1 _17147_ (.A1(_10042_),
    .A2(_10165_),
    .B1(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__and2_1 _17148_ (.A(_09373_),
    .B(_09600_),
    .X(_10168_));
 sky130_fd_sc_hd__xnor2_1 _17149_ (.A(_10167_),
    .B(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__a21oi_1 _17150_ (.A1(_10164_),
    .A2(_10065_),
    .B1(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__and3_1 _17151_ (.A(_10164_),
    .B(_10065_),
    .C(_10169_),
    .X(_10171_));
 sky130_fd_sc_hd__nor2_1 _17152_ (.A(_10170_),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__xnor2_1 _17153_ (.A(_10162_),
    .B(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__a21oi_1 _17154_ (.A1(_10039_),
    .A2(_10048_),
    .B1(_10046_),
    .Y(_10174_));
 sky130_fd_sc_hd__nor2_1 _17155_ (.A(_10173_),
    .B(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__and2_1 _17156_ (.A(_10173_),
    .B(_10174_),
    .X(_10176_));
 sky130_fd_sc_hd__nor2_1 _17157_ (.A(_10175_),
    .B(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__xnor2_1 _17158_ (.A(_10161_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__a21o_1 _17159_ (.A1(_10079_),
    .A2(_10148_),
    .B1(_10178_),
    .X(_10179_));
 sky130_fd_sc_hd__nand3_1 _17160_ (.A(_10079_),
    .B(_10148_),
    .C(_10178_),
    .Y(_10180_));
 sky130_fd_sc_hd__nand2_1 _17161_ (.A(_10179_),
    .B(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__xnor2_2 _17162_ (.A(_10147_),
    .B(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__a21o_1 _17163_ (.A1(_10067_),
    .A2(_10076_),
    .B1(_10075_),
    .X(_10183_));
 sky130_fd_sc_hd__a21o_1 _17164_ (.A1(_10083_),
    .A2(_10092_),
    .B1(_10091_),
    .X(_10184_));
 sky130_fd_sc_hd__a2bb2o_1 _17165_ (.A1_N(_08338_),
    .A2_N(_08472_),
    .B1(_09135_),
    .B2(_08366_),
    .X(_10185_));
 sky130_fd_sc_hd__nand2_1 _17166_ (.A(_08408_),
    .B(_08409_),
    .Y(_10186_));
 sky130_fd_sc_hd__nor2_1 _17167_ (.A(_08140_),
    .B(_10186_),
    .Y(_10187_));
 sky130_fd_sc_hd__nand2_1 _17168_ (.A(_10063_),
    .B(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__and2_1 _17169_ (.A(_10185_),
    .B(_10188_),
    .X(_10189_));
 sky130_fd_sc_hd__clkbuf_4 _17170_ (.A(_08374_),
    .X(_10190_));
 sky130_fd_sc_hd__nor2_1 _17171_ (.A(_10190_),
    .B(_08616_),
    .Y(_10191_));
 sky130_fd_sc_hd__xnor2_1 _17172_ (.A(_10189_),
    .B(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__or2_1 _17173_ (.A(_08309_),
    .B(_09165_),
    .X(_10193_));
 sky130_fd_sc_hd__nor2_1 _17174_ (.A(_08326_),
    .B(_09170_),
    .Y(_10194_));
 sky130_fd_sc_hd__xnor2_1 _17175_ (.A(_10193_),
    .B(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__nor2_1 _17176_ (.A(_09262_),
    .B(_09025_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand2_1 _17177_ (.A(_10195_),
    .B(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__or2_1 _17178_ (.A(_10195_),
    .B(_10196_),
    .X(_10198_));
 sky130_fd_sc_hd__nand2_1 _17179_ (.A(_10197_),
    .B(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__and2_1 _17180_ (.A(_10070_),
    .B(_10071_),
    .X(_10200_));
 sky130_fd_sc_hd__a21oi_2 _17181_ (.A1(_10068_),
    .A2(_10069_),
    .B1(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__xor2_1 _17182_ (.A(_10199_),
    .B(_10201_),
    .X(_10202_));
 sky130_fd_sc_hd__xnor2_1 _17183_ (.A(_10192_),
    .B(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__nand2_1 _17184_ (.A(_10184_),
    .B(_10203_),
    .Y(_10204_));
 sky130_fd_sc_hd__or2_1 _17185_ (.A(_10184_),
    .B(_10203_),
    .X(_10205_));
 sky130_fd_sc_hd__nand2_1 _17186_ (.A(_10204_),
    .B(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__xnor2_1 _17187_ (.A(_10183_),
    .B(_10206_),
    .Y(_10207_));
 sky130_fd_sc_hd__o21ai_2 _17188_ (.A1(_10088_),
    .A2(_10089_),
    .B1(_10086_),
    .Y(_10208_));
 sky130_fd_sc_hd__and2b_1 _17189_ (.A_N(_10098_),
    .B(_10099_),
    .X(_10209_));
 sky130_fd_sc_hd__a21o_1 _17190_ (.A1(_10097_),
    .A2(_10100_),
    .B1(_10209_),
    .X(_10210_));
 sky130_fd_sc_hd__clkbuf_4 _17191_ (.A(_08391_),
    .X(_10211_));
 sky130_fd_sc_hd__or4_2 _17192_ (.A(_08880_),
    .B(_10211_),
    .C(_09411_),
    .D(_10096_),
    .X(_10212_));
 sky130_fd_sc_hd__o22ai_2 _17193_ (.A1(_10211_),
    .A2(_09664_),
    .B1(_10096_),
    .B2(_08918_),
    .Y(_10213_));
 sky130_fd_sc_hd__nand2_1 _17194_ (.A(_10212_),
    .B(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__nor2_1 _17195_ (.A(_09272_),
    .B(_09403_),
    .Y(_10215_));
 sky130_fd_sc_hd__xnor2_2 _17196_ (.A(_10214_),
    .B(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__xnor2_2 _17197_ (.A(_10210_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__xnor2_2 _17198_ (.A(_10208_),
    .B(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__and2_1 _17199_ (.A(_09666_),
    .B(_09667_),
    .X(_10219_));
 sky130_fd_sc_hd__clkbuf_4 _17200_ (.A(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__nor2_1 _17201_ (.A(_09537_),
    .B(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__o22ai_1 _17202_ (.A1(_08948_),
    .A2(_09970_),
    .B1(_09976_),
    .B2(_08916_),
    .Y(_10222_));
 sky130_fd_sc_hd__or4_1 _17203_ (.A(_08948_),
    .B(_08916_),
    .C(_09970_),
    .D(_09976_),
    .X(_10223_));
 sky130_fd_sc_hd__nand3_1 _17204_ (.A(_10221_),
    .B(_10222_),
    .C(_10223_),
    .Y(_10224_));
 sky130_fd_sc_hd__a21o_1 _17205_ (.A1(_10222_),
    .A2(_10223_),
    .B1(_10221_),
    .X(_10225_));
 sky130_fd_sc_hd__nand3_1 _17206_ (.A(_10106_),
    .B(_10224_),
    .C(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__a21o_1 _17207_ (.A1(_10224_),
    .A2(_10225_),
    .B1(_10106_),
    .X(_10227_));
 sky130_fd_sc_hd__a21bo_1 _17208_ (.A1(_10101_),
    .A2(_10106_),
    .B1_N(_10105_),
    .X(_10228_));
 sky130_fd_sc_hd__nand3_1 _17209_ (.A(_10226_),
    .B(_10227_),
    .C(_10228_),
    .Y(_10229_));
 sky130_fd_sc_hd__a21o_1 _17210_ (.A1(_10226_),
    .A2(_10227_),
    .B1(_10228_),
    .X(_10230_));
 sky130_fd_sc_hd__and2_1 _17211_ (.A(_10229_),
    .B(_10230_),
    .X(_10231_));
 sky130_fd_sc_hd__xor2_1 _17212_ (.A(_10218_),
    .B(_10231_),
    .X(_10232_));
 sky130_fd_sc_hd__a21oi_2 _17213_ (.A1(_10094_),
    .A2(_10110_),
    .B1(_10108_),
    .Y(_10233_));
 sky130_fd_sc_hd__xnor2_1 _17214_ (.A(_10232_),
    .B(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__nand2_1 _17215_ (.A(_10207_),
    .B(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__or2_1 _17216_ (.A(_10207_),
    .B(_10234_),
    .X(_10236_));
 sky130_fd_sc_hd__nand2_2 _17217_ (.A(_10235_),
    .B(_10236_),
    .Y(_10237_));
 sky130_fd_sc_hd__nor2_1 _17218_ (.A(_10111_),
    .B(_10112_),
    .Y(_10238_));
 sky130_fd_sc_hd__a21oi_2 _17219_ (.A1(_10082_),
    .A2(_10113_),
    .B1(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__xor2_2 _17220_ (.A(_10237_),
    .B(_10239_),
    .X(_10240_));
 sky130_fd_sc_hd__xnor2_1 _17221_ (.A(_10182_),
    .B(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__a21oi_1 _17222_ (.A1(_10058_),
    .A2(_10118_),
    .B1(_10117_),
    .Y(_10242_));
 sky130_fd_sc_hd__nor2_1 _17223_ (.A(_10241_),
    .B(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__nand2_1 _17224_ (.A(_10241_),
    .B(_10242_),
    .Y(_10244_));
 sky130_fd_sc_hd__and2b_1 _17225_ (.A_N(_10243_),
    .B(_10244_),
    .X(_10245_));
 sky130_fd_sc_hd__xnor2_4 _17226_ (.A(_10146_),
    .B(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__nor2_1 _17227_ (.A(_10120_),
    .B(_10121_),
    .Y(_10247_));
 sky130_fd_sc_hd__a21oi_2 _17228_ (.A1(_10023_),
    .A2(_10122_),
    .B1(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__xor2_4 _17229_ (.A(_10246_),
    .B(_10248_),
    .X(_10249_));
 sky130_fd_sc_hd__xnor2_4 _17230_ (.A(_10021_),
    .B(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__nor2_1 _17231_ (.A(_10123_),
    .B(_10125_),
    .Y(_10251_));
 sky130_fd_sc_hd__a21oi_2 _17232_ (.A1(_09891_),
    .A2(_10126_),
    .B1(_10251_),
    .Y(_10252_));
 sky130_fd_sc_hd__xor2_4 _17233_ (.A(_10250_),
    .B(_10252_),
    .X(_10253_));
 sky130_fd_sc_hd__a21o_1 _17234_ (.A1(_10017_),
    .A2(_10018_),
    .B1(_10127_),
    .X(_10254_));
 sky130_fd_sc_hd__a21o_1 _17235_ (.A1(_10004_),
    .A2(_10254_),
    .B1(_10129_),
    .X(_10255_));
 sky130_fd_sc_hd__o31a_4 _17236_ (.A1(_10006_),
    .A2(_10008_),
    .A3(_10130_),
    .B1(_10255_),
    .X(_10256_));
 sky130_fd_sc_hd__xnor2_4 _17237_ (.A(_10253_),
    .B(_10256_),
    .Y(_10257_));
 sky130_fd_sc_hd__and2_1 _17238_ (.A(_08103_),
    .B(_10257_),
    .X(_10258_));
 sky130_fd_sc_hd__a31o_1 _17239_ (.A1(_09788_),
    .A2(_10139_),
    .A3(_10140_),
    .B1(_10258_),
    .X(_10259_));
 sky130_fd_sc_hd__clkbuf_8 _17240_ (.A(net4648),
    .X(_10260_));
 sky130_fd_sc_hd__mux2_1 _17241_ (.A0(_10259_),
    .A1(net4657),
    .S(_10260_),
    .X(_10261_));
 sky130_fd_sc_hd__clkbuf_1 _17242_ (.A(_10261_),
    .X(_00541_));
 sky130_fd_sc_hd__and2_1 _17243_ (.A(net4610),
    .B(net4405),
    .X(_10262_));
 sky130_fd_sc_hd__nor2_1 _17244_ (.A(net4610),
    .B(net4405),
    .Y(_10263_));
 sky130_fd_sc_hd__a211oi_1 _17245_ (.A1(_10136_),
    .A2(_10140_),
    .B1(_10262_),
    .C1(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__o211a_1 _17246_ (.A1(_10262_),
    .A2(_10263_),
    .B1(_10136_),
    .C1(_10140_),
    .X(_10265_));
 sky130_fd_sc_hd__or2_1 _17247_ (.A(_10250_),
    .B(_10252_),
    .X(_10266_));
 sky130_fd_sc_hd__inv_2 _17248_ (.A(_10253_),
    .Y(_10267_));
 sky130_fd_sc_hd__or2_1 _17249_ (.A(_10267_),
    .B(_10256_),
    .X(_10268_));
 sky130_fd_sc_hd__or2_1 _17250_ (.A(_10246_),
    .B(_10248_),
    .X(_10269_));
 sky130_fd_sc_hd__nand2_1 _17251_ (.A(_10021_),
    .B(_10249_),
    .Y(_10270_));
 sky130_fd_sc_hd__or2b_1 _17252_ (.A(_10181_),
    .B_N(_10147_),
    .X(_10271_));
 sky130_fd_sc_hd__a21oi_1 _17253_ (.A1(_10159_),
    .A2(_10160_),
    .B1(_10157_),
    .Y(_10272_));
 sky130_fd_sc_hd__a21oi_2 _17254_ (.A1(_10179_),
    .A2(_10271_),
    .B1(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__and3_1 _17255_ (.A(_10179_),
    .B(_10271_),
    .C(_10272_),
    .X(_10274_));
 sky130_fd_sc_hd__nor2_1 _17256_ (.A(_10273_),
    .B(_10274_),
    .Y(_10275_));
 sky130_fd_sc_hd__a21o_1 _17257_ (.A1(_10161_),
    .A2(_10177_),
    .B1(_10175_),
    .X(_10276_));
 sky130_fd_sc_hd__or2b_1 _17258_ (.A(_10206_),
    .B_N(_10183_),
    .X(_10277_));
 sky130_fd_sc_hd__and2_1 _17259_ (.A(_09373_),
    .B(net4909),
    .X(_10278_));
 sky130_fd_sc_hd__xnor2_1 _17260_ (.A(_10150_),
    .B(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__nor2_1 _17261_ (.A(_08226_),
    .B(_09472_),
    .Y(_10280_));
 sky130_fd_sc_hd__and2_1 _17262_ (.A(_10279_),
    .B(_10280_),
    .X(_10281_));
 sky130_fd_sc_hd__nor2_1 _17263_ (.A(_10279_),
    .B(_10280_),
    .Y(_10282_));
 sky130_fd_sc_hd__or2_1 _17264_ (.A(_10281_),
    .B(_10282_),
    .X(_10283_));
 sky130_fd_sc_hd__a21boi_1 _17265_ (.A1(_10153_),
    .A2(_10154_),
    .B1_N(_10152_),
    .Y(_10284_));
 sky130_fd_sc_hd__nor2_1 _17266_ (.A(_10283_),
    .B(_10284_),
    .Y(_10285_));
 sky130_fd_sc_hd__and2_1 _17267_ (.A(_10283_),
    .B(_10284_),
    .X(_10286_));
 sky130_fd_sc_hd__nor2_1 _17268_ (.A(_10285_),
    .B(_10286_),
    .Y(_10287_));
 sky130_fd_sc_hd__or3_1 _17269_ (.A(net8035),
    .B(_06124_),
    .C(_09413_),
    .X(_10288_));
 sky130_fd_sc_hd__buf_2 _17270_ (.A(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__nor2_1 _17271_ (.A(_09133_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__xor2_1 _17272_ (.A(_10287_),
    .B(_10290_),
    .X(_10291_));
 sky130_fd_sc_hd__a21bo_1 _17273_ (.A1(_10167_),
    .A2(_10168_),
    .B1_N(_10166_),
    .X(_10292_));
 sky130_fd_sc_hd__o22a_1 _17274_ (.A1(_10190_),
    .A2(_08614_),
    .B1(_09062_),
    .B2(_08383_),
    .X(_10293_));
 sky130_fd_sc_hd__or4_1 _17275_ (.A(_10190_),
    .B(_08383_),
    .C(_08614_),
    .D(_09062_),
    .X(_10294_));
 sky130_fd_sc_hd__and2b_1 _17276_ (.A_N(_10293_),
    .B(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__nor2_1 _17277_ (.A(_08661_),
    .B(_09116_),
    .Y(_10296_));
 sky130_fd_sc_hd__xnor2_1 _17278_ (.A(_10295_),
    .B(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__a21bo_1 _17279_ (.A1(_10189_),
    .A2(_10191_),
    .B1_N(_10188_),
    .X(_10298_));
 sky130_fd_sc_hd__and2b_1 _17280_ (.A_N(_10297_),
    .B(_10298_),
    .X(_10299_));
 sky130_fd_sc_hd__and2b_1 _17281_ (.A_N(_10298_),
    .B(_10297_),
    .X(_10300_));
 sky130_fd_sc_hd__nor2_1 _17282_ (.A(_10299_),
    .B(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__xnor2_1 _17283_ (.A(_10292_),
    .B(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__a21oi_1 _17284_ (.A1(_10162_),
    .A2(_10172_),
    .B1(_10170_),
    .Y(_10303_));
 sky130_fd_sc_hd__nor2_1 _17285_ (.A(_10302_),
    .B(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__and2_1 _17286_ (.A(_10302_),
    .B(_10303_),
    .X(_10305_));
 sky130_fd_sc_hd__nor2_1 _17287_ (.A(_10304_),
    .B(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__xnor2_1 _17288_ (.A(_10291_),
    .B(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__a21o_1 _17289_ (.A1(_10204_),
    .A2(_10277_),
    .B1(_10307_),
    .X(_10308_));
 sky130_fd_sc_hd__nand3_1 _17290_ (.A(_10204_),
    .B(_10277_),
    .C(_10307_),
    .Y(_10309_));
 sky130_fd_sc_hd__nand2_1 _17291_ (.A(_10308_),
    .B(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__xnor2_2 _17292_ (.A(_10276_),
    .B(_10310_),
    .Y(_10311_));
 sky130_fd_sc_hd__or2b_1 _17293_ (.A(_10192_),
    .B_N(_10202_),
    .X(_10312_));
 sky130_fd_sc_hd__o21ai_1 _17294_ (.A1(_10199_),
    .A2(_10201_),
    .B1(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand2_1 _17295_ (.A(_10210_),
    .B(_10216_),
    .Y(_10314_));
 sky130_fd_sc_hd__or2b_1 _17296_ (.A(_10217_),
    .B_N(_10208_),
    .X(_10315_));
 sky130_fd_sc_hd__a21oi_4 _17297_ (.A1(_08421_),
    .A2(_08424_),
    .B1(_08426_),
    .Y(_10316_));
 sky130_fd_sc_hd__nor2_1 _17298_ (.A(_08338_),
    .B(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__xnor2_1 _17299_ (.A(_10187_),
    .B(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__or3_1 _17300_ (.A(_10163_),
    .B(net8008),
    .C(_10318_),
    .X(_10319_));
 sky130_fd_sc_hd__o21ai_1 _17301_ (.A1(_10163_),
    .A2(net8008),
    .B1(_10318_),
    .Y(_10320_));
 sky130_fd_sc_hd__and2_1 _17302_ (.A(_10319_),
    .B(_10320_),
    .X(_10321_));
 sky130_fd_sc_hd__or2_1 _17303_ (.A(_08309_),
    .B(_09170_),
    .X(_10322_));
 sky130_fd_sc_hd__nor2_1 _17304_ (.A(_08326_),
    .B(_09403_),
    .Y(_10323_));
 sky130_fd_sc_hd__xor2_2 _17305_ (.A(_10322_),
    .B(_10323_),
    .X(_10324_));
 sky130_fd_sc_hd__or2_1 _17306_ (.A(_09262_),
    .B(_09165_),
    .X(_10325_));
 sky130_fd_sc_hd__xnor2_2 _17307_ (.A(_10324_),
    .B(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__clkbuf_4 _17308_ (.A(_08326_),
    .X(_10327_));
 sky130_fd_sc_hd__o31a_1 _17309_ (.A1(_10327_),
    .A2(_09170_),
    .A3(_10193_),
    .B1(_10197_),
    .X(_10328_));
 sky130_fd_sc_hd__xor2_1 _17310_ (.A(_10326_),
    .B(_10328_),
    .X(_10329_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(_10321_),
    .B(_10329_),
    .Y(_10330_));
 sky130_fd_sc_hd__or2_1 _17312_ (.A(_10321_),
    .B(_10329_),
    .X(_10331_));
 sky130_fd_sc_hd__nand2_1 _17313_ (.A(_10330_),
    .B(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__a21o_1 _17314_ (.A1(_10314_),
    .A2(_10315_),
    .B1(_10332_),
    .X(_10333_));
 sky130_fd_sc_hd__nand3_1 _17315_ (.A(_10314_),
    .B(_10315_),
    .C(_10332_),
    .Y(_10334_));
 sky130_fd_sc_hd__nand2_1 _17316_ (.A(_10333_),
    .B(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__xnor2_1 _17317_ (.A(_10313_),
    .B(_10335_),
    .Y(_10336_));
 sky130_fd_sc_hd__a21bo_1 _17318_ (.A1(_10213_),
    .A2(_10215_),
    .B1_N(_10212_),
    .X(_10337_));
 sky130_fd_sc_hd__nand2_1 _17319_ (.A(_10223_),
    .B(_10224_),
    .Y(_10338_));
 sky130_fd_sc_hd__or4_1 _17320_ (.A(_08918_),
    .B(_10211_),
    .C(_10096_),
    .D(_10220_),
    .X(_10339_));
 sky130_fd_sc_hd__o22ai_1 _17321_ (.A1(_10211_),
    .A2(_10096_),
    .B1(_10220_),
    .B2(_08918_),
    .Y(_10340_));
 sky130_fd_sc_hd__nand2_1 _17322_ (.A(_10339_),
    .B(_10340_),
    .Y(_10341_));
 sky130_fd_sc_hd__nor2_1 _17323_ (.A(_09272_),
    .B(_09664_),
    .Y(_10342_));
 sky130_fd_sc_hd__xor2_1 _17324_ (.A(_10341_),
    .B(_10342_),
    .X(_10343_));
 sky130_fd_sc_hd__xor2_1 _17325_ (.A(_10338_),
    .B(_10343_),
    .X(_10344_));
 sky130_fd_sc_hd__xnor2_1 _17326_ (.A(_10337_),
    .B(_10344_),
    .Y(_10345_));
 sky130_fd_sc_hd__buf_2 _17327_ (.A(_09976_),
    .X(_10346_));
 sky130_fd_sc_hd__nor2_1 _17328_ (.A(_09537_),
    .B(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__or3_2 _17329_ (.A(_08948_),
    .B(_08916_),
    .C(_09970_),
    .X(_10348_));
 sky130_fd_sc_hd__a21oi_1 _17330_ (.A1(_08948_),
    .A2(_08916_),
    .B1(_09970_),
    .Y(_10349_));
 sky130_fd_sc_hd__nand2_2 _17331_ (.A(_10348_),
    .B(_10349_),
    .Y(_10350_));
 sky130_fd_sc_hd__xnor2_2 _17332_ (.A(_10347_),
    .B(_10350_),
    .Y(_10351_));
 sky130_fd_sc_hd__xnor2_1 _17333_ (.A(_10106_),
    .B(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__and2_1 _17334_ (.A(_10105_),
    .B(_10226_),
    .X(_10353_));
 sky130_fd_sc_hd__xor2_1 _17335_ (.A(_10352_),
    .B(_10353_),
    .X(_10354_));
 sky130_fd_sc_hd__xnor2_1 _17336_ (.A(_10345_),
    .B(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__a21boi_1 _17337_ (.A1(_10218_),
    .A2(_10230_),
    .B1_N(_10229_),
    .Y(_10356_));
 sky130_fd_sc_hd__nor2_1 _17338_ (.A(_10355_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__and2_1 _17339_ (.A(_10355_),
    .B(_10356_),
    .X(_10358_));
 sky130_fd_sc_hd__nor2_1 _17340_ (.A(_10357_),
    .B(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__xnor2_1 _17341_ (.A(_10336_),
    .B(_10359_),
    .Y(_10360_));
 sky130_fd_sc_hd__and2_1 _17342_ (.A(_10218_),
    .B(_10231_),
    .X(_10361_));
 sky130_fd_sc_hd__nor2_1 _17343_ (.A(_10218_),
    .B(_10231_),
    .Y(_10362_));
 sky130_fd_sc_hd__o31a_1 _17344_ (.A1(_10361_),
    .A2(_10362_),
    .A3(_10233_),
    .B1(_10235_),
    .X(_10363_));
 sky130_fd_sc_hd__nor2_1 _17345_ (.A(_10360_),
    .B(_10363_),
    .Y(_10364_));
 sky130_fd_sc_hd__and2_1 _17346_ (.A(_10360_),
    .B(_10363_),
    .X(_10365_));
 sky130_fd_sc_hd__nor2_1 _17347_ (.A(_10364_),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__xnor2_2 _17348_ (.A(_10311_),
    .B(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__nor2_1 _17349_ (.A(_10237_),
    .B(_10239_),
    .Y(_10368_));
 sky130_fd_sc_hd__a21oi_2 _17350_ (.A1(_10182_),
    .A2(_10240_),
    .B1(_10368_),
    .Y(_10369_));
 sky130_fd_sc_hd__xor2_2 _17351_ (.A(_10367_),
    .B(_10369_),
    .X(_10370_));
 sky130_fd_sc_hd__xnor2_2 _17352_ (.A(_10275_),
    .B(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__a21oi_2 _17353_ (.A1(_10146_),
    .A2(_10244_),
    .B1(_10243_),
    .Y(_10372_));
 sky130_fd_sc_hd__xor2_2 _17354_ (.A(_10371_),
    .B(_10372_),
    .X(_10373_));
 sky130_fd_sc_hd__xnor2_2 _17355_ (.A(_10144_),
    .B(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__a21oi_1 _17356_ (.A1(_10269_),
    .A2(_10270_),
    .B1(_10374_),
    .Y(_10375_));
 sky130_fd_sc_hd__and3_1 _17357_ (.A(_10269_),
    .B(_10270_),
    .C(_10374_),
    .X(_10376_));
 sky130_fd_sc_hd__or2_1 _17358_ (.A(_10375_),
    .B(_10376_),
    .X(_10377_));
 sky130_fd_sc_hd__a21o_1 _17359_ (.A1(_10266_),
    .A2(_10268_),
    .B1(_10377_),
    .X(_10378_));
 sky130_fd_sc_hd__nand2_1 _17360_ (.A(_08103_),
    .B(_10378_),
    .Y(_10379_));
 sky130_fd_sc_hd__a31o_2 _17361_ (.A1(_10266_),
    .A2(_10268_),
    .A3(_10377_),
    .B1(_10379_),
    .X(_10380_));
 sky130_fd_sc_hd__o31ai_1 _17362_ (.A1(_09809_),
    .A2(_10264_),
    .A3(_10265_),
    .B1(_10380_),
    .Y(_10381_));
 sky130_fd_sc_hd__mux2_1 _17363_ (.A0(_10381_),
    .A1(net4610),
    .S(_10260_),
    .X(_10382_));
 sky130_fd_sc_hd__clkbuf_1 _17364_ (.A(_10382_),
    .X(_00542_));
 sky130_fd_sc_hd__nand2_1 _17365_ (.A(net4651),
    .B(net4522),
    .Y(_10383_));
 sky130_fd_sc_hd__or2_1 _17366_ (.A(net4651),
    .B(net4522),
    .X(_10384_));
 sky130_fd_sc_hd__nand2_1 _17367_ (.A(_10383_),
    .B(_10384_),
    .Y(_10385_));
 sky130_fd_sc_hd__nor2_1 _17368_ (.A(_10262_),
    .B(_10264_),
    .Y(_10386_));
 sky130_fd_sc_hd__xnor2_1 _17369_ (.A(_10385_),
    .B(_10386_),
    .Y(_10387_));
 sky130_fd_sc_hd__or2b_1 _17370_ (.A(_10310_),
    .B_N(_10276_),
    .X(_10388_));
 sky130_fd_sc_hd__a21oi_1 _17371_ (.A1(_10287_),
    .A2(_10290_),
    .B1(_10285_),
    .Y(_10389_));
 sky130_fd_sc_hd__a21oi_2 _17372_ (.A1(_10308_),
    .A2(_10388_),
    .B1(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__and3_1 _17373_ (.A(_10308_),
    .B(_10388_),
    .C(_10389_),
    .X(_10391_));
 sky130_fd_sc_hd__nor2_1 _17374_ (.A(_10390_),
    .B(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__a21o_1 _17375_ (.A1(_10291_),
    .A2(_10306_),
    .B1(_10304_),
    .X(_10393_));
 sky130_fd_sc_hd__or2b_1 _17376_ (.A(_10335_),
    .B_N(_10313_),
    .X(_10394_));
 sky130_fd_sc_hd__nand2_1 _17377_ (.A(_08167_),
    .B(net4909),
    .Y(_10395_));
 sky130_fd_sc_hd__nand2_1 _17378_ (.A(_09373_),
    .B(net4914),
    .Y(_10396_));
 sky130_fd_sc_hd__and3_1 _17379_ (.A(_08167_),
    .B(net4914),
    .C(_10278_),
    .X(_10397_));
 sky130_fd_sc_hd__a21oi_1 _17380_ (.A1(_10395_),
    .A2(_10396_),
    .B1(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__and2b_1 _17381_ (.A_N(_09612_),
    .B(_09249_),
    .X(_10399_));
 sky130_fd_sc_hd__xnor2_1 _17382_ (.A(_10398_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__a21oi_1 _17383_ (.A1(_10151_),
    .A2(_10278_),
    .B1(_10281_),
    .Y(_10401_));
 sky130_fd_sc_hd__nor2_1 _17384_ (.A(_10400_),
    .B(_10401_),
    .Y(_10402_));
 sky130_fd_sc_hd__and2_1 _17385_ (.A(_10400_),
    .B(_10401_),
    .X(_10403_));
 sky130_fd_sc_hd__nor2_1 _17386_ (.A(_10402_),
    .B(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__nor2_1 _17387_ (.A(_08864_),
    .B(_10289_),
    .Y(_10405_));
 sky130_fd_sc_hd__xor2_1 _17388_ (.A(_10404_),
    .B(_10405_),
    .X(_10406_));
 sky130_fd_sc_hd__a21bo_1 _17389_ (.A1(_10295_),
    .A2(_10296_),
    .B1_N(_10294_),
    .X(_10407_));
 sky130_fd_sc_hd__o21a_2 _17390_ (.A1(_08115_),
    .A2(_08369_),
    .B1(_08371_),
    .X(_10408_));
 sky130_fd_sc_hd__nor2_1 _17391_ (.A(_10408_),
    .B(_09062_),
    .Y(_10409_));
 sky130_fd_sc_hd__nor2_1 _17392_ (.A(_08413_),
    .B(_08612_),
    .Y(_10410_));
 sky130_fd_sc_hd__xnor2_1 _17393_ (.A(_10409_),
    .B(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__or3_1 _17394_ (.A(_09915_),
    .B(_09116_),
    .C(_10411_),
    .X(_10412_));
 sky130_fd_sc_hd__o21ai_1 _17395_ (.A1(_09915_),
    .A2(_09116_),
    .B1(_10411_),
    .Y(_10413_));
 sky130_fd_sc_hd__nand2_1 _17396_ (.A(_10412_),
    .B(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__a21bo_1 _17397_ (.A1(_10187_),
    .A2(_10317_),
    .B1_N(_10319_),
    .X(_10415_));
 sky130_fd_sc_hd__and2b_1 _17398_ (.A_N(_10414_),
    .B(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__and2b_1 _17399_ (.A_N(_10415_),
    .B(_10414_),
    .X(_10417_));
 sky130_fd_sc_hd__nor2_1 _17400_ (.A(_10416_),
    .B(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__xnor2_1 _17401_ (.A(_10407_),
    .B(_10418_),
    .Y(_10419_));
 sky130_fd_sc_hd__a21oi_1 _17402_ (.A1(_10292_),
    .A2(_10301_),
    .B1(_10299_),
    .Y(_10420_));
 sky130_fd_sc_hd__nor2_1 _17403_ (.A(_10419_),
    .B(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__and2_1 _17404_ (.A(_10419_),
    .B(_10420_),
    .X(_10422_));
 sky130_fd_sc_hd__nor2_1 _17405_ (.A(_10421_),
    .B(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__xnor2_1 _17406_ (.A(_10406_),
    .B(_10423_),
    .Y(_10424_));
 sky130_fd_sc_hd__a21o_1 _17407_ (.A1(_10333_),
    .A2(_10394_),
    .B1(_10424_),
    .X(_10425_));
 sky130_fd_sc_hd__nand3_1 _17408_ (.A(_10333_),
    .B(_10394_),
    .C(_10424_),
    .Y(_10426_));
 sky130_fd_sc_hd__nand2_1 _17409_ (.A(_10425_),
    .B(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__xnor2_1 _17410_ (.A(_10393_),
    .B(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__o21ai_2 _17411_ (.A1(_10326_),
    .A2(_10328_),
    .B1(_10330_),
    .Y(_10429_));
 sky130_fd_sc_hd__or2b_1 _17412_ (.A(_10343_),
    .B_N(_10338_),
    .X(_10430_));
 sky130_fd_sc_hd__or2b_1 _17413_ (.A(_10344_),
    .B_N(_10337_),
    .X(_10431_));
 sky130_fd_sc_hd__nand2_1 _17414_ (.A(_08427_),
    .B(_08428_),
    .Y(_10432_));
 sky130_fd_sc_hd__or2_1 _17415_ (.A(_08140_),
    .B(_10432_),
    .X(_10433_));
 sky130_fd_sc_hd__nor2_1 _17416_ (.A(_10062_),
    .B(_08461_),
    .Y(_10434_));
 sky130_fd_sc_hd__xnor2_1 _17417_ (.A(_10433_),
    .B(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__nor2_1 _17418_ (.A(_08472_),
    .B(_08616_),
    .Y(_10436_));
 sky130_fd_sc_hd__nand2_1 _17419_ (.A(_10435_),
    .B(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__or2_1 _17420_ (.A(_10435_),
    .B(_10436_),
    .X(_10438_));
 sky130_fd_sc_hd__and2_1 _17421_ (.A(_10437_),
    .B(_10438_),
    .X(_01663_));
 sky130_fd_sc_hd__or2_1 _17422_ (.A(_08799_),
    .B(_09403_),
    .X(_01664_));
 sky130_fd_sc_hd__nor2_1 _17423_ (.A(_08326_),
    .B(_09664_),
    .Y(_01665_));
 sky130_fd_sc_hd__xnor2_1 _17424_ (.A(_01664_),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__nor2_1 _17425_ (.A(_09262_),
    .B(_09170_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _17426_ (.A(_01666_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__or2_1 _17427_ (.A(_01666_),
    .B(_01667_),
    .X(_01669_));
 sky130_fd_sc_hd__nand2_1 _17428_ (.A(_01668_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__or2_1 _17429_ (.A(_10324_),
    .B(_10325_),
    .X(_01671_));
 sky130_fd_sc_hd__o31a_1 _17430_ (.A1(_10327_),
    .A2(_09403_),
    .A3(_10322_),
    .B1(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__xor2_1 _17431_ (.A(_01670_),
    .B(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__nand2_1 _17432_ (.A(_01663_),
    .B(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__or2_1 _17433_ (.A(_01663_),
    .B(_01673_),
    .X(_01675_));
 sky130_fd_sc_hd__nand2_1 _17434_ (.A(_01674_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21o_1 _17435_ (.A1(_10430_),
    .A2(_10431_),
    .B1(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__nand3_1 _17436_ (.A(_10430_),
    .B(_10431_),
    .C(_01676_),
    .Y(_01678_));
 sky130_fd_sc_hd__nand2_1 _17437_ (.A(_01677_),
    .B(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__xnor2_1 _17438_ (.A(_10429_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__a21bo_1 _17439_ (.A1(_10340_),
    .A2(_10342_),
    .B1_N(_10339_),
    .X(_01681_));
 sky130_fd_sc_hd__or3_1 _17440_ (.A(_09537_),
    .B(_10346_),
    .C(_10350_),
    .X(_01682_));
 sky130_fd_sc_hd__or4_1 _17441_ (.A(_08918_),
    .B(_10211_),
    .C(_10220_),
    .D(_10346_),
    .X(_01683_));
 sky130_fd_sc_hd__o22ai_1 _17442_ (.A1(_10211_),
    .A2(_10220_),
    .B1(_10346_),
    .B2(_08918_),
    .Y(_01684_));
 sky130_fd_sc_hd__nand2_1 _17443_ (.A(_01683_),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__nor2_1 _17444_ (.A(_09272_),
    .B(_10096_),
    .Y(_01686_));
 sky130_fd_sc_hd__xor2_1 _17445_ (.A(_01685_),
    .B(_01686_),
    .X(_01687_));
 sky130_fd_sc_hd__a21o_1 _17446_ (.A1(_10348_),
    .A2(_01682_),
    .B1(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__nand3_1 _17447_ (.A(_10348_),
    .B(_01682_),
    .C(_01687_),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _17448_ (.A(_01688_),
    .B(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__xnor2_1 _17449_ (.A(_01681_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _17450_ (.A(_10106_),
    .B(_10351_),
    .Y(_01692_));
 sky130_fd_sc_hd__buf_2 _17451_ (.A(_09970_),
    .X(_01693_));
 sky130_fd_sc_hd__nor2_1 _17452_ (.A(_09537_),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__mux2_1 _17453_ (.A0(_09537_),
    .A1(_01694_),
    .S(_10350_),
    .X(_01695_));
 sky130_fd_sc_hd__xnor2_1 _17454_ (.A(_10106_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__a21oi_1 _17455_ (.A1(_10105_),
    .A2(_01692_),
    .B1(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__and3_1 _17456_ (.A(_10105_),
    .B(_01692_),
    .C(_01696_),
    .X(_01698_));
 sky130_fd_sc_hd__nor2_1 _17457_ (.A(_01697_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__xnor2_1 _17458_ (.A(_01691_),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__nor2_1 _17459_ (.A(_10352_),
    .B(_10353_),
    .Y(_01701_));
 sky130_fd_sc_hd__a21oi_1 _17460_ (.A1(_10345_),
    .A2(_10354_),
    .B1(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nor2_1 _17461_ (.A(_01700_),
    .B(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__and2_1 _17462_ (.A(_01700_),
    .B(_01702_),
    .X(_01704_));
 sky130_fd_sc_hd__nor2_1 _17463_ (.A(_01703_),
    .B(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__xnor2_1 _17464_ (.A(_01680_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__a21oi_1 _17465_ (.A1(_10336_),
    .A2(_10359_),
    .B1(_10357_),
    .Y(_01707_));
 sky130_fd_sc_hd__xor2_1 _17466_ (.A(_01706_),
    .B(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__xnor2_1 _17467_ (.A(_10428_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__a21oi_1 _17468_ (.A1(_10311_),
    .A2(_10366_),
    .B1(_10364_),
    .Y(_01710_));
 sky130_fd_sc_hd__nor2_1 _17469_ (.A(_01709_),
    .B(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hd__and2_1 _17470_ (.A(_01709_),
    .B(_01710_),
    .X(_01712_));
 sky130_fd_sc_hd__nor2_1 _17471_ (.A(_01711_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__xnor2_1 _17472_ (.A(_10392_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__nor2_1 _17473_ (.A(_10367_),
    .B(_10369_),
    .Y(_01715_));
 sky130_fd_sc_hd__a21oi_1 _17474_ (.A1(_10275_),
    .A2(_10370_),
    .B1(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__xor2_1 _17475_ (.A(_01714_),
    .B(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__xnor2_1 _17476_ (.A(_10273_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__nor2_1 _17477_ (.A(_10371_),
    .B(_10372_),
    .Y(_01719_));
 sky130_fd_sc_hd__a21oi_1 _17478_ (.A1(_10144_),
    .A2(_10373_),
    .B1(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor2_1 _17479_ (.A(_01718_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__and2_1 _17480_ (.A(_01718_),
    .B(_01720_),
    .X(_01722_));
 sky130_fd_sc_hd__or2_1 _17481_ (.A(_01721_),
    .B(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__a21o_1 _17482_ (.A1(_10269_),
    .A2(_10270_),
    .B1(_10374_),
    .X(_01724_));
 sky130_fd_sc_hd__a21o_1 _17483_ (.A1(_10266_),
    .A2(_01724_),
    .B1(_10376_),
    .X(_01725_));
 sky130_fd_sc_hd__o31a_4 _17484_ (.A1(_10267_),
    .A2(_10256_),
    .A3(_10377_),
    .B1(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__and2_1 _17485_ (.A(_01723_),
    .B(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__nor2_1 _17486_ (.A(_01723_),
    .B(_01726_),
    .Y(_01728_));
 sky130_fd_sc_hd__or3_4 _17487_ (.A(net90),
    .B(_01727_),
    .C(_01728_),
    .X(_01729_));
 sky130_fd_sc_hd__o21ai_1 _17488_ (.A1(_06058_),
    .A2(_10387_),
    .B1(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__mux2_1 _17489_ (.A0(_01730_),
    .A1(net4651),
    .S(_10260_),
    .X(_01731_));
 sky130_fd_sc_hd__clkbuf_1 _17490_ (.A(_01731_),
    .X(_00543_));
 sky130_fd_sc_hd__nor2_1 _17491_ (.A(net4659),
    .B(net4653),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_1 _17492_ (.A(net4659),
    .B(net4653),
    .Y(_01733_));
 sky130_fd_sc_hd__or2b_1 _17493_ (.A(_01732_),
    .B_N(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__o21a_1 _17494_ (.A1(_10385_),
    .A2(_10386_),
    .B1(_10383_),
    .X(_01735_));
 sky130_fd_sc_hd__xnor2_1 _17495_ (.A(_01734_),
    .B(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__or2_1 _17496_ (.A(_01714_),
    .B(_01716_),
    .X(_01737_));
 sky130_fd_sc_hd__nand2_1 _17497_ (.A(_10273_),
    .B(_01717_),
    .Y(_01738_));
 sky130_fd_sc_hd__or2b_1 _17498_ (.A(_10427_),
    .B_N(_10393_),
    .X(_01739_));
 sky130_fd_sc_hd__a21oi_1 _17499_ (.A1(_10404_),
    .A2(_10405_),
    .B1(_10402_),
    .Y(_01740_));
 sky130_fd_sc_hd__a21oi_2 _17500_ (.A1(_10425_),
    .A2(_01739_),
    .B1(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__and3_1 _17501_ (.A(_10425_),
    .B(_01739_),
    .C(_01740_),
    .X(_01742_));
 sky130_fd_sc_hd__nor2_1 _17502_ (.A(_01741_),
    .B(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__a21o_1 _17503_ (.A1(_10406_),
    .A2(_10423_),
    .B1(_10421_),
    .X(_01744_));
 sky130_fd_sc_hd__or2b_1 _17504_ (.A(_01679_),
    .B_N(_10429_),
    .X(_01745_));
 sky130_fd_sc_hd__nand2_1 _17505_ (.A(_08167_),
    .B(net4914),
    .Y(_01746_));
 sky130_fd_sc_hd__or2_1 _17506_ (.A(_09915_),
    .B(_09225_),
    .X(_01747_));
 sky130_fd_sc_hd__or2_1 _17507_ (.A(_09915_),
    .B(_09345_),
    .X(_01748_));
 sky130_fd_sc_hd__nor2_1 _17508_ (.A(_10395_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__a21oi_1 _17509_ (.A1(_01746_),
    .A2(_01747_),
    .B1(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__and2b_1 _17510_ (.A_N(_09612_),
    .B(_09373_),
    .X(_01751_));
 sky130_fd_sc_hd__xnor2_1 _17511_ (.A(_01750_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__a21oi_1 _17512_ (.A1(_10398_),
    .A2(_10399_),
    .B1(_10397_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_1 _17513_ (.A(_01752_),
    .B(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__and2_1 _17514_ (.A(_01752_),
    .B(_01753_),
    .X(_01755_));
 sky130_fd_sc_hd__nor2_1 _17515_ (.A(_01754_),
    .B(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__nor2_1 _17516_ (.A(_09249_),
    .B(_10289_),
    .Y(_01757_));
 sky130_fd_sc_hd__xor2_1 _17517_ (.A(_01756_),
    .B(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__a21bo_1 _17518_ (.A1(_10409_),
    .A2(_10410_),
    .B1_N(_10412_),
    .X(_01759_));
 sky130_fd_sc_hd__buf_2 _17519_ (.A(_08461_),
    .X(_01760_));
 sky130_fd_sc_hd__or3_1 _17520_ (.A(_10062_),
    .B(_01760_),
    .C(_10433_),
    .X(_01761_));
 sky130_fd_sc_hd__or2_1 _17521_ (.A(_08472_),
    .B(_08614_),
    .X(_01762_));
 sky130_fd_sc_hd__or3_1 _17522_ (.A(_10163_),
    .B(_09060_),
    .C(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__o21ai_1 _17523_ (.A1(_10163_),
    .A2(_09060_),
    .B1(_01762_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(_01763_),
    .B(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_1 _17525_ (.A(_10190_),
    .B(_09116_),
    .Y(_01766_));
 sky130_fd_sc_hd__xor2_1 _17526_ (.A(_01765_),
    .B(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__a21oi_1 _17527_ (.A1(_01761_),
    .A2(_10437_),
    .B1(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__and3_1 _17528_ (.A(_01761_),
    .B(_10437_),
    .C(_01767_),
    .X(_01769_));
 sky130_fd_sc_hd__nor2_1 _17529_ (.A(_01768_),
    .B(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__xnor2_1 _17530_ (.A(_01759_),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__a21oi_1 _17531_ (.A1(_10407_),
    .A2(_10418_),
    .B1(_10416_),
    .Y(_01772_));
 sky130_fd_sc_hd__nor2_1 _17532_ (.A(_01771_),
    .B(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__and2_1 _17533_ (.A(_01771_),
    .B(_01772_),
    .X(_01774_));
 sky130_fd_sc_hd__nor2_1 _17534_ (.A(_01773_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__xnor2_1 _17535_ (.A(_01758_),
    .B(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__a21o_1 _17536_ (.A1(_01677_),
    .A2(_01745_),
    .B1(_01776_),
    .X(_01777_));
 sky130_fd_sc_hd__nand3_1 _17537_ (.A(_01677_),
    .B(_01745_),
    .C(_01776_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand2_1 _17538_ (.A(_01777_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__xnor2_1 _17539_ (.A(_01744_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__o21ai_1 _17540_ (.A1(_01670_),
    .A2(_01672_),
    .B1(_01674_),
    .Y(_01781_));
 sky130_fd_sc_hd__or2b_1 _17541_ (.A(_01690_),
    .B_N(_01681_),
    .X(_01782_));
 sky130_fd_sc_hd__or2_1 _17542_ (.A(_10062_),
    .B(_09040_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_2 _17543_ (.A(_08140_),
    .X(_01784_));
 sky130_fd_sc_hd__nor2_1 _17544_ (.A(_01784_),
    .B(_01760_),
    .Y(_01785_));
 sky130_fd_sc_hd__xnor2_1 _17545_ (.A(_01783_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__nor2_1 _17546_ (.A(_10316_),
    .B(_08616_),
    .Y(_01787_));
 sky130_fd_sc_hd__nand2_1 _17547_ (.A(_01786_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__or2_1 _17548_ (.A(_01786_),
    .B(_01787_),
    .X(_01789_));
 sky130_fd_sc_hd__and2_1 _17549_ (.A(_01788_),
    .B(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__nor2_1 _17550_ (.A(_08799_),
    .B(_09664_),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _17551_ (.A(_10327_),
    .B(_10096_),
    .Y(_01792_));
 sky130_fd_sc_hd__xnor2_1 _17552_ (.A(_01791_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__buf_2 _17553_ (.A(_09262_),
    .X(_01794_));
 sky130_fd_sc_hd__nor2_1 _17554_ (.A(_01794_),
    .B(_09403_),
    .Y(_01795_));
 sky130_fd_sc_hd__xor2_1 _17555_ (.A(_01793_),
    .B(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__o31a_1 _17556_ (.A1(_10327_),
    .A2(_09664_),
    .A3(_01664_),
    .B1(_01668_),
    .X(_01797_));
 sky130_fd_sc_hd__nor2_1 _17557_ (.A(_01796_),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__and2_1 _17558_ (.A(_01796_),
    .B(_01797_),
    .X(_01799_));
 sky130_fd_sc_hd__nor2_1 _17559_ (.A(_01798_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__xnor2_1 _17560_ (.A(_01790_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__a21o_1 _17561_ (.A1(_01688_),
    .A2(_01782_),
    .B1(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__nand3_1 _17562_ (.A(_01688_),
    .B(_01782_),
    .C(_01801_),
    .Y(_01803_));
 sky130_fd_sc_hd__nand2_1 _17563_ (.A(_01802_),
    .B(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__xnor2_1 _17564_ (.A(_01781_),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__a21bo_1 _17565_ (.A1(_01684_),
    .A2(_01686_),
    .B1_N(_01683_),
    .X(_01806_));
 sky130_fd_sc_hd__o21ai_4 _17566_ (.A1(_09537_),
    .A2(_10350_),
    .B1(_10348_),
    .Y(_01807_));
 sky130_fd_sc_hd__o22ai_2 _17567_ (.A1(_08918_),
    .A2(_01693_),
    .B1(_10346_),
    .B2(_10211_),
    .Y(_01808_));
 sky130_fd_sc_hd__or4_1 _17568_ (.A(_08918_),
    .B(_10211_),
    .C(_01693_),
    .D(_10346_),
    .X(_01809_));
 sky130_fd_sc_hd__nand2_1 _17569_ (.A(_01808_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _17570_ (.A(_09272_),
    .B(_10220_),
    .Y(_01811_));
 sky130_fd_sc_hd__xnor2_1 _17571_ (.A(_01810_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__xnor2_1 _17572_ (.A(_01807_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__xnor2_1 _17573_ (.A(_01806_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nand2b_2 _17574_ (.A_N(_10105_),
    .B(_01695_),
    .Y(_01815_));
 sky130_fd_sc_hd__or3_1 _17575_ (.A(_10102_),
    .B(_10103_),
    .C(_01695_),
    .X(_01816_));
 sky130_fd_sc_hd__and2_1 _17576_ (.A(_01815_),
    .B(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__clkbuf_2 _17577_ (.A(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__nand2_1 _17578_ (.A(_01814_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__or2_1 _17579_ (.A(_01814_),
    .B(_01818_),
    .X(_01820_));
 sky130_fd_sc_hd__nand2_1 _17580_ (.A(_01819_),
    .B(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__a21oi_1 _17581_ (.A1(_01691_),
    .A2(_01699_),
    .B1(_01697_),
    .Y(_01822_));
 sky130_fd_sc_hd__nor2_1 _17582_ (.A(_01821_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__and2_1 _17583_ (.A(_01821_),
    .B(_01822_),
    .X(_01824_));
 sky130_fd_sc_hd__nor2_1 _17584_ (.A(_01823_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__xnor2_1 _17585_ (.A(_01805_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__a21oi_1 _17586_ (.A1(_01680_),
    .A2(_01705_),
    .B1(_01703_),
    .Y(_01827_));
 sky130_fd_sc_hd__nor2_1 _17587_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__and2_1 _17588_ (.A(_01826_),
    .B(_01827_),
    .X(_01829_));
 sky130_fd_sc_hd__nor2_1 _17589_ (.A(_01828_),
    .B(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__xnor2_1 _17590_ (.A(_01780_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__nor2_1 _17591_ (.A(_01706_),
    .B(_01707_),
    .Y(_01832_));
 sky130_fd_sc_hd__a21oi_1 _17592_ (.A1(_10428_),
    .A2(_01708_),
    .B1(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__xor2_1 _17593_ (.A(_01831_),
    .B(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__xnor2_1 _17594_ (.A(_01743_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__a21oi_1 _17595_ (.A1(_10392_),
    .A2(_01713_),
    .B1(_01711_),
    .Y(_01836_));
 sky130_fd_sc_hd__xor2_1 _17596_ (.A(_01835_),
    .B(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__xnor2_1 _17597_ (.A(_10390_),
    .B(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand3_1 _17598_ (.A(_01737_),
    .B(_01738_),
    .C(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__a21o_1 _17599_ (.A1(_01737_),
    .A2(_01738_),
    .B1(_01838_),
    .X(_01840_));
 sky130_fd_sc_hd__nand2_1 _17600_ (.A(_01839_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__nor2_1 _17601_ (.A(_01721_),
    .B(_01728_),
    .Y(_01842_));
 sky130_fd_sc_hd__o21ai_1 _17602_ (.A1(_01841_),
    .A2(_01842_),
    .B1(_06057_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21o_2 _17603_ (.A1(_01841_),
    .A2(_01842_),
    .B1(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__o21ai_1 _17604_ (.A1(_06058_),
    .A2(_01736_),
    .B1(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__mux2_1 _17605_ (.A0(_01845_),
    .A1(net4659),
    .S(_10260_),
    .X(_01846_));
 sky130_fd_sc_hd__clkbuf_1 _17606_ (.A(_01846_),
    .X(_00544_));
 sky130_fd_sc_hd__nor2_1 _17607_ (.A(net3875),
    .B(net4624),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _17608_ (.A(net3875),
    .B(net4624),
    .Y(_01848_));
 sky130_fd_sc_hd__or2b_1 _17609_ (.A(_01847_),
    .B_N(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__o21a_1 _17610_ (.A1(_01732_),
    .A2(_01735_),
    .B1(_01733_),
    .X(_01850_));
 sky130_fd_sc_hd__nor2_1 _17611_ (.A(_01849_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__a21o_1 _17612_ (.A1(_01849_),
    .A2(_01850_),
    .B1(_09845_),
    .X(_01852_));
 sky130_fd_sc_hd__or2b_1 _17613_ (.A(_01779_),
    .B_N(_01744_),
    .X(_01853_));
 sky130_fd_sc_hd__a21oi_2 _17614_ (.A1(_01756_),
    .A2(_01757_),
    .B1(_01754_),
    .Y(_01854_));
 sky130_fd_sc_hd__a21oi_2 _17615_ (.A1(_01777_),
    .A2(_01853_),
    .B1(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__and3_1 _17616_ (.A(_01777_),
    .B(_01853_),
    .C(_01854_),
    .X(_01856_));
 sky130_fd_sc_hd__nor2_1 _17617_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__a21o_1 _17618_ (.A1(_01758_),
    .A2(_01775_),
    .B1(_01773_),
    .X(_01858_));
 sky130_fd_sc_hd__or2b_1 _17619_ (.A(_01804_),
    .B_N(_01781_),
    .X(_01859_));
 sky130_fd_sc_hd__nor2_1 _17620_ (.A(_10190_),
    .B(_09225_),
    .Y(_01860_));
 sky130_fd_sc_hd__xnor2_1 _17621_ (.A(_01748_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _17622_ (.A(_08661_),
    .B(_09612_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_1 _17623_ (.A(_01861_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__or2_1 _17624_ (.A(_01861_),
    .B(_01862_),
    .X(_01864_));
 sky130_fd_sc_hd__nand2_1 _17625_ (.A(_01863_),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__a21oi_1 _17626_ (.A1(_01750_),
    .A2(_01751_),
    .B1(_01749_),
    .Y(_01866_));
 sky130_fd_sc_hd__nor2_1 _17627_ (.A(_01865_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__and2_1 _17628_ (.A(_01865_),
    .B(_01866_),
    .X(_01868_));
 sky130_fd_sc_hd__nor2_1 _17629_ (.A(_01867_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _17630_ (.A(_09373_),
    .B(_10289_),
    .Y(_01870_));
 sky130_fd_sc_hd__xor2_2 _17631_ (.A(_01869_),
    .B(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__o31ai_2 _17632_ (.A1(_10190_),
    .A2(_09116_),
    .A3(_01765_),
    .B1(_01763_),
    .Y(_01872_));
 sky130_fd_sc_hd__or3_1 _17633_ (.A(_01784_),
    .B(_01760_),
    .C(_01783_),
    .X(_01873_));
 sky130_fd_sc_hd__or2_1 _17634_ (.A(_10432_),
    .B(_08612_),
    .X(_01874_));
 sky130_fd_sc_hd__nor2_1 _17635_ (.A(_10186_),
    .B(_09060_),
    .Y(_01875_));
 sky130_fd_sc_hd__xnor2_1 _17636_ (.A(_01874_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__nor2_1 _17637_ (.A(_10163_),
    .B(_09114_),
    .Y(_01877_));
 sky130_fd_sc_hd__xnor2_1 _17638_ (.A(_01876_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__a21oi_1 _17639_ (.A1(_01873_),
    .A2(_01788_),
    .B1(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__and3_1 _17640_ (.A(_01873_),
    .B(_01788_),
    .C(_01878_),
    .X(_01880_));
 sky130_fd_sc_hd__nor2_1 _17641_ (.A(_01879_),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__xnor2_1 _17642_ (.A(_01872_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21oi_1 _17643_ (.A1(_01759_),
    .A2(_01770_),
    .B1(_01768_),
    .Y(_01883_));
 sky130_fd_sc_hd__nor2_1 _17644_ (.A(_01882_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__and2_1 _17645_ (.A(_01882_),
    .B(_01883_),
    .X(_01885_));
 sky130_fd_sc_hd__nor2_1 _17646_ (.A(_01884_),
    .B(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__xnor2_1 _17647_ (.A(_01871_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__a21o_1 _17648_ (.A1(_01802_),
    .A2(_01859_),
    .B1(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__nand3_1 _17649_ (.A(_01802_),
    .B(_01859_),
    .C(_01887_),
    .Y(_01889_));
 sky130_fd_sc_hd__nand2_1 _17650_ (.A(_01888_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__xnor2_1 _17651_ (.A(_01858_),
    .B(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__a21o_1 _17652_ (.A1(_01790_),
    .A2(_01800_),
    .B1(_01798_),
    .X(_01892_));
 sky130_fd_sc_hd__nand2_1 _17653_ (.A(_01807_),
    .B(_01812_),
    .Y(_01893_));
 sky130_fd_sc_hd__or2b_1 _17654_ (.A(_01813_),
    .B_N(_01806_),
    .X(_01894_));
 sky130_fd_sc_hd__or2_1 _17655_ (.A(_10062_),
    .B(_09181_),
    .X(_01895_));
 sky130_fd_sc_hd__or3_1 _17656_ (.A(_01784_),
    .B(_09040_),
    .C(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__o21ai_1 _17657_ (.A1(_01784_),
    .A2(_09040_),
    .B1(_01895_),
    .Y(_01897_));
 sky130_fd_sc_hd__and2_1 _17658_ (.A(_01896_),
    .B(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__nor2_1 _17659_ (.A(_01760_),
    .B(net8008),
    .Y(_01899_));
 sky130_fd_sc_hd__nand2_1 _17660_ (.A(_01898_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__or2_1 _17661_ (.A(_01898_),
    .B(_01899_),
    .X(_01901_));
 sky130_fd_sc_hd__and2_1 _17662_ (.A(_01900_),
    .B(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__nor2_1 _17663_ (.A(_08799_),
    .B(_10096_),
    .Y(_01903_));
 sky130_fd_sc_hd__nor2_1 _17664_ (.A(_10327_),
    .B(_10220_),
    .Y(_01904_));
 sky130_fd_sc_hd__xnor2_1 _17665_ (.A(_01903_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__or2_1 _17666_ (.A(_01794_),
    .B(_09664_),
    .X(_01906_));
 sky130_fd_sc_hd__xnor2_1 _17667_ (.A(_01905_),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _17668_ (.A(_01791_),
    .B(_01792_),
    .Y(_01908_));
 sky130_fd_sc_hd__o31a_1 _17669_ (.A1(_01794_),
    .A2(_09403_),
    .A3(_01793_),
    .B1(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__nor2_1 _17670_ (.A(_01907_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__and2_1 _17671_ (.A(_01907_),
    .B(_01909_),
    .X(_01911_));
 sky130_fd_sc_hd__nor2_1 _17672_ (.A(_01910_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__xnor2_1 _17673_ (.A(_01902_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__a21o_1 _17674_ (.A1(_01893_),
    .A2(_01894_),
    .B1(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__nand3_1 _17675_ (.A(_01893_),
    .B(_01894_),
    .C(_01913_),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _17676_ (.A(_01914_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_1 _17677_ (.A(_01892_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__a21bo_1 _17678_ (.A1(_01808_),
    .A2(_01811_),
    .B1_N(_01809_),
    .X(_01918_));
 sky130_fd_sc_hd__or2_1 _17679_ (.A(_09272_),
    .B(_10346_),
    .X(_01919_));
 sky130_fd_sc_hd__or3_1 _17680_ (.A(_08918_),
    .B(_10211_),
    .C(_09970_),
    .X(_01920_));
 sky130_fd_sc_hd__a21oi_1 _17681_ (.A1(_08918_),
    .A2(_10211_),
    .B1(_01693_),
    .Y(_01921_));
 sky130_fd_sc_hd__nand2_2 _17682_ (.A(_01920_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__xor2_1 _17683_ (.A(_01919_),
    .B(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__xnor2_1 _17684_ (.A(_01807_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__xnor2_1 _17685_ (.A(_01918_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__xnor2_1 _17686_ (.A(_01818_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__a21oi_1 _17687_ (.A1(_01815_),
    .A2(_01819_),
    .B1(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__and3_1 _17688_ (.A(_01815_),
    .B(_01819_),
    .C(_01926_),
    .X(_01928_));
 sky130_fd_sc_hd__nor2_1 _17689_ (.A(_01927_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__xnor2_1 _17690_ (.A(_01917_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__a21oi_1 _17691_ (.A1(_01805_),
    .A2(_01825_),
    .B1(_01823_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _17692_ (.A(_01930_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__and2_1 _17693_ (.A(_01930_),
    .B(_01931_),
    .X(_01933_));
 sky130_fd_sc_hd__nor2_1 _17694_ (.A(_01932_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__xnor2_1 _17695_ (.A(_01891_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__a21oi_1 _17696_ (.A1(_01780_),
    .A2(_01830_),
    .B1(_01828_),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _17697_ (.A(_01935_),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__nand2_1 _17698_ (.A(_01935_),
    .B(_01936_),
    .Y(_01938_));
 sky130_fd_sc_hd__and2b_1 _17699_ (.A_N(_01937_),
    .B(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__xnor2_1 _17700_ (.A(_01857_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__nor2_1 _17701_ (.A(_01831_),
    .B(_01833_),
    .Y(_01941_));
 sky130_fd_sc_hd__a21oi_1 _17702_ (.A1(_01743_),
    .A2(_01834_),
    .B1(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__xor2_1 _17703_ (.A(_01940_),
    .B(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_01741_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__nor2_1 _17705_ (.A(_01835_),
    .B(_01836_),
    .Y(_01945_));
 sky130_fd_sc_hd__a21oi_1 _17706_ (.A1(_10390_),
    .A2(_01837_),
    .B1(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__or2_1 _17707_ (.A(_01944_),
    .B(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__nand2_1 _17708_ (.A(_01944_),
    .B(_01946_),
    .Y(_01948_));
 sky130_fd_sc_hd__nand2_2 _17709_ (.A(_01947_),
    .B(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__a311o_1 _17710_ (.A1(_01737_),
    .A2(_01738_),
    .A3(_01838_),
    .B1(_01720_),
    .C1(_01718_),
    .X(_01950_));
 sky130_fd_sc_hd__o311a_4 _17711_ (.A1(_01723_),
    .A2(_01726_),
    .A3(_01841_),
    .B1(_01950_),
    .C1(_01840_),
    .X(_01951_));
 sky130_fd_sc_hd__o21ai_1 _17712_ (.A1(_01949_),
    .A2(_01951_),
    .B1(_08103_),
    .Y(_01952_));
 sky130_fd_sc_hd__a21o_1 _17713_ (.A1(_01949_),
    .A2(_01951_),
    .B1(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__o21ai_1 _17714_ (.A1(_01851_),
    .A2(_01852_),
    .B1(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__mux2_1 _17715_ (.A0(_01954_),
    .A1(net3875),
    .S(_10260_),
    .X(_01955_));
 sky130_fd_sc_hd__clkbuf_1 _17716_ (.A(_01955_),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _17717_ (.A(net4723),
    .B(net4520),
    .Y(_01956_));
 sky130_fd_sc_hd__nand2_1 _17718_ (.A(net4723),
    .B(net4520),
    .Y(_01957_));
 sky130_fd_sc_hd__or2b_1 _17719_ (.A(_01956_),
    .B_N(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__o21a_1 _17720_ (.A1(_01847_),
    .A2(_01850_),
    .B1(_01848_),
    .X(_01959_));
 sky130_fd_sc_hd__nor2_1 _17721_ (.A(_01958_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__a21o_1 _17722_ (.A1(_01958_),
    .A2(_01959_),
    .B1(_09845_),
    .X(_01961_));
 sky130_fd_sc_hd__or2_1 _17723_ (.A(_01940_),
    .B(_01942_),
    .X(_01962_));
 sky130_fd_sc_hd__nand2_1 _17724_ (.A(_01741_),
    .B(_01943_),
    .Y(_01963_));
 sky130_fd_sc_hd__or2b_1 _17725_ (.A(_01890_),
    .B_N(_01858_),
    .X(_01964_));
 sky130_fd_sc_hd__a21oi_2 _17726_ (.A1(_01869_),
    .A2(_01870_),
    .B1(_01867_),
    .Y(_01965_));
 sky130_fd_sc_hd__a21oi_2 _17727_ (.A1(_01888_),
    .A2(_01964_),
    .B1(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__and3_1 _17728_ (.A(_01888_),
    .B(_01964_),
    .C(_01965_),
    .X(_01967_));
 sky130_fd_sc_hd__nor2_1 _17729_ (.A(_01966_),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__a21o_1 _17730_ (.A1(_01871_),
    .A2(_01886_),
    .B1(_01884_),
    .X(_01969_));
 sky130_fd_sc_hd__or2b_1 _17731_ (.A(_01916_),
    .B_N(_01892_),
    .X(_01970_));
 sky130_fd_sc_hd__nor2_1 _17732_ (.A(_10408_),
    .B(_09345_),
    .Y(_01971_));
 sky130_fd_sc_hd__nor2_1 _17733_ (.A(_10163_),
    .B(net4908),
    .Y(_01972_));
 sky130_fd_sc_hd__xnor2_1 _17734_ (.A(_01971_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_1 _17735_ (.A(_09915_),
    .B(_09612_),
    .Y(_01974_));
 sky130_fd_sc_hd__xor2_1 _17736_ (.A(_01973_),
    .B(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__o31a_1 _17737_ (.A1(_10190_),
    .A2(_09225_),
    .A3(_01748_),
    .B1(_01863_),
    .X(_01976_));
 sky130_fd_sc_hd__nor2_1 _17738_ (.A(_01975_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__and2_1 _17739_ (.A(_01975_),
    .B(_01976_),
    .X(_01978_));
 sky130_fd_sc_hd__nor2_1 _17740_ (.A(_01977_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _17741_ (.A(_08167_),
    .B(_10289_),
    .Y(_01980_));
 sky130_fd_sc_hd__xor2_1 _17742_ (.A(_01979_),
    .B(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__nand2_1 _17743_ (.A(_08465_),
    .B(_09354_),
    .Y(_01982_));
 sky130_fd_sc_hd__o2bb2ai_2 _17744_ (.A1_N(_01876_),
    .A2_N(_01877_),
    .B1(_01982_),
    .B2(_01762_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _17745_ (.A(_01760_),
    .B(_08612_),
    .Y(_01984_));
 sky130_fd_sc_hd__xnor2_1 _17746_ (.A(_01982_),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__nor2_1 _17747_ (.A(_10186_),
    .B(_09114_),
    .Y(_01986_));
 sky130_fd_sc_hd__xnor2_1 _17748_ (.A(_01985_),
    .B(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__a21oi_1 _17749_ (.A1(_01896_),
    .A2(_01900_),
    .B1(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__and3_1 _17750_ (.A(_01896_),
    .B(_01900_),
    .C(_01987_),
    .X(_01989_));
 sky130_fd_sc_hd__nor2_1 _17751_ (.A(_01988_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__xnor2_1 _17752_ (.A(_01983_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__a21oi_1 _17753_ (.A1(_01872_),
    .A2(_01881_),
    .B1(_01879_),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _17754_ (.A(_01991_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__and2_1 _17755_ (.A(_01991_),
    .B(_01992_),
    .X(_01994_));
 sky130_fd_sc_hd__nor2_1 _17756_ (.A(_01993_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__xnor2_1 _17757_ (.A(_01981_),
    .B(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__a21o_1 _17758_ (.A1(_01914_),
    .A2(_01970_),
    .B1(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__nand3_1 _17759_ (.A(_01914_),
    .B(_01970_),
    .C(_01996_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_1 _17760_ (.A(_01997_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__xnor2_2 _17761_ (.A(_01969_),
    .B(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__o21ai_1 _17762_ (.A1(_01919_),
    .A2(_01922_),
    .B1(_01920_),
    .Y(_02001_));
 sky130_fd_sc_hd__nor2_1 _17763_ (.A(_09272_),
    .B(_01693_),
    .Y(_02002_));
 sky130_fd_sc_hd__mux2_2 _17764_ (.A0(_09272_),
    .A1(_02002_),
    .S(_01922_),
    .X(_02003_));
 sky130_fd_sc_hd__xnor2_4 _17765_ (.A(_01807_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__xnor2_1 _17766_ (.A(_02001_),
    .B(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _17767_ (.A(_01818_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__or2_1 _17768_ (.A(_01818_),
    .B(_02005_),
    .X(_02007_));
 sky130_fd_sc_hd__nand2_1 _17769_ (.A(_02006_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__a21boi_1 _17770_ (.A1(_01818_),
    .A2(_01925_),
    .B1_N(_01815_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _17771_ (.A(_02008_),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__and2_1 _17772_ (.A(_02008_),
    .B(_02009_),
    .X(_02011_));
 sky130_fd_sc_hd__nor2_1 _17773_ (.A(_02010_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__a21o_1 _17774_ (.A1(_01902_),
    .A2(_01912_),
    .B1(_01910_),
    .X(_02013_));
 sky130_fd_sc_hd__nand2_1 _17775_ (.A(_01807_),
    .B(_01923_),
    .Y(_02014_));
 sky130_fd_sc_hd__or2b_1 _17776_ (.A(_01924_),
    .B_N(_01918_),
    .X(_02015_));
 sky130_fd_sc_hd__nor2_1 _17777_ (.A(_10062_),
    .B(_09410_),
    .Y(_02016_));
 sky130_fd_sc_hd__nor2_1 _17778_ (.A(_01784_),
    .B(_09181_),
    .Y(_02017_));
 sky130_fd_sc_hd__xnor2_1 _17779_ (.A(_02016_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__or3_1 _17780_ (.A(_09040_),
    .B(net8008),
    .C(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__o21ai_1 _17781_ (.A1(_09040_),
    .A2(net8008),
    .B1(_02018_),
    .Y(_02020_));
 sky130_fd_sc_hd__and2_1 _17782_ (.A(_02019_),
    .B(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__nor2_1 _17783_ (.A(_08799_),
    .B(_10220_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_1 _17784_ (.A(_10327_),
    .B(_10346_),
    .Y(_02023_));
 sky130_fd_sc_hd__xnor2_1 _17785_ (.A(_02022_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__nor2_1 _17786_ (.A(_01794_),
    .B(_10096_),
    .Y(_02025_));
 sky130_fd_sc_hd__xor2_1 _17787_ (.A(_02024_),
    .B(_02025_),
    .X(_02026_));
 sky130_fd_sc_hd__nand2_1 _17788_ (.A(_01903_),
    .B(_01904_),
    .Y(_02027_));
 sky130_fd_sc_hd__o31a_1 _17789_ (.A1(_01794_),
    .A2(_09664_),
    .A3(_01905_),
    .B1(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__xor2_1 _17790_ (.A(_02026_),
    .B(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__xnor2_1 _17791_ (.A(_02021_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__a21o_1 _17792_ (.A1(_02014_),
    .A2(_02015_),
    .B1(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__nand3_1 _17793_ (.A(_02014_),
    .B(_02015_),
    .C(_02030_),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_1 _17794_ (.A(_02031_),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__xnor2_2 _17795_ (.A(_02013_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__xnor2_1 _17796_ (.A(_02012_),
    .B(_02034_),
    .Y(_02035_));
 sky130_fd_sc_hd__a21oi_1 _17797_ (.A1(_01917_),
    .A2(_01929_),
    .B1(_01927_),
    .Y(_02036_));
 sky130_fd_sc_hd__nor2_1 _17798_ (.A(_02035_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__and2_1 _17799_ (.A(_02035_),
    .B(_02036_),
    .X(_02038_));
 sky130_fd_sc_hd__nor2_1 _17800_ (.A(_02037_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__xnor2_2 _17801_ (.A(_02000_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__a21oi_2 _17802_ (.A1(_01891_),
    .A2(_01934_),
    .B1(_01932_),
    .Y(_02041_));
 sky130_fd_sc_hd__xor2_2 _17803_ (.A(_02040_),
    .B(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__xnor2_1 _17804_ (.A(_01968_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21oi_1 _17805_ (.A1(_01857_),
    .A2(_01938_),
    .B1(_01937_),
    .Y(_02044_));
 sky130_fd_sc_hd__xor2_1 _17806_ (.A(_02043_),
    .B(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__xnor2_1 _17807_ (.A(_01855_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__a21oi_1 _17808_ (.A1(_01962_),
    .A2(_01963_),
    .B1(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__and3_1 _17809_ (.A(_01962_),
    .B(_01963_),
    .C(_02046_),
    .X(_02048_));
 sky130_fd_sc_hd__or2_2 _17810_ (.A(_02047_),
    .B(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__o21a_1 _17811_ (.A1(_01949_),
    .A2(_01951_),
    .B1(_01947_),
    .X(_02050_));
 sky130_fd_sc_hd__o21ai_1 _17812_ (.A1(_02049_),
    .A2(_02050_),
    .B1(_08103_),
    .Y(_02051_));
 sky130_fd_sc_hd__a21o_1 _17813_ (.A1(_02049_),
    .A2(_02050_),
    .B1(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__o21ai_1 _17814_ (.A1(_01960_),
    .A2(_01961_),
    .B1(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__mux2_1 _17815_ (.A0(_02053_),
    .A1(net4723),
    .S(_10260_),
    .X(_02054_));
 sky130_fd_sc_hd__clkbuf_1 _17816_ (.A(_02054_),
    .X(_00546_));
 sky130_fd_sc_hd__or2_1 _17817_ (.A(net4655),
    .B(net4756),
    .X(_02055_));
 sky130_fd_sc_hd__nand2_1 _17818_ (.A(net4655),
    .B(net4756),
    .Y(_02056_));
 sky130_fd_sc_hd__nand2_1 _17819_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__o21ai_1 _17820_ (.A1(_01956_),
    .A2(_01959_),
    .B1(_01957_),
    .Y(_02058_));
 sky130_fd_sc_hd__xnor2_1 _17821_ (.A(_02057_),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__or2b_1 _17822_ (.A(_01999_),
    .B_N(_01969_),
    .X(_02060_));
 sky130_fd_sc_hd__a21oi_1 _17823_ (.A1(_01979_),
    .A2(_01980_),
    .B1(_01977_),
    .Y(_02061_));
 sky130_fd_sc_hd__a21oi_2 _17824_ (.A1(_01997_),
    .A2(_02060_),
    .B1(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__and3_1 _17825_ (.A(_01997_),
    .B(_02060_),
    .C(_02061_),
    .X(_02063_));
 sky130_fd_sc_hd__nor2_1 _17826_ (.A(_02062_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__o21a_1 _17827_ (.A1(_09272_),
    .A2(_01922_),
    .B1(_01920_),
    .X(_02065_));
 sky130_fd_sc_hd__xor2_2 _17828_ (.A(_02004_),
    .B(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__xnor2_1 _17829_ (.A(_01818_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__a21o_1 _17830_ (.A1(_01815_),
    .A2(_02006_),
    .B1(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__nand3_1 _17831_ (.A(_01815_),
    .B(_02006_),
    .C(_02067_),
    .Y(_02069_));
 sky130_fd_sc_hd__and2_1 _17832_ (.A(_02068_),
    .B(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__nor2_1 _17833_ (.A(_02026_),
    .B(_02028_),
    .Y(_02071_));
 sky130_fd_sc_hd__a21o_1 _17834_ (.A1(_02021_),
    .A2(_02029_),
    .B1(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__nand2_1 _17835_ (.A(_01807_),
    .B(_02003_),
    .Y(_02073_));
 sky130_fd_sc_hd__or2b_1 _17836_ (.A(_02004_),
    .B_N(_02001_),
    .X(_02074_));
 sky130_fd_sc_hd__nand2_1 _17837_ (.A(_02073_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__or2_1 _17838_ (.A(_10062_),
    .B(_09540_),
    .X(_02076_));
 sky130_fd_sc_hd__nor2_1 _17839_ (.A(_01784_),
    .B(_09410_),
    .Y(_02077_));
 sky130_fd_sc_hd__xnor2_1 _17840_ (.A(_02076_),
    .B(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__nor2_1 _17841_ (.A(net8008),
    .B(_09181_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _17842_ (.A(_02078_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__or4_1 _17843_ (.A(_10327_),
    .B(_08799_),
    .C(_01693_),
    .D(_09976_),
    .X(_02081_));
 sky130_fd_sc_hd__o22ai_1 _17844_ (.A1(_10327_),
    .A2(_01693_),
    .B1(_10346_),
    .B2(_08799_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _17845_ (.A(_02081_),
    .B(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_1 _17846_ (.A(_01794_),
    .B(_10220_),
    .Y(_02084_));
 sky130_fd_sc_hd__xor2_1 _17847_ (.A(_02083_),
    .B(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__nand2_1 _17848_ (.A(_02022_),
    .B(_02023_),
    .Y(_02086_));
 sky130_fd_sc_hd__o31a_1 _17849_ (.A1(_01794_),
    .A2(_10096_),
    .A3(_02024_),
    .B1(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__xor2_1 _17850_ (.A(_02085_),
    .B(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__xnor2_1 _17851_ (.A(_02080_),
    .B(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__xnor2_1 _17852_ (.A(_02075_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__xnor2_1 _17853_ (.A(_02072_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2_1 _17854_ (.A(_02070_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__or2_1 _17855_ (.A(_02070_),
    .B(_02091_),
    .X(_02093_));
 sky130_fd_sc_hd__nand2_1 _17856_ (.A(_02092_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__a21oi_1 _17857_ (.A1(_02012_),
    .A2(_02034_),
    .B1(_02010_),
    .Y(_02095_));
 sky130_fd_sc_hd__xor2_1 _17858_ (.A(_02094_),
    .B(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__a21o_1 _17859_ (.A1(_01981_),
    .A2(_01995_),
    .B1(_01993_),
    .X(_02097_));
 sky130_fd_sc_hd__or2b_1 _17860_ (.A(_02033_),
    .B_N(_02013_),
    .X(_02098_));
 sky130_fd_sc_hd__or2_1 _17861_ (.A(_08472_),
    .B(_09225_),
    .X(_02099_));
 sky130_fd_sc_hd__or3_1 _17862_ (.A(_10163_),
    .B(net4913),
    .C(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__o21ai_1 _17863_ (.A1(_10163_),
    .A2(net4913),
    .B1(_02099_),
    .Y(_02101_));
 sky130_fd_sc_hd__nand2_1 _17864_ (.A(_02100_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _17865_ (.A(_10190_),
    .B(_09612_),
    .Y(_02103_));
 sky130_fd_sc_hd__xor2_1 _17866_ (.A(_02102_),
    .B(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__nand2_1 _17867_ (.A(_01971_),
    .B(_01972_),
    .Y(_02105_));
 sky130_fd_sc_hd__o31a_1 _17868_ (.A1(_09915_),
    .A2(_09612_),
    .A3(_01973_),
    .B1(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__nor2_1 _17869_ (.A(_02104_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__and2_1 _17870_ (.A(_02104_),
    .B(_02106_),
    .X(_02108_));
 sky130_fd_sc_hd__nor2_1 _17871_ (.A(_02107_),
    .B(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__and2_1 _17872_ (.A(_09915_),
    .B(net4891),
    .X(_02110_));
 sky130_fd_sc_hd__xor2_1 _17873_ (.A(_02109_),
    .B(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__or3_1 _17874_ (.A(_01760_),
    .B(_08612_),
    .C(_01982_),
    .X(_02112_));
 sky130_fd_sc_hd__a21bo_1 _17875_ (.A1(_01985_),
    .A2(_01986_),
    .B1_N(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(_02016_),
    .B(_02017_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _17877_ (.A(_01760_),
    .B(_09060_),
    .Y(_02115_));
 sky130_fd_sc_hd__nor2_1 _17878_ (.A(_09040_),
    .B(_08612_),
    .Y(_02116_));
 sky130_fd_sc_hd__xnor2_1 _17879_ (.A(_02115_),
    .B(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__or3_1 _17880_ (.A(_10432_),
    .B(_09114_),
    .C(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__o21ai_1 _17881_ (.A1(_10432_),
    .A2(_09114_),
    .B1(_02117_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _17882_ (.A(_02118_),
    .B(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21oi_1 _17883_ (.A1(_02114_),
    .A2(_02019_),
    .B1(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__and3_1 _17884_ (.A(_02114_),
    .B(_02019_),
    .C(_02120_),
    .X(_02122_));
 sky130_fd_sc_hd__nor2_1 _17885_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__xnor2_1 _17886_ (.A(_02113_),
    .B(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__a21oi_1 _17887_ (.A1(_01983_),
    .A2(_01990_),
    .B1(_01988_),
    .Y(_02125_));
 sky130_fd_sc_hd__nor2_1 _17888_ (.A(_02124_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__and2_1 _17889_ (.A(_02124_),
    .B(_02125_),
    .X(_02127_));
 sky130_fd_sc_hd__nor2_1 _17890_ (.A(_02126_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__xnor2_1 _17891_ (.A(_02111_),
    .B(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__a21oi_1 _17892_ (.A1(_02031_),
    .A2(_02098_),
    .B1(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__and3_1 _17893_ (.A(_02031_),
    .B(_02098_),
    .C(_02129_),
    .X(_02131_));
 sky130_fd_sc_hd__or2_1 _17894_ (.A(_02130_),
    .B(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__xnor2_1 _17895_ (.A(_02097_),
    .B(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand2_1 _17896_ (.A(_02096_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__or2_1 _17897_ (.A(_02096_),
    .B(_02133_),
    .X(_02135_));
 sky130_fd_sc_hd__nand2_1 _17898_ (.A(_02134_),
    .B(_02135_),
    .Y(_02136_));
 sky130_fd_sc_hd__a21oi_1 _17899_ (.A1(_02000_),
    .A2(_02039_),
    .B1(_02037_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _17900_ (.A(_02136_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__and2_1 _17901_ (.A(_02136_),
    .B(_02137_),
    .X(_02139_));
 sky130_fd_sc_hd__nor2_1 _17902_ (.A(_02138_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__xnor2_1 _17903_ (.A(_02064_),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nor2_1 _17904_ (.A(_02040_),
    .B(_02041_),
    .Y(_02142_));
 sky130_fd_sc_hd__a21oi_2 _17905_ (.A1(_01968_),
    .A2(_02042_),
    .B1(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__xor2_1 _17906_ (.A(_02141_),
    .B(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__xnor2_1 _17907_ (.A(_01966_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nor2_1 _17908_ (.A(_02043_),
    .B(_02044_),
    .Y(_02146_));
 sky130_fd_sc_hd__a21oi_2 _17909_ (.A1(_01855_),
    .A2(_02045_),
    .B1(_02146_),
    .Y(_02147_));
 sky130_fd_sc_hd__or2_1 _17910_ (.A(_02145_),
    .B(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__nand2_1 _17911_ (.A(_02145_),
    .B(_02147_),
    .Y(_02149_));
 sky130_fd_sc_hd__and2_1 _17912_ (.A(_02148_),
    .B(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__a21o_1 _17913_ (.A1(_01962_),
    .A2(_01963_),
    .B1(_02046_),
    .X(_02151_));
 sky130_fd_sc_hd__a21o_1 _17914_ (.A1(_01947_),
    .A2(_02151_),
    .B1(_02048_),
    .X(_02152_));
 sky130_fd_sc_hd__o31ai_4 _17915_ (.A1(_01949_),
    .A2(_01951_),
    .A3(_02049_),
    .B1(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__a21oi_1 _17916_ (.A1(_02150_),
    .A2(_02153_),
    .B1(net90),
    .Y(_02154_));
 sky130_fd_sc_hd__o21a_1 _17917_ (.A1(_02150_),
    .A2(_02153_),
    .B1(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__a21o_1 _17918_ (.A1(_09788_),
    .A2(_02059_),
    .B1(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__mux2_1 _17919_ (.A0(_02156_),
    .A1(net4655),
    .S(_10260_),
    .X(_02157_));
 sky130_fd_sc_hd__clkbuf_1 _17920_ (.A(_02157_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _17921_ (.A(_02141_),
    .B(_02143_),
    .X(_02158_));
 sky130_fd_sc_hd__nand2_1 _17922_ (.A(_01966_),
    .B(_02144_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _17923_ (.A(_01816_),
    .B(_02066_),
    .Y(_02160_));
 sky130_fd_sc_hd__and2b_1 _17924_ (.A_N(_01815_),
    .B(_02066_),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_1 _17925_ (.A(_02160_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__or2b_1 _17926_ (.A(_02080_),
    .B_N(_02088_),
    .X(_02163_));
 sky130_fd_sc_hd__o21a_1 _17927_ (.A1(_02085_),
    .A2(_02087_),
    .B1(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__o21ai_2 _17928_ (.A1(_02004_),
    .A2(_02065_),
    .B1(_02073_),
    .Y(_02165_));
 sky130_fd_sc_hd__or2_1 _17929_ (.A(_10062_),
    .B(_09666_),
    .X(_02166_));
 sky130_fd_sc_hd__nor2_1 _17930_ (.A(_01784_),
    .B(_09540_),
    .Y(_02167_));
 sky130_fd_sc_hd__xnor2_1 _17931_ (.A(_02166_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__nor2_1 _17932_ (.A(net8008),
    .B(_09410_),
    .Y(_02169_));
 sky130_fd_sc_hd__nand2_1 _17933_ (.A(_02168_),
    .B(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__or2_1 _17934_ (.A(_02168_),
    .B(_02169_),
    .X(_02171_));
 sky130_fd_sc_hd__and2_1 _17935_ (.A(_02170_),
    .B(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__o31a_1 _17936_ (.A1(_01794_),
    .A2(_10220_),
    .A3(_02083_),
    .B1(_02081_),
    .X(_02173_));
 sky130_fd_sc_hd__a21o_1 _17937_ (.A1(_10327_),
    .A2(_08799_),
    .B1(_01693_),
    .X(_02174_));
 sky130_fd_sc_hd__nor3_1 _17938_ (.A(_10327_),
    .B(_08799_),
    .C(_01693_),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _17939_ (.A(_02174_),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _17940_ (.A(_01794_),
    .B(_10346_),
    .Y(_02177_));
 sky130_fd_sc_hd__xnor2_1 _17941_ (.A(_02176_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__xor2_1 _17942_ (.A(_02173_),
    .B(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__xor2_1 _17943_ (.A(_02172_),
    .B(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__and2_1 _17944_ (.A(_02165_),
    .B(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__nor2_1 _17945_ (.A(_02165_),
    .B(_02180_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_1 _17946_ (.A(_02181_),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__xnor2_1 _17947_ (.A(_02164_),
    .B(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__xnor2_1 _17948_ (.A(_02162_),
    .B(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__a21o_1 _17949_ (.A1(_02068_),
    .A2(_02092_),
    .B1(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__nand3_1 _17950_ (.A(_02068_),
    .B(_02092_),
    .C(_02185_),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _17951_ (.A(_02186_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__a21o_1 _17952_ (.A1(_02111_),
    .A2(_02128_),
    .B1(_02126_),
    .X(_02189_));
 sky130_fd_sc_hd__or2b_1 _17953_ (.A(_02090_),
    .B_N(_02072_),
    .X(_02190_));
 sky130_fd_sc_hd__a21bo_1 _17954_ (.A1(_02075_),
    .A2(_02089_),
    .B1_N(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__o22a_1 _17955_ (.A1(_10316_),
    .A2(_09225_),
    .B1(_09345_),
    .B2(_08472_),
    .X(_02192_));
 sky130_fd_sc_hd__or3_1 _17956_ (.A(_10316_),
    .B(_09345_),
    .C(_02099_),
    .X(_02193_));
 sky130_fd_sc_hd__or2b_1 _17957_ (.A(_02192_),
    .B_N(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__or3b_1 _17958_ (.A(_09413_),
    .B(_10163_),
    .C_N(net7837),
    .X(_02195_));
 sky130_fd_sc_hd__xnor2_1 _17959_ (.A(_02194_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__o31a_1 _17960_ (.A1(_10190_),
    .A2(_09612_),
    .A3(_02102_),
    .B1(_02100_),
    .X(_02197_));
 sky130_fd_sc_hd__xnor2_1 _17961_ (.A(_02196_),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__nand2_1 _17962_ (.A(_10190_),
    .B(net7818),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _17963_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__a21bo_1 _17964_ (.A1(_02115_),
    .A2(_02116_),
    .B1_N(_02118_),
    .X(_02201_));
 sky130_fd_sc_hd__or3_1 _17965_ (.A(_01784_),
    .B(_09410_),
    .C(_02076_),
    .X(_02202_));
 sky130_fd_sc_hd__a21bo_1 _17966_ (.A1(_02078_),
    .A2(_02079_),
    .B1_N(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__nor2_1 _17967_ (.A(_09040_),
    .B(_09060_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _17968_ (.A(_08612_),
    .B(_09181_),
    .Y(_02205_));
 sky130_fd_sc_hd__xnor2_1 _17969_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__nor2_1 _17970_ (.A(_01760_),
    .B(_09114_),
    .Y(_02207_));
 sky130_fd_sc_hd__xnor2_1 _17971_ (.A(_02206_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__nand2_1 _17972_ (.A(_02203_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__or2_1 _17973_ (.A(_02203_),
    .B(_02208_),
    .X(_02210_));
 sky130_fd_sc_hd__and2_1 _17974_ (.A(_02209_),
    .B(_02210_),
    .X(_02211_));
 sky130_fd_sc_hd__xnor2_2 _17975_ (.A(_02201_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__a21oi_1 _17976_ (.A1(_02113_),
    .A2(_02123_),
    .B1(_02121_),
    .Y(_02213_));
 sky130_fd_sc_hd__xor2_1 _17977_ (.A(_02212_),
    .B(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__xnor2_1 _17978_ (.A(_02200_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__xor2_1 _17979_ (.A(_02191_),
    .B(_02215_),
    .X(_02216_));
 sky130_fd_sc_hd__and2_1 _17980_ (.A(_02189_),
    .B(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__nor2_1 _17981_ (.A(_02189_),
    .B(_02216_),
    .Y(_02218_));
 sky130_fd_sc_hd__nor2_1 _17982_ (.A(_02217_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__xor2_1 _17983_ (.A(_02188_),
    .B(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__o21a_1 _17984_ (.A1(_02094_),
    .A2(_02095_),
    .B1(_02134_),
    .X(_02221_));
 sky130_fd_sc_hd__xor2_1 _17985_ (.A(_02220_),
    .B(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__and2b_1 _17986_ (.A_N(_02132_),
    .B(_02097_),
    .X(_02223_));
 sky130_fd_sc_hd__a21oi_1 _17987_ (.A1(_02109_),
    .A2(_02110_),
    .B1(_02107_),
    .Y(_02224_));
 sky130_fd_sc_hd__o21ba_1 _17988_ (.A1(_02130_),
    .A2(_02223_),
    .B1_N(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__or3b_1 _17989_ (.A(_02130_),
    .B(_02223_),
    .C_N(_02224_),
    .X(_02226_));
 sky130_fd_sc_hd__and2b_1 _17990_ (.A_N(_02225_),
    .B(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__nand2_1 _17991_ (.A(_02222_),
    .B(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__or2_1 _17992_ (.A(_02222_),
    .B(_02227_),
    .X(_02229_));
 sky130_fd_sc_hd__nand2_1 _17993_ (.A(_02228_),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__a21oi_1 _17994_ (.A1(_02064_),
    .A2(_02140_),
    .B1(_02138_),
    .Y(_02231_));
 sky130_fd_sc_hd__xor2_1 _17995_ (.A(_02230_),
    .B(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__xnor2_1 _17996_ (.A(_02062_),
    .B(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__a21oi_1 _17997_ (.A1(_02158_),
    .A2(_02159_),
    .B1(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__and3_1 _17998_ (.A(_02158_),
    .B(_02159_),
    .C(_02233_),
    .X(_02235_));
 sky130_fd_sc_hd__nor2_1 _17999_ (.A(_02234_),
    .B(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__a21bo_1 _18000_ (.A1(_02150_),
    .A2(_02153_),
    .B1_N(_02148_),
    .X(_02237_));
 sky130_fd_sc_hd__or2_1 _18001_ (.A(_02236_),
    .B(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__a21oi_2 _18002_ (.A1(_02236_),
    .A2(_02237_),
    .B1(net90),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_1 _18003_ (.A(net4762),
    .B(net4388),
    .Y(_02240_));
 sky130_fd_sc_hd__or2_1 _18004_ (.A(net4762),
    .B(net4388),
    .X(_02241_));
 sky130_fd_sc_hd__nand2_1 _18005_ (.A(_02240_),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__a21bo_1 _18006_ (.A1(_02055_),
    .A2(_02058_),
    .B1_N(_02056_),
    .X(_02243_));
 sky130_fd_sc_hd__xnor2_1 _18007_ (.A(_02242_),
    .B(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__clkbuf_8 _18008_ (.A(net89),
    .X(_02245_));
 sky130_fd_sc_hd__a22o_1 _18009_ (.A1(_02238_),
    .A2(_02239_),
    .B1(_02244_),
    .B2(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_2 _18010_ (.A0(_02246_),
    .A1(net4762),
    .S(_10260_),
    .X(_02247_));
 sky130_fd_sc_hd__clkbuf_1 _18011_ (.A(_02247_),
    .X(_00548_));
 sky130_fd_sc_hd__a21bo_1 _18012_ (.A1(_02241_),
    .A2(_02243_),
    .B1_N(_02240_),
    .X(_02248_));
 sky130_fd_sc_hd__xor2_1 _18013_ (.A(net4742),
    .B(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__nor2_1 _18014_ (.A(net4622),
    .B(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21o_1 _18015_ (.A1(net4622),
    .A2(_02249_),
    .B1(_09845_),
    .X(_02251_));
 sky130_fd_sc_hd__a21o_1 _18016_ (.A1(_02158_),
    .A2(_02159_),
    .B1(_02233_),
    .X(_02252_));
 sky130_fd_sc_hd__a21oi_1 _18017_ (.A1(_02148_),
    .A2(_02252_),
    .B1(_02235_),
    .Y(_02253_));
 sky130_fd_sc_hd__a31o_1 _18018_ (.A1(_02150_),
    .A2(_02153_),
    .A3(_02236_),
    .B1(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__nor2_1 _18019_ (.A(_02230_),
    .B(_02231_),
    .Y(_02255_));
 sky130_fd_sc_hd__a21oi_1 _18020_ (.A1(_02062_),
    .A2(_02232_),
    .B1(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__o22a_1 _18021_ (.A1(_02196_),
    .A2(_02197_),
    .B1(_02198_),
    .B2(_02199_),
    .X(_02257_));
 sky130_fd_sc_hd__xnor2_1 _18022_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__o21a_1 _18023_ (.A1(_02220_),
    .A2(_02221_),
    .B1(_02228_),
    .X(_02259_));
 sky130_fd_sc_hd__o21bai_1 _18024_ (.A1(_02174_),
    .A2(_02177_),
    .B1_N(_02175_),
    .Y(_02260_));
 sky130_fd_sc_hd__a21oi_1 _18025_ (.A1(_02191_),
    .A2(_02215_),
    .B1(_02217_),
    .Y(_02261_));
 sky130_fd_sc_hd__o31a_1 _18026_ (.A1(_02188_),
    .A2(_02217_),
    .A3(_02218_),
    .B1(_02186_),
    .X(_02262_));
 sky130_fd_sc_hd__xnor2_1 _18027_ (.A(_02261_),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__xnor2_1 _18028_ (.A(_02260_),
    .B(_02263_),
    .Y(_02264_));
 sky130_fd_sc_hd__o21ba_1 _18029_ (.A1(_02160_),
    .A2(_02184_),
    .B1_N(_02161_),
    .X(_02265_));
 sky130_fd_sc_hd__xnor2_1 _18030_ (.A(_02165_),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_1 _18031_ (.A(_02173_),
    .B(_02178_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21oi_1 _18032_ (.A1(_02172_),
    .A2(_02179_),
    .B1(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__nor2_1 _18033_ (.A(net8008),
    .B(_09540_),
    .Y(_02269_));
 sky130_fd_sc_hd__xor2_1 _18034_ (.A(_02268_),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__or2b_1 _18035_ (.A(_02200_),
    .B_N(_02214_),
    .X(_02271_));
 sky130_fd_sc_hd__o21a_1 _18036_ (.A1(_02212_),
    .A2(_02213_),
    .B1(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__nor2_1 _18037_ (.A(_08366_),
    .B(_10289_),
    .Y(_02273_));
 sky130_fd_sc_hd__xnor2_1 _18038_ (.A(_02272_),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _18039_ (.A(_09181_),
    .B(_09060_),
    .Y(_02275_));
 sky130_fd_sc_hd__a21bo_1 _18040_ (.A1(_02201_),
    .A2(_02211_),
    .B1_N(_02209_),
    .X(_02276_));
 sky130_fd_sc_hd__xor2_1 _18041_ (.A(_02275_),
    .B(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__xnor2_1 _18042_ (.A(_02274_),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__o31a_1 _18043_ (.A1(_01784_),
    .A2(_09540_),
    .A3(_02166_),
    .B1(_02170_),
    .X(_02279_));
 sky130_fd_sc_hd__nand2_1 _18044_ (.A(_02204_),
    .B(_02205_),
    .Y(_02280_));
 sky130_fd_sc_hd__o31a_1 _18045_ (.A1(_01760_),
    .A2(_09114_),
    .A3(_02206_),
    .B1(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__or2_1 _18046_ (.A(_09040_),
    .B(_09114_),
    .X(_02282_));
 sky130_fd_sc_hd__xnor2_1 _18047_ (.A(_02281_),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__o21bai_2 _18048_ (.A1(_02164_),
    .A2(_02182_),
    .B1_N(_02181_),
    .Y(_02284_));
 sky130_fd_sc_hd__nor2_1 _18049_ (.A(_10316_),
    .B(_09345_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _18050_ (.A(_01760_),
    .B(net4908),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _18051_ (.A(_02285_),
    .B(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__xnor2_1 _18052_ (.A(_02284_),
    .B(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__o21a_1 _18053_ (.A1(_02192_),
    .A2(_02195_),
    .B1(_02193_),
    .X(_02289_));
 sky130_fd_sc_hd__nor2_1 _18054_ (.A(_08472_),
    .B(_09612_),
    .Y(_02290_));
 sky130_fd_sc_hd__xnor2_1 _18055_ (.A(_02289_),
    .B(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__xnor2_1 _18056_ (.A(_02288_),
    .B(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__xnor2_1 _18057_ (.A(_02283_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__xnor2_1 _18058_ (.A(_02279_),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__nor2_1 _18059_ (.A(_08612_),
    .B(_09410_),
    .Y(_02295_));
 sky130_fd_sc_hd__xnor2_1 _18060_ (.A(_02294_),
    .B(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__xnor2_1 _18061_ (.A(_02278_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _18062_ (.A(_01794_),
    .B(_01693_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _18063_ (.A(_01784_),
    .B(_09666_),
    .Y(_02299_));
 sky130_fd_sc_hd__nor2_1 _18064_ (.A(_10062_),
    .B(_09974_),
    .Y(_02300_));
 sky130_fd_sc_hd__xnor2_1 _18065_ (.A(_02299_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__xnor2_1 _18066_ (.A(_02298_),
    .B(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hd__xnor2_1 _18067_ (.A(_02297_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__xnor2_1 _18068_ (.A(_02270_),
    .B(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__xnor2_1 _18069_ (.A(_02266_),
    .B(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__xnor2_1 _18070_ (.A(_02225_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__xor2_1 _18071_ (.A(_02264_),
    .B(_02306_),
    .X(_02307_));
 sky130_fd_sc_hd__xnor2_1 _18072_ (.A(_02259_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__nand2_1 _18073_ (.A(_02258_),
    .B(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__or2_1 _18074_ (.A(_02258_),
    .B(_02308_),
    .X(_02310_));
 sky130_fd_sc_hd__and2_1 _18075_ (.A(_02309_),
    .B(_02310_),
    .X(_02311_));
 sky130_fd_sc_hd__a311oi_1 _18076_ (.A1(_02150_),
    .A2(_02153_),
    .A3(_02236_),
    .B1(_02253_),
    .C1(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__a311o_1 _18077_ (.A1(_02254_),
    .A2(_02309_),
    .A3(_02310_),
    .B1(_02312_),
    .C1(net90),
    .X(_02313_));
 sky130_fd_sc_hd__o21ai_1 _18078_ (.A1(_02250_),
    .A2(_02251_),
    .B1(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__mux2_4 _18079_ (.A0(_02314_),
    .A1(net4742),
    .S(_10260_),
    .X(_02315_));
 sky130_fd_sc_hd__clkbuf_1 _18080_ (.A(_02315_),
    .X(_00549_));
 sky130_fd_sc_hd__nand2_1 _18081_ (.A(net3749),
    .B(net4381),
    .Y(_02316_));
 sky130_fd_sc_hd__or2_1 _18082_ (.A(net3749),
    .B(net4381),
    .X(_02317_));
 sky130_fd_sc_hd__a31o_1 _18083_ (.A1(_09788_),
    .A2(net3700),
    .A3(_02317_),
    .B1(_09793_),
    .X(_02318_));
 sky130_fd_sc_hd__o211ai_1 _18084_ (.A1(net4646),
    .A2(_09413_),
    .B1(_06239_),
    .C1(net4781),
    .Y(_02319_));
 sky130_fd_sc_hd__buf_4 _18085_ (.A(net4782),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _18086_ (.A0(_02318_),
    .A1(net3749),
    .S(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__clkbuf_1 _18087_ (.A(_02321_),
    .X(_00550_));
 sky130_fd_sc_hd__or2_1 _18088_ (.A(net4518),
    .B(net4351),
    .X(_02322_));
 sky130_fd_sc_hd__nand2_1 _18089_ (.A(net4518),
    .B(net4351),
    .Y(_02323_));
 sky130_fd_sc_hd__nand2_1 _18090_ (.A(_02322_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_1 _18091_ (.A(net3700),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__o21ai_1 _18092_ (.A1(_06058_),
    .A2(net3701),
    .B1(_09801_),
    .Y(_02326_));
 sky130_fd_sc_hd__mux2_1 _18093_ (.A0(_02326_),
    .A1(net4518),
    .S(_02320_),
    .X(_02327_));
 sky130_fd_sc_hd__clkbuf_1 _18094_ (.A(_02327_),
    .X(_00551_));
 sky130_fd_sc_hd__o21a_1 _18095_ (.A1(net3700),
    .A2(_02324_),
    .B1(_02323_),
    .X(_02328_));
 sky130_fd_sc_hd__nor2_1 _18096_ (.A(net3932),
    .B(net4399),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _18097_ (.A(net3932),
    .B(net4399),
    .Y(_02330_));
 sky130_fd_sc_hd__or2b_1 _18098_ (.A(_02329_),
    .B_N(net3730),
    .X(_02331_));
 sky130_fd_sc_hd__xnor2_1 _18099_ (.A(_02328_),
    .B(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__o21ai_1 _18100_ (.A1(_06058_),
    .A2(_02332_),
    .B1(_09810_),
    .Y(_02333_));
 sky130_fd_sc_hd__mux2_1 _18101_ (.A0(_02333_),
    .A1(net3932),
    .S(_02320_),
    .X(_02334_));
 sky130_fd_sc_hd__clkbuf_1 _18102_ (.A(_02334_),
    .X(_00552_));
 sky130_fd_sc_hd__o21a_1 _18103_ (.A1(_02328_),
    .A2(_02329_),
    .B1(net3730),
    .X(_02335_));
 sky130_fd_sc_hd__nor2_1 _18104_ (.A(net3787),
    .B(net4539),
    .Y(_02336_));
 sky130_fd_sc_hd__nand2_1 _18105_ (.A(net3787),
    .B(net4539),
    .Y(_02337_));
 sky130_fd_sc_hd__or2b_1 _18106_ (.A(_02336_),
    .B_N(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__nor2_1 _18107_ (.A(net3731),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__a21o_1 _18108_ (.A1(net3731),
    .A2(_02338_),
    .B1(_09845_),
    .X(_02340_));
 sky130_fd_sc_hd__o21ai_1 _18109_ (.A1(_02339_),
    .A2(_02340_),
    .B1(_09820_),
    .Y(_02341_));
 sky130_fd_sc_hd__mux2_1 _18110_ (.A0(_02341_),
    .A1(net3787),
    .S(_02320_),
    .X(_02342_));
 sky130_fd_sc_hd__clkbuf_1 _18111_ (.A(_02342_),
    .X(_00553_));
 sky130_fd_sc_hd__or2_1 _18112_ (.A(net4565),
    .B(net4403),
    .X(_02343_));
 sky130_fd_sc_hd__nand2_1 _18113_ (.A(net4565),
    .B(net4403),
    .Y(_02344_));
 sky130_fd_sc_hd__o21ai_1 _18114_ (.A1(net3731),
    .A2(_02336_),
    .B1(_02337_),
    .Y(_02345_));
 sky130_fd_sc_hd__a21oi_1 _18115_ (.A1(_02343_),
    .A2(_02344_),
    .B1(net3732),
    .Y(_02346_));
 sky130_fd_sc_hd__a31o_1 _18116_ (.A1(net3732),
    .A2(_02343_),
    .A3(_02344_),
    .B1(_06057_),
    .X(_02347_));
 sky130_fd_sc_hd__o21ai_1 _18117_ (.A1(_02346_),
    .A2(net3733),
    .B1(_09829_),
    .Y(_02348_));
 sky130_fd_sc_hd__mux2_1 _18118_ (.A0(_02348_),
    .A1(net4565),
    .S(_02320_),
    .X(_02349_));
 sky130_fd_sc_hd__clkbuf_1 _18119_ (.A(_02349_),
    .X(_00554_));
 sky130_fd_sc_hd__a21boi_1 _18120_ (.A1(net3732),
    .A2(_02343_),
    .B1_N(_02344_),
    .Y(_02350_));
 sky130_fd_sc_hd__nor2_1 _18121_ (.A(net3847),
    .B(net4415),
    .Y(_02351_));
 sky130_fd_sc_hd__nand2_1 _18122_ (.A(net3847),
    .B(net4415),
    .Y(_02352_));
 sky130_fd_sc_hd__or2b_1 _18123_ (.A(_02351_),
    .B_N(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__xnor2_1 _18124_ (.A(_02350_),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__o21ai_1 _18125_ (.A1(_09809_),
    .A2(_02354_),
    .B1(_09837_),
    .Y(_02355_));
 sky130_fd_sc_hd__mux2_1 _18126_ (.A0(_02355_),
    .A1(net3847),
    .S(_02320_),
    .X(_02356_));
 sky130_fd_sc_hd__clkbuf_1 _18127_ (.A(_02356_),
    .X(_00555_));
 sky130_fd_sc_hd__o21a_1 _18128_ (.A1(_02350_),
    .A2(_02351_),
    .B1(_02352_),
    .X(_02357_));
 sky130_fd_sc_hd__nor2_1 _18129_ (.A(net3757),
    .B(net4379),
    .Y(_02358_));
 sky130_fd_sc_hd__nand2_1 _18130_ (.A(net3757),
    .B(net4379),
    .Y(_02359_));
 sky130_fd_sc_hd__or2b_1 _18131_ (.A(_02358_),
    .B_N(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__nor2_1 _18132_ (.A(net8039),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__a21o_1 _18133_ (.A1(net8039),
    .A2(_02360_),
    .B1(_09845_),
    .X(_02362_));
 sky130_fd_sc_hd__o21ai_1 _18134_ (.A1(_02361_),
    .A2(_02362_),
    .B1(_09847_),
    .Y(_02363_));
 sky130_fd_sc_hd__mux2_1 _18135_ (.A0(_02363_),
    .A1(net3757),
    .S(_02320_),
    .X(_02364_));
 sky130_fd_sc_hd__clkbuf_1 _18136_ (.A(_02364_),
    .X(_00556_));
 sky130_fd_sc_hd__o21a_1 _18137_ (.A1(net8039),
    .A2(_02358_),
    .B1(_02359_),
    .X(_02365_));
 sky130_fd_sc_hd__nor2_1 _18138_ (.A(net3768),
    .B(net4392),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _18139_ (.A(net3768),
    .B(net4392),
    .Y(_02367_));
 sky130_fd_sc_hd__or2b_1 _18140_ (.A(_02366_),
    .B_N(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__xnor2_1 _18141_ (.A(_02365_),
    .B(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__o21ai_1 _18142_ (.A1(_09809_),
    .A2(_02369_),
    .B1(_09855_),
    .Y(_02370_));
 sky130_fd_sc_hd__mux2_1 _18143_ (.A0(_02370_),
    .A1(net3768),
    .S(_02320_),
    .X(_02371_));
 sky130_fd_sc_hd__clkbuf_1 _18144_ (.A(_02371_),
    .X(_00557_));
 sky130_fd_sc_hd__o21a_1 _18145_ (.A1(_02365_),
    .A2(_02366_),
    .B1(_02367_),
    .X(_02372_));
 sky130_fd_sc_hd__nor2_1 _18146_ (.A(net3785),
    .B(net4390),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_1 _18147_ (.A(net3785),
    .B(net4390),
    .Y(_02374_));
 sky130_fd_sc_hd__or2b_1 _18148_ (.A(_02373_),
    .B_N(_02374_),
    .X(_02375_));
 sky130_fd_sc_hd__nor2_1 _18149_ (.A(_02372_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _18150_ (.A1(_02372_),
    .A2(_02375_),
    .B1(_09845_),
    .X(_02377_));
 sky130_fd_sc_hd__o21ai_1 _18151_ (.A1(_02376_),
    .A2(_02377_),
    .B1(_09864_),
    .Y(_02378_));
 sky130_fd_sc_hd__mux2_1 _18152_ (.A0(_02378_),
    .A1(net3785),
    .S(_02320_),
    .X(_02379_));
 sky130_fd_sc_hd__clkbuf_1 _18153_ (.A(_02379_),
    .X(_00558_));
 sky130_fd_sc_hd__or2_1 _18154_ (.A(net4567),
    .B(net4461),
    .X(_02380_));
 sky130_fd_sc_hd__nand2_1 _18155_ (.A(net4567),
    .B(net4461),
    .Y(_02381_));
 sky130_fd_sc_hd__o21ai_2 _18156_ (.A1(_02372_),
    .A2(_02373_),
    .B1(_02374_),
    .Y(_02382_));
 sky130_fd_sc_hd__a21oi_1 _18157_ (.A1(_02380_),
    .A2(_02381_),
    .B1(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__a31o_1 _18158_ (.A1(_02382_),
    .A2(_02380_),
    .A3(_02381_),
    .B1(_06057_),
    .X(_02384_));
 sky130_fd_sc_hd__o21ai_1 _18159_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_09872_),
    .Y(_02385_));
 sky130_fd_sc_hd__mux2_1 _18160_ (.A0(_02385_),
    .A1(net4567),
    .S(_02320_),
    .X(_02386_));
 sky130_fd_sc_hd__clkbuf_1 _18161_ (.A(_02386_),
    .X(_00559_));
 sky130_fd_sc_hd__nand2_1 _18162_ (.A(_02382_),
    .B(_02380_),
    .Y(_02387_));
 sky130_fd_sc_hd__and2_1 _18163_ (.A(net3790),
    .B(net3777),
    .X(_02388_));
 sky130_fd_sc_hd__nor2_1 _18164_ (.A(net3790),
    .B(net3777),
    .Y(_02389_));
 sky130_fd_sc_hd__a211oi_2 _18165_ (.A1(_02381_),
    .A2(_02387_),
    .B1(net3666),
    .C1(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__o211a_1 _18166_ (.A1(_02389_),
    .A2(net3666),
    .B1(_02387_),
    .C1(_02381_),
    .X(_02391_));
 sky130_fd_sc_hd__o31ai_1 _18167_ (.A1(_09809_),
    .A2(_02390_),
    .A3(_02391_),
    .B1(_09880_),
    .Y(_02392_));
 sky130_fd_sc_hd__buf_4 _18168_ (.A(net4782),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _18169_ (.A0(_02392_),
    .A1(net3790),
    .S(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__clkbuf_1 _18170_ (.A(_02394_),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _18171_ (.A(net4526),
    .B(net4496),
    .X(_02395_));
 sky130_fd_sc_hd__nand2_1 _18172_ (.A(net4526),
    .B(net4496),
    .Y(_02396_));
 sky130_fd_sc_hd__a211o_1 _18173_ (.A1(_02395_),
    .A2(_02396_),
    .B1(net3666),
    .C1(_02390_),
    .X(_02397_));
 sky130_fd_sc_hd__o211ai_2 _18174_ (.A1(net3666),
    .A2(_02390_),
    .B1(_02395_),
    .C1(_02396_),
    .Y(_02398_));
 sky130_fd_sc_hd__a31o_1 _18175_ (.A1(_02245_),
    .A2(net3667),
    .A3(_02398_),
    .B1(_10010_),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _18176_ (.A0(_02399_),
    .A1(net4526),
    .S(_02393_),
    .X(_02400_));
 sky130_fd_sc_hd__clkbuf_1 _18177_ (.A(_02400_),
    .X(_00561_));
 sky130_fd_sc_hd__and2_1 _18178_ (.A(net3751),
    .B(net4435),
    .X(_02401_));
 sky130_fd_sc_hd__nor2_1 _18179_ (.A(net3751),
    .B(net4435),
    .Y(_02402_));
 sky130_fd_sc_hd__a211o_1 _18180_ (.A1(_02396_),
    .A2(_02398_),
    .B1(_02401_),
    .C1(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__o211ai_1 _18181_ (.A1(_02401_),
    .A2(_02402_),
    .B1(_02396_),
    .C1(_02398_),
    .Y(_02404_));
 sky130_fd_sc_hd__a31o_1 _18182_ (.A1(_02245_),
    .A2(_02403_),
    .A3(_02404_),
    .B1(_10133_),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _18183_ (.A0(_02405_),
    .A1(net3751),
    .S(_02393_),
    .X(_02406_));
 sky130_fd_sc_hd__clkbuf_1 _18184_ (.A(_02406_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_2 _18185_ (.A(net3766),
    .B(net4481),
    .Y(_02407_));
 sky130_fd_sc_hd__or2_1 _18186_ (.A(net3766),
    .B(net4481),
    .X(_02408_));
 sky130_fd_sc_hd__inv_2 _18187_ (.A(_02403_),
    .Y(_02409_));
 sky130_fd_sc_hd__a211o_1 _18188_ (.A1(_02407_),
    .A2(_02408_),
    .B1(_02401_),
    .C1(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__o211ai_2 _18189_ (.A1(_02401_),
    .A2(_02409_),
    .B1(_02407_),
    .C1(_02408_),
    .Y(_02411_));
 sky130_fd_sc_hd__a31o_1 _18190_ (.A1(_02245_),
    .A2(_02410_),
    .A3(_02411_),
    .B1(_10258_),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _18191_ (.A0(_02412_),
    .A1(net3766),
    .S(_02393_),
    .X(_02413_));
 sky130_fd_sc_hd__clkbuf_1 _18192_ (.A(_02413_),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _18193_ (.A(net3811),
    .B(net4430),
    .X(_02414_));
 sky130_fd_sc_hd__nor2_1 _18194_ (.A(net3811),
    .B(net4430),
    .Y(_02415_));
 sky130_fd_sc_hd__a211oi_2 _18195_ (.A1(_02407_),
    .A2(_02411_),
    .B1(_02414_),
    .C1(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__o211a_1 _18196_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_02407_),
    .C1(_02411_),
    .X(_02417_));
 sky130_fd_sc_hd__o31ai_1 _18197_ (.A1(_09809_),
    .A2(_02416_),
    .A3(_02417_),
    .B1(_10380_),
    .Y(_02418_));
 sky130_fd_sc_hd__mux2_1 _18198_ (.A0(_02418_),
    .A1(net3811),
    .S(_02393_),
    .X(_02419_));
 sky130_fd_sc_hd__clkbuf_1 _18199_ (.A(_02419_),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _18200_ (.A(net3669),
    .B(net4459),
    .Y(_02420_));
 sky130_fd_sc_hd__or2_1 _18201_ (.A(net3669),
    .B(net4459),
    .X(_02421_));
 sky130_fd_sc_hd__nand2_1 _18202_ (.A(_02420_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__nor2_1 _18203_ (.A(_02414_),
    .B(_02416_),
    .Y(_02423_));
 sky130_fd_sc_hd__xnor2_1 _18204_ (.A(_02422_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__o21ai_1 _18205_ (.A1(_09809_),
    .A2(_02424_),
    .B1(_01729_),
    .Y(_02425_));
 sky130_fd_sc_hd__mux2_1 _18206_ (.A0(_02425_),
    .A1(net3669),
    .S(_02393_),
    .X(_02426_));
 sky130_fd_sc_hd__clkbuf_1 _18207_ (.A(_02426_),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _18208_ (.A(net3803),
    .B(net4440),
    .Y(_02427_));
 sky130_fd_sc_hd__nand2_1 _18209_ (.A(net3803),
    .B(net4440),
    .Y(_02428_));
 sky130_fd_sc_hd__or2b_1 _18210_ (.A(_02427_),
    .B_N(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__o21a_1 _18211_ (.A1(_02422_),
    .A2(_02423_),
    .B1(_02420_),
    .X(_02430_));
 sky130_fd_sc_hd__xnor2_1 _18212_ (.A(_02429_),
    .B(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__o21ai_1 _18213_ (.A1(_09809_),
    .A2(_02431_),
    .B1(_01844_),
    .Y(_02432_));
 sky130_fd_sc_hd__mux2_1 _18214_ (.A0(_02432_),
    .A1(net3803),
    .S(_02393_),
    .X(_02433_));
 sky130_fd_sc_hd__clkbuf_1 _18215_ (.A(_02433_),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_1 _18216_ (.A(net4575),
    .B(net4428),
    .Y(_02434_));
 sky130_fd_sc_hd__nand2_1 _18217_ (.A(net4575),
    .B(net4428),
    .Y(_02435_));
 sky130_fd_sc_hd__or2b_1 _18218_ (.A(_02434_),
    .B_N(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__o21a_1 _18219_ (.A1(_02427_),
    .A2(_02430_),
    .B1(_02428_),
    .X(_02437_));
 sky130_fd_sc_hd__nor2_1 _18220_ (.A(_02436_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__a21o_1 _18221_ (.A1(_02436_),
    .A2(_02437_),
    .B1(_09845_),
    .X(_02439_));
 sky130_fd_sc_hd__o21ai_1 _18222_ (.A1(_02438_),
    .A2(_02439_),
    .B1(_01953_),
    .Y(_02440_));
 sky130_fd_sc_hd__mux2_1 _18223_ (.A0(_02440_),
    .A1(net4575),
    .S(_02393_),
    .X(_02441_));
 sky130_fd_sc_hd__clkbuf_1 _18224_ (.A(_02441_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _18225_ (.A(net3820),
    .B(net4537),
    .Y(_02442_));
 sky130_fd_sc_hd__nand2_1 _18226_ (.A(net3820),
    .B(net4537),
    .Y(_02443_));
 sky130_fd_sc_hd__or2b_1 _18227_ (.A(_02442_),
    .B_N(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__o21a_1 _18228_ (.A1(_02434_),
    .A2(_02437_),
    .B1(_02435_),
    .X(_02445_));
 sky130_fd_sc_hd__nor2_1 _18229_ (.A(_02444_),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__a21o_1 _18230_ (.A1(_02444_),
    .A2(_02445_),
    .B1(_09845_),
    .X(_02447_));
 sky130_fd_sc_hd__o21ai_1 _18231_ (.A1(_02446_),
    .A2(_02447_),
    .B1(_02052_),
    .Y(_02448_));
 sky130_fd_sc_hd__mux2_1 _18232_ (.A0(_02448_),
    .A1(net3820),
    .S(_02393_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_1 _18233_ (.A(_02449_),
    .X(_00568_));
 sky130_fd_sc_hd__or2_1 _18234_ (.A(net3835),
    .B(net4524),
    .X(_02450_));
 sky130_fd_sc_hd__nand2_1 _18235_ (.A(net3835),
    .B(net4524),
    .Y(_02451_));
 sky130_fd_sc_hd__nand2_1 _18236_ (.A(_02450_),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__o21ai_1 _18237_ (.A1(_02442_),
    .A2(_02445_),
    .B1(_02443_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_1 _18238_ (.A(_02452_),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__a21o_1 _18239_ (.A1(_09788_),
    .A2(_02454_),
    .B1(_02155_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _18240_ (.A0(_02455_),
    .A1(net3835),
    .S(_02393_),
    .X(_02456_));
 sky130_fd_sc_hd__clkbuf_1 _18241_ (.A(_02456_),
    .X(_00569_));
 sky130_fd_sc_hd__nand2_1 _18242_ (.A(net3926),
    .B(net4608),
    .Y(_02457_));
 sky130_fd_sc_hd__or2_1 _18243_ (.A(net3926),
    .B(net4608),
    .X(_02458_));
 sky130_fd_sc_hd__nand2_1 _18244_ (.A(_02457_),
    .B(net3588),
    .Y(_02459_));
 sky130_fd_sc_hd__a21bo_1 _18245_ (.A1(_02450_),
    .A2(_02453_),
    .B1_N(_02451_),
    .X(_02460_));
 sky130_fd_sc_hd__xnor2_1 _18246_ (.A(_02459_),
    .B(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__a22o_1 _18247_ (.A1(_02238_),
    .A2(_02239_),
    .B1(_02461_),
    .B2(_02245_),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_4 _18248_ (.A0(_02462_),
    .A1(net3926),
    .S(net4782),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_1 _18249_ (.A(_02463_),
    .X(_00570_));
 sky130_fd_sc_hd__a21bo_1 _18250_ (.A1(net3588),
    .A2(_02460_),
    .B1_N(_02457_),
    .X(_02464_));
 sky130_fd_sc_hd__xnor2_1 _18251_ (.A(_06162_),
    .B(net3589),
    .Y(_02465_));
 sky130_fd_sc_hd__nor2_1 _18252_ (.A(net4413),
    .B(net3590),
    .Y(_02466_));
 sky130_fd_sc_hd__a21o_1 _18253_ (.A1(net4413),
    .A2(net3590),
    .B1(_06057_),
    .X(_02467_));
 sky130_fd_sc_hd__o21ai_1 _18254_ (.A1(net3591),
    .A2(_02467_),
    .B1(_02313_),
    .Y(_02468_));
 sky130_fd_sc_hd__mux2_4 _18255_ (.A0(_02468_),
    .A1(net4498),
    .S(net4782),
    .X(_02469_));
 sky130_fd_sc_hd__clkbuf_1 _18256_ (.A(_02469_),
    .X(_00571_));
 sky130_fd_sc_hd__clkbuf_1 _18257_ (.A(net3897),
    .X(_02470_));
 sky130_fd_sc_hd__inv_2 _18258_ (.A(net3770),
    .Y(_02471_));
 sky130_fd_sc_hd__clkbuf_4 _18259_ (.A(net4832),
    .X(_02472_));
 sky130_fd_sc_hd__nor2_1 _18260_ (.A(net1879),
    .B(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__and3b_1 _18261_ (.A_N(net3940),
    .B(net4814),
    .C(net3906),
    .X(_02474_));
 sky130_fd_sc_hd__nand2_2 _18262_ (.A(net1880),
    .B(net4815),
    .Y(_02475_));
 sky130_fd_sc_hd__nor2_4 _18263_ (.A(_04458_),
    .B(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__buf_4 _18264_ (.A(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _18265_ (.A0(net6355),
    .A1(net1622),
    .S(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__clkbuf_1 _18266_ (.A(net1287),
    .X(_00572_));
 sky130_fd_sc_hd__clkbuf_1 _18267_ (.A(net4028),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _18268_ (.A0(net6393),
    .A1(net1396),
    .S(_02477_),
    .X(_02480_));
 sky130_fd_sc_hd__clkbuf_1 _18269_ (.A(net1397),
    .X(_00573_));
 sky130_fd_sc_hd__buf_1 _18270_ (.A(net6476),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _18271_ (.A0(net6335),
    .A1(net1493),
    .S(_02477_),
    .X(_02482_));
 sky130_fd_sc_hd__clkbuf_1 _18272_ (.A(net6337),
    .X(_00574_));
 sky130_fd_sc_hd__clkbuf_1 _18273_ (.A(net4074),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _18274_ (.A0(net6291),
    .A1(net1426),
    .S(_02477_),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_1 _18275_ (.A(net1282),
    .X(_00575_));
 sky130_fd_sc_hd__buf_1 _18276_ (.A(net4038),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _18277_ (.A0(net6299),
    .A1(net4016),
    .S(_02477_),
    .X(_02486_));
 sky130_fd_sc_hd__clkbuf_1 _18278_ (.A(net1242),
    .X(_00576_));
 sky130_fd_sc_hd__clkbuf_1 _18279_ (.A(net2204),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _18280_ (.A0(net6390),
    .A1(net2205),
    .S(_02477_),
    .X(_02488_));
 sky130_fd_sc_hd__clkbuf_1 _18281_ (.A(net1420),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _18282_ (.A0(net6492),
    .A1(net3863),
    .S(_02477_),
    .X(_02489_));
 sky130_fd_sc_hd__clkbuf_1 _18283_ (.A(net1539),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _18284_ (.A0(net6454),
    .A1(net3816),
    .S(_02477_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _18285_ (.A(net1632),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _18286_ (.A0(net6405),
    .A1(net3402),
    .S(_02477_),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_1 _18287_ (.A(net1509),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _18288_ (.A0(net6363),
    .A1(net2953),
    .S(_02477_),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_1 _18289_ (.A(net6365),
    .X(_00581_));
 sky130_fd_sc_hd__buf_4 _18290_ (.A(_02476_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _18291_ (.A0(net6307),
    .A1(net3838),
    .S(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__clkbuf_1 _18292_ (.A(net1436),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _18293_ (.A0(net6558),
    .A1(net3745),
    .S(_02493_),
    .X(_02495_));
 sky130_fd_sc_hd__clkbuf_1 _18294_ (.A(net1860),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _18295_ (.A0(net6407),
    .A1(net3596),
    .S(_02493_),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_1 _18296_ (.A(net1457),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _18297_ (.A0(net6585),
    .A1(net3562),
    .S(_02493_),
    .X(_02497_));
 sky130_fd_sc_hd__clkbuf_1 _18298_ (.A(net1678),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _18299_ (.A0(net6339),
    .A1(net3738),
    .S(_02493_),
    .X(_02498_));
 sky130_fd_sc_hd__clkbuf_1 _18300_ (.A(net1381),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _18301_ (.A0(net6380),
    .A1(net3592),
    .S(_02493_),
    .X(_02499_));
 sky130_fd_sc_hd__clkbuf_1 _18302_ (.A(net6382),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _18303_ (.A0(net6384),
    .A1(net3556),
    .S(_02493_),
    .X(_02500_));
 sky130_fd_sc_hd__clkbuf_1 _18304_ (.A(net6386),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _18305_ (.A0(net6603),
    .A1(net3674),
    .S(_02493_),
    .X(_02501_));
 sky130_fd_sc_hd__clkbuf_1 _18306_ (.A(net6605),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _18307_ (.A0(net6528),
    .A1(net3866),
    .S(_02493_),
    .X(_02502_));
 sky130_fd_sc_hd__clkbuf_1 _18308_ (.A(net6530),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _18309_ (.A0(net6426),
    .A1(net1447),
    .S(_02493_),
    .X(_02503_));
 sky130_fd_sc_hd__clkbuf_1 _18310_ (.A(net6428),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _18311_ (.A0(net6191),
    .A1(net3478),
    .S(_02476_),
    .X(_02504_));
 sky130_fd_sc_hd__clkbuf_1 _18312_ (.A(net6193),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _18313_ (.A0(net6148),
    .A1(net3481),
    .S(_02476_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _18314_ (.A(net6150),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _18315_ (.A0(net6160),
    .A1(net3583),
    .S(_02476_),
    .X(_02506_));
 sky130_fd_sc_hd__clkbuf_1 _18316_ (.A(net6162),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _18317_ (.A0(net6331),
    .A1(net3631),
    .S(_02476_),
    .X(_02507_));
 sky130_fd_sc_hd__clkbuf_1 _18318_ (.A(net6333),
    .X(_00595_));
 sky130_fd_sc_hd__clkbuf_4 _18319_ (.A(_09735_),
    .X(_02508_));
 sky130_fd_sc_hd__nor2_1 _18320_ (.A(net4501),
    .B(net4852),
    .Y(_02509_));
 sky130_fd_sc_hd__nor2_1 _18321_ (.A(net4733),
    .B(net4887),
    .Y(_02510_));
 sky130_fd_sc_hd__nand2_1 _18322_ (.A(_05155_),
    .B(net693),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2_1 _18323_ (.A(net3565),
    .B(net5033),
    .Y(_02512_));
 sky130_fd_sc_hd__or2_1 _18324_ (.A(net4713),
    .B(net693),
    .X(_02513_));
 sky130_fd_sc_hd__nand3b_1 _18325_ (.A_N(_02512_),
    .B(net4714),
    .C(_02511_),
    .Y(_02514_));
 sky130_fd_sc_hd__and2_1 _18326_ (.A(_02511_),
    .B(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__nand2_1 _18327_ (.A(net4733),
    .B(net4887),
    .Y(_02516_));
 sky130_fd_sc_hd__o21a_1 _18328_ (.A1(_02510_),
    .A2(_02515_),
    .B1(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__nand2_1 _18329_ (.A(net4501),
    .B(net4852),
    .Y(_02518_));
 sky130_fd_sc_hd__o21a_1 _18330_ (.A1(_02509_),
    .A2(_02517_),
    .B1(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__nor2_1 _18331_ (.A(net3660),
    .B(net4883),
    .Y(_02520_));
 sky130_fd_sc_hd__nand2_1 _18332_ (.A(net3661),
    .B(net4883),
    .Y(_02521_));
 sky130_fd_sc_hd__or2b_1 _18333_ (.A(_02520_),
    .B_N(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__xor2_1 _18334_ (.A(_02519_),
    .B(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__inv_2 _18335_ (.A(net3565),
    .Y(_02524_));
 sky130_fd_sc_hd__nor2_1 _18336_ (.A(_02524_),
    .B(_08038_),
    .Y(_02525_));
 sky130_fd_sc_hd__a221o_1 _18337_ (.A1(net4883),
    .A2(_02508_),
    .B1(_09739_),
    .B2(net8255),
    .C1(_02525_),
    .X(_00596_));
 sky130_fd_sc_hd__buf_4 _18338_ (.A(_04478_),
    .X(_02526_));
 sky130_fd_sc_hd__nand2_1 _18339_ (.A(_05155_),
    .B(net3565),
    .Y(_02527_));
 sky130_fd_sc_hd__or2_1 _18340_ (.A(_05155_),
    .B(net3565),
    .X(_02528_));
 sky130_fd_sc_hd__o21a_1 _18341_ (.A1(_02519_),
    .A2(_02520_),
    .B1(_02521_),
    .X(_02529_));
 sky130_fd_sc_hd__nor2_1 _18342_ (.A(net3509),
    .B(net5961),
    .Y(_02530_));
 sky130_fd_sc_hd__nand2_1 _18343_ (.A(net3509),
    .B(net5961),
    .Y(_02531_));
 sky130_fd_sc_hd__or2b_1 _18344_ (.A(_02530_),
    .B_N(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__or2_1 _18345_ (.A(_02529_),
    .B(_02532_),
    .X(_02533_));
 sky130_fd_sc_hd__a21oi_1 _18346_ (.A1(_02529_),
    .A2(_02532_),
    .B1(_04489_),
    .Y(_02534_));
 sky130_fd_sc_hd__a32o_1 _18347_ (.A1(_02526_),
    .A2(_02527_),
    .A3(_02528_),
    .B1(_02533_),
    .B2(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__nand2_1 _18348_ (.A(_04480_),
    .B(_09734_),
    .Y(_02536_));
 sky130_fd_sc_hd__buf_4 _18349_ (.A(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _18350_ (.A0(net5961),
    .A1(_02535_),
    .S(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_1 _18351_ (.A(net5963),
    .X(_00597_));
 sky130_fd_sc_hd__nand2_1 _18352_ (.A(net4733),
    .B(_02528_),
    .Y(_02539_));
 sky130_fd_sc_hd__or2_1 _18353_ (.A(net4733),
    .B(_02528_),
    .X(_02540_));
 sky130_fd_sc_hd__o21a_1 _18354_ (.A1(_02529_),
    .A2(_02530_),
    .B1(_02531_),
    .X(_02541_));
 sky130_fd_sc_hd__nor2_1 _18355_ (.A(net4698),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_1 _18356_ (.A(net4698),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02543_));
 sky130_fd_sc_hd__or2b_1 _18357_ (.A(_02542_),
    .B_N(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__or2_1 _18358_ (.A(_02541_),
    .B(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__a21oi_1 _18359_ (.A1(_02541_),
    .A2(_02544_),
    .B1(_04489_),
    .Y(_02546_));
 sky130_fd_sc_hd__a32o_1 _18360_ (.A1(_02526_),
    .A2(_02539_),
    .A3(_02540_),
    .B1(_02545_),
    .B2(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__mux2_1 _18361_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_02547_),
    .S(_02537_),
    .X(_02548_));
 sky130_fd_sc_hd__clkbuf_1 _18362_ (.A(net5823),
    .X(_00598_));
 sky130_fd_sc_hd__or4_1 _18363_ (.A(net4501),
    .B(net4733),
    .C(_05155_),
    .D(net3565),
    .X(_02549_));
 sky130_fd_sc_hd__a21oi_1 _18364_ (.A1(net4501),
    .A2(_02540_),
    .B1(_04480_),
    .Y(_02550_));
 sky130_fd_sc_hd__o21ai_2 _18365_ (.A1(_02541_),
    .A2(_02542_),
    .B1(_02543_),
    .Y(_02551_));
 sky130_fd_sc_hd__clkbuf_1 _18366_ (.A(net3493),
    .X(_02552_));
 sky130_fd_sc_hd__nor2_1 _18367_ (.A(net3494),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_02553_));
 sky130_fd_sc_hd__and2_1 _18368_ (.A(net3493),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02554_));
 sky130_fd_sc_hd__or2_1 _18369_ (.A(_02553_),
    .B(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__xnor2_1 _18370_ (.A(_02551_),
    .B(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__a22o_1 _18371_ (.A1(_02549_),
    .A2(_02550_),
    .B1(_02556_),
    .B2(_04481_),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _18372_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_02557_),
    .S(_02537_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_1 _18373_ (.A(net5832),
    .X(_00599_));
 sky130_fd_sc_hd__buf_4 _18374_ (.A(_09738_),
    .X(_02559_));
 sky130_fd_sc_hd__o21a_1 _18375_ (.A1(net3494),
    .A2(\rbzero.wall_tracer.rayAddendX[-2] ),
    .B1(_02551_),
    .X(_02560_));
 sky130_fd_sc_hd__nand2_1 _18376_ (.A(net4554),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_02561_));
 sky130_fd_sc_hd__or2_1 _18377_ (.A(net4554),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02562_));
 sky130_fd_sc_hd__o211a_1 _18378_ (.A1(_02554_),
    .A2(_02560_),
    .B1(net4784),
    .C1(net8047),
    .X(_02563_));
 sky130_fd_sc_hd__inv_2 _18379_ (.A(net8048),
    .Y(_02564_));
 sky130_fd_sc_hd__a211o_1 _18380_ (.A1(net8047),
    .A2(net4784),
    .B1(_02560_),
    .C1(_02554_),
    .X(_02565_));
 sky130_fd_sc_hd__o31a_1 _18381_ (.A1(net4501),
    .A2(net4733),
    .A3(_05155_),
    .B1(_02524_),
    .X(_02566_));
 sky130_fd_sc_hd__or2_1 _18382_ (.A(net3661),
    .B(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__nand2_1 _18383_ (.A(net3661),
    .B(_02566_),
    .Y(_02568_));
 sky130_fd_sc_hd__a32o_1 _18384_ (.A1(_04490_),
    .A2(_02567_),
    .A3(_02568_),
    .B1(_09736_),
    .B2(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02569_));
 sky130_fd_sc_hd__a31o_1 _18385_ (.A1(_02559_),
    .A2(net8049),
    .A3(net4785),
    .B1(net3514),
    .X(_00600_));
 sky130_fd_sc_hd__xor2_1 _18386_ (.A(net3509),
    .B(_05155_),
    .X(_02570_));
 sky130_fd_sc_hd__nand2_1 _18387_ (.A(net3661),
    .B(net3565),
    .Y(_02571_));
 sky130_fd_sc_hd__o21ai_1 _18388_ (.A1(net3661),
    .A2(_02549_),
    .B1(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__xnor2_1 _18389_ (.A(_02570_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__nand2_1 _18390_ (.A(net4784),
    .B(_02564_),
    .Y(_02574_));
 sky130_fd_sc_hd__or2_1 _18391_ (.A(net4603),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_1 _18392_ (.A(net4603),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_02576_));
 sky130_fd_sc_hd__nand2_1 _18393_ (.A(_02575_),
    .B(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__xnor2_1 _18394_ (.A(_02574_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__mux2_1 _18395_ (.A0(_02573_),
    .A1(_02578_),
    .S(_04480_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _18396_ (.A0(\rbzero.wall_tracer.rayAddendX[0] ),
    .A1(_02579_),
    .S(_02537_),
    .X(_02580_));
 sky130_fd_sc_hd__clkbuf_1 _18397_ (.A(net5884),
    .X(_00601_));
 sky130_fd_sc_hd__nand2_1 _18398_ (.A(net4724),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_02581_));
 sky130_fd_sc_hd__or2_1 _18399_ (.A(net4724),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02582_));
 sky130_fd_sc_hd__a21bo_1 _18400_ (.A1(_02574_),
    .A2(_02575_),
    .B1_N(_02576_),
    .X(_02583_));
 sky130_fd_sc_hd__a21o_1 _18401_ (.A1(net4725),
    .A2(net8074),
    .B1(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__and3_1 _18402_ (.A(net4725),
    .B(net8074),
    .C(_02583_),
    .X(_02585_));
 sky130_fd_sc_hd__inv_2 _18403_ (.A(net8075),
    .Y(_02586_));
 sky130_fd_sc_hd__nor2_1 _18404_ (.A(net4698),
    .B(net4733),
    .Y(_02587_));
 sky130_fd_sc_hd__and2_1 _18405_ (.A(net4698),
    .B(net4733),
    .X(_02588_));
 sky130_fd_sc_hd__nor4_2 _18406_ (.A(net3509),
    .B(_05155_),
    .C(_02587_),
    .D(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__o22a_1 _18407_ (.A1(net3509),
    .A2(_05155_),
    .B1(_02587_),
    .B2(_02588_),
    .X(_02590_));
 sky130_fd_sc_hd__or2_1 _18408_ (.A(_02589_),
    .B(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__o2bb2a_1 _18409_ (.A1_N(_02570_),
    .A2_N(_02571_),
    .B1(net3661),
    .B2(_02549_),
    .X(_02592_));
 sky130_fd_sc_hd__nor2_1 _18410_ (.A(_02591_),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__a21o_1 _18411_ (.A1(_02591_),
    .A2(_02592_),
    .B1(_04481_),
    .X(_02594_));
 sky130_fd_sc_hd__a2bb2o_1 _18412_ (.A1_N(_02593_),
    .A2_N(_02594_),
    .B1(\rbzero.wall_tracer.rayAddendX[1] ),
    .B2(_09736_),
    .X(_02595_));
 sky130_fd_sc_hd__a31o_1 _18413_ (.A1(_02559_),
    .A2(net4726),
    .A3(net8076),
    .B1(net3639),
    .X(_00602_));
 sky130_fd_sc_hd__xor2_1 _18414_ (.A(net4724),
    .B(net3604),
    .X(_02596_));
 sky130_fd_sc_hd__and2_1 _18415_ (.A(net4725),
    .B(_02586_),
    .X(_02597_));
 sky130_fd_sc_hd__xnor2_1 _18416_ (.A(_02596_),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__xor2_2 _18417_ (.A(net3494),
    .B(net4501),
    .X(_02599_));
 sky130_fd_sc_hd__or3_1 _18418_ (.A(_02589_),
    .B(_02593_),
    .C(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__o21ai_2 _18419_ (.A1(_02589_),
    .A2(_02593_),
    .B1(_02599_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand2_1 _18420_ (.A(_02600_),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__xnor2_1 _18421_ (.A(_02587_),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__mux2_1 _18422_ (.A0(_02598_),
    .A1(_02603_),
    .S(_02526_),
    .X(_02604_));
 sky130_fd_sc_hd__mux2_1 _18423_ (.A0(net3604),
    .A1(_02604_),
    .S(_02537_),
    .X(_02605_));
 sky130_fd_sc_hd__clkbuf_1 _18424_ (.A(net5972),
    .X(_00603_));
 sky130_fd_sc_hd__inv_2 _18425_ (.A(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02606_));
 sky130_fd_sc_hd__or2_1 _18426_ (.A(net4554),
    .B(net3661),
    .X(_02607_));
 sky130_fd_sc_hd__nand2_1 _18427_ (.A(net4554),
    .B(net3661),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_1 _18428_ (.A(_02607_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__or3_1 _18429_ (.A(net3494),
    .B(net4501),
    .C(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__o21ai_1 _18430_ (.A1(net3494),
    .A2(net4501),
    .B1(_02609_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand2_1 _18431_ (.A(_02610_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__o21ai_1 _18432_ (.A1(_02593_),
    .A2(_02599_),
    .B1(_02587_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21o_1 _18433_ (.A1(_02601_),
    .A2(_02613_),
    .B1(_02612_),
    .X(_02614_));
 sky130_fd_sc_hd__nand2_1 _18434_ (.A(_04490_),
    .B(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__a31o_1 _18435_ (.A1(_02601_),
    .A2(_02612_),
    .A3(_02613_),
    .B1(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__clkbuf_4 _18436_ (.A(net4724),
    .X(_02617_));
 sky130_fd_sc_hd__nand2_1 _18437_ (.A(_02617_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02618_));
 sky130_fd_sc_hd__or2_1 _18438_ (.A(net4724),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02619_));
 sky130_fd_sc_hd__o21a_1 _18439_ (.A1(net3604),
    .A2(\rbzero.wall_tracer.rayAddendX[1] ),
    .B1(net4724),
    .X(_02620_));
 sky130_fd_sc_hd__a21o_1 _18440_ (.A1(_02585_),
    .A2(_02596_),
    .B1(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__a21oi_1 _18441_ (.A1(net4791),
    .A2(_02619_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__and3_1 _18442_ (.A(net4791),
    .B(_02619_),
    .C(_02621_),
    .X(_02623_));
 sky130_fd_sc_hd__or3_1 _18443_ (.A(_09747_),
    .B(net4792),
    .C(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__o211ai_1 _18444_ (.A1(net8109),
    .A2(_02537_),
    .B1(_02616_),
    .C1(net4793),
    .Y(_00604_));
 sky130_fd_sc_hd__xor2_1 _18445_ (.A(_02617_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_02625_));
 sky130_fd_sc_hd__buf_2 _18446_ (.A(_02617_),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_4 _18447_ (.A(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__a21oi_1 _18448_ (.A1(_02627_),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02623_),
    .Y(_02628_));
 sky130_fd_sc_hd__xnor2_1 _18449_ (.A(_02625_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__nor2_1 _18450_ (.A(net4603),
    .B(net3509),
    .Y(_02630_));
 sky130_fd_sc_hd__and2_1 _18451_ (.A(net4603),
    .B(net3509),
    .X(_02631_));
 sky130_fd_sc_hd__or2_1 _18452_ (.A(_02630_),
    .B(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__nand3_1 _18453_ (.A(_02610_),
    .B(_02614_),
    .C(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__a21o_1 _18454_ (.A1(_02610_),
    .A2(_02614_),
    .B1(_02632_),
    .X(_02634_));
 sky130_fd_sc_hd__a21oi_1 _18455_ (.A1(_02633_),
    .A2(_02634_),
    .B1(_02607_),
    .Y(_02635_));
 sky130_fd_sc_hd__and3_1 _18456_ (.A(_02607_),
    .B(_02633_),
    .C(_02634_),
    .X(_02636_));
 sky130_fd_sc_hd__or2_1 _18457_ (.A(_02635_),
    .B(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _18458_ (.A0(_02629_),
    .A1(_02637_),
    .S(_02526_),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_1 _18459_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02638_),
    .S(_02537_),
    .X(_02639_));
 sky130_fd_sc_hd__clkbuf_1 _18460_ (.A(net5874),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _18461_ (.A(_02617_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02640_));
 sky130_fd_sc_hd__or2_1 _18462_ (.A(_02617_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_02641_));
 sky130_fd_sc_hd__and2_1 _18463_ (.A(net8084),
    .B(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__and2_1 _18464_ (.A(_02623_),
    .B(_02625_),
    .X(_02643_));
 sky130_fd_sc_hd__o21a_1 _18465_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02617_),
    .X(_02644_));
 sky130_fd_sc_hd__or3_1 _18466_ (.A(net8085),
    .B(_02643_),
    .C(net4820),
    .X(_02645_));
 sky130_fd_sc_hd__o21ai_2 _18467_ (.A1(_02643_),
    .A2(net4820),
    .B1(net8085),
    .Y(_02646_));
 sky130_fd_sc_hd__a21o_1 _18468_ (.A1(_02614_),
    .A2(_02632_),
    .B1(_02607_),
    .X(_02647_));
 sky130_fd_sc_hd__xor2_1 _18469_ (.A(_02617_),
    .B(net4698),
    .X(_02648_));
 sky130_fd_sc_hd__xnor2_1 _18470_ (.A(_02630_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__a21oi_1 _18471_ (.A1(_02634_),
    .A2(_02647_),
    .B1(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__a31o_1 _18472_ (.A1(_02634_),
    .A2(_02649_),
    .A3(_02647_),
    .B1(_04481_),
    .X(_02651_));
 sky130_fd_sc_hd__a2bb2o_1 _18473_ (.A1_N(_02650_),
    .A2_N(_02651_),
    .B1(\rbzero.wall_tracer.rayAddendX[5] ),
    .B2(_09735_),
    .X(_02652_));
 sky130_fd_sc_hd__a31o_1 _18474_ (.A1(_02559_),
    .A2(net4821),
    .A3(net8086),
    .B1(net3947),
    .X(_00606_));
 sky130_fd_sc_hd__xnor2_2 _18475_ (.A(_02617_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_02653_));
 sky130_fd_sc_hd__a21oi_1 _18476_ (.A1(_02640_),
    .A2(_02646_),
    .B1(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__a31o_1 _18477_ (.A1(_02640_),
    .A2(_02646_),
    .A3(_02653_),
    .B1(_04489_),
    .X(_02655_));
 sky130_fd_sc_hd__or2_1 _18478_ (.A(_02617_),
    .B(net3494),
    .X(_02656_));
 sky130_fd_sc_hd__nand2_1 _18479_ (.A(_02626_),
    .B(net3494),
    .Y(_02657_));
 sky130_fd_sc_hd__a2bb2o_1 _18480_ (.A1_N(_02626_),
    .A2_N(net4698),
    .B1(_02656_),
    .B2(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__or3b_1 _18481_ (.A(_02626_),
    .B(net4698),
    .C_N(net3494),
    .X(_02659_));
 sky130_fd_sc_hd__nand2_1 _18482_ (.A(_02658_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__a21o_1 _18483_ (.A1(_02630_),
    .A2(_02648_),
    .B1(_02650_),
    .X(_02661_));
 sky130_fd_sc_hd__xnor2_1 _18484_ (.A(_02660_),
    .B(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__a2bb2o_1 _18485_ (.A1_N(_02654_),
    .A2_N(_02655_),
    .B1(_02662_),
    .B2(_02526_),
    .X(_02663_));
 sky130_fd_sc_hd__buf_4 _18486_ (.A(_02536_),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _18487_ (.A0(\rbzero.wall_tracer.rayAddendX[6] ),
    .A1(_02663_),
    .S(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__clkbuf_1 _18488_ (.A(net5892),
    .X(_00607_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(_02626_),
    .B(net3614),
    .Y(_02666_));
 sky130_fd_sc_hd__or2_1 _18490_ (.A(_02626_),
    .B(net3614),
    .X(_02667_));
 sky130_fd_sc_hd__inv_2 _18491_ (.A(_02653_),
    .Y(_02668_));
 sky130_fd_sc_hd__o21a_1 _18492_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .B1(_02617_),
    .X(_02669_));
 sky130_fd_sc_hd__a311o_1 _18493_ (.A1(_02642_),
    .A2(_02643_),
    .A3(_02668_),
    .B1(net4867),
    .C1(net4820),
    .X(_02670_));
 sky130_fd_sc_hd__a21o_1 _18494_ (.A1(_02666_),
    .A2(_02667_),
    .B1(net4868),
    .X(_02671_));
 sky130_fd_sc_hd__nand3_1 _18495_ (.A(net8257),
    .B(_02667_),
    .C(net4868),
    .Y(_02672_));
 sky130_fd_sc_hd__or2_1 _18496_ (.A(_02626_),
    .B(net4554),
    .X(_02673_));
 sky130_fd_sc_hd__nand2_1 _18497_ (.A(_02626_),
    .B(net4554),
    .Y(_02674_));
 sky130_fd_sc_hd__a21bo_1 _18498_ (.A1(_02673_),
    .A2(_02674_),
    .B1_N(_02656_),
    .X(_02675_));
 sky130_fd_sc_hd__or3b_2 _18499_ (.A(_02626_),
    .B(net3494),
    .C_N(net4554),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_1 _18500_ (.A(_02675_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__a21bo_1 _18501_ (.A1(_02658_),
    .A2(_02661_),
    .B1_N(_02659_),
    .X(_02678_));
 sky130_fd_sc_hd__xnor2_1 _18502_ (.A(_02677_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__a22o_1 _18503_ (.A1(net3614),
    .A2(_09736_),
    .B1(_02679_),
    .B2(_04490_),
    .X(_02680_));
 sky130_fd_sc_hd__a31o_1 _18504_ (.A1(_02559_),
    .A2(net4869),
    .A3(net8258),
    .B1(net3615),
    .X(_00608_));
 sky130_fd_sc_hd__nand2_1 _18505_ (.A(_02627_),
    .B(net6015),
    .Y(_02681_));
 sky130_fd_sc_hd__or2_1 _18506_ (.A(_02626_),
    .B(net6015),
    .X(_02682_));
 sky130_fd_sc_hd__nand2_1 _18507_ (.A(_02681_),
    .B(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__a21oi_1 _18508_ (.A1(_02666_),
    .A2(_02672_),
    .B1(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__a31o_1 _18509_ (.A1(_02666_),
    .A2(_02672_),
    .A3(_02683_),
    .B1(_04489_),
    .X(_02685_));
 sky130_fd_sc_hd__or2b_1 _18510_ (.A(_02677_),
    .B_N(_02678_),
    .X(_02686_));
 sky130_fd_sc_hd__or2_1 _18511_ (.A(_02627_),
    .B(net4603),
    .X(_02687_));
 sky130_fd_sc_hd__nand2_1 _18512_ (.A(_02627_),
    .B(net4603),
    .Y(_02688_));
 sky130_fd_sc_hd__nand2_1 _18513_ (.A(_02687_),
    .B(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__xnor2_1 _18514_ (.A(_02673_),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__a21oi_2 _18515_ (.A1(_02676_),
    .A2(_02686_),
    .B1(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__a31o_1 _18516_ (.A1(_02676_),
    .A2(_02686_),
    .A3(_02690_),
    .B1(_04480_),
    .X(_02692_));
 sky130_fd_sc_hd__o22ai_1 _18517_ (.A1(_02684_),
    .A2(_02685_),
    .B1(_02691_),
    .B2(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__mux2_1 _18518_ (.A0(net6015),
    .A1(_02693_),
    .S(_02664_),
    .X(_02694_));
 sky130_fd_sc_hd__clkbuf_1 _18519_ (.A(net6017),
    .X(_00609_));
 sky130_fd_sc_hd__or2_1 _18520_ (.A(_02627_),
    .B(net4828),
    .X(_02695_));
 sky130_fd_sc_hd__nand2_1 _18521_ (.A(_02627_),
    .B(net4828),
    .Y(_02696_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(_02695_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__o211a_1 _18523_ (.A1(net8258),
    .A2(_02683_),
    .B1(_02681_),
    .C1(net8257),
    .X(_02698_));
 sky130_fd_sc_hd__xor2_1 _18524_ (.A(_02697_),
    .B(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__a211oi_1 _18525_ (.A1(net4603),
    .A2(net4554),
    .B1(_02691_),
    .C1(_02627_),
    .Y(_02700_));
 sky130_fd_sc_hd__a211o_1 _18526_ (.A1(_02687_),
    .A2(_02691_),
    .B1(net8260),
    .C1(_04482_),
    .X(_02701_));
 sky130_fd_sc_hd__o221a_1 _18527_ (.A1(net4828),
    .A2(_02537_),
    .B1(_09747_),
    .B2(_02699_),
    .C1(_02701_),
    .X(_00610_));
 sky130_fd_sc_hd__o21ai_1 _18528_ (.A1(_02697_),
    .A2(_02698_),
    .B1(_02696_),
    .Y(_02702_));
 sky130_fd_sc_hd__xor2_1 _18529_ (.A(_02627_),
    .B(net5952),
    .X(_02703_));
 sky130_fd_sc_hd__xnor2_1 _18530_ (.A(_02702_),
    .B(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__inv_2 _18531_ (.A(net4603),
    .Y(_02705_));
 sky130_fd_sc_hd__a211o_1 _18532_ (.A1(_02705_),
    .A2(_02691_),
    .B1(_04480_),
    .C1(_02627_),
    .X(_02706_));
 sky130_fd_sc_hd__o21ai_1 _18533_ (.A1(_04490_),
    .A2(_02704_),
    .B1(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__mux2_1 _18534_ (.A0(net5952),
    .A1(_02707_),
    .S(_02664_),
    .X(_02708_));
 sky130_fd_sc_hd__clkbuf_1 _18535_ (.A(net5954),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _18536_ (.A0(net7690),
    .A1(_06061_),
    .S(_02245_),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_1 _18537_ (.A0(_02709_),
    .A1(net5974),
    .S(_06242_),
    .X(_02710_));
 sky130_fd_sc_hd__clkbuf_1 _18538_ (.A(net3894),
    .X(_00612_));
 sky130_fd_sc_hd__nor2_1 _18539_ (.A(net3893),
    .B(_06041_),
    .Y(_02711_));
 sky130_fd_sc_hd__or3_1 _18540_ (.A(_08103_),
    .B(_06042_),
    .C(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_1 _18541_ (.A1(net4053),
    .A2(_09788_),
    .B1(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__mux2_1 _18542_ (.A0(net4054),
    .A1(_06039_),
    .S(_06242_),
    .X(_02714_));
 sky130_fd_sc_hd__clkbuf_1 _18543_ (.A(net4055),
    .X(_00613_));
 sky130_fd_sc_hd__or3_1 _18544_ (.A(_06038_),
    .B(_06042_),
    .C(_06044_),
    .X(_02715_));
 sky130_fd_sc_hd__nor2_1 _18545_ (.A(_06057_),
    .B(_06045_),
    .Y(_02716_));
 sky130_fd_sc_hd__a22o_1 _18546_ (.A1(net4436),
    .A2(_09818_),
    .B1(_02715_),
    .B2(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__mux2_1 _18547_ (.A0(_02717_),
    .A1(net5933),
    .S(_06242_),
    .X(_02718_));
 sky130_fd_sc_hd__clkbuf_1 _18548_ (.A(net5935),
    .X(_00614_));
 sky130_fd_sc_hd__or2b_1 _18549_ (.A(_06034_),
    .B_N(_06036_),
    .X(_02719_));
 sky130_fd_sc_hd__xnor2_1 _18550_ (.A(_06046_),
    .B(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__mux2_1 _18551_ (.A0(net7635),
    .A1(_02720_),
    .S(_02245_),
    .X(_02721_));
 sky130_fd_sc_hd__mux2_1 _18552_ (.A0(net7636),
    .A1(net4044),
    .S(_06242_),
    .X(_02722_));
 sky130_fd_sc_hd__clkbuf_1 _18553_ (.A(net4045),
    .X(_00615_));
 sky130_fd_sc_hd__or3_1 _18554_ (.A(_06049_),
    .B(_06034_),
    .C(_06047_),
    .X(_02723_));
 sky130_fd_sc_hd__nor2_1 _18555_ (.A(_06057_),
    .B(_06050_),
    .Y(_02724_));
 sky130_fd_sc_hd__a22o_1 _18556_ (.A1(net3552),
    .A2(_09818_),
    .B1(_02723_),
    .B2(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__mux2_1 _18557_ (.A0(_02725_),
    .A1(net7669),
    .S(_06242_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_1 _18558_ (.A(net7671),
    .X(_00616_));
 sky130_fd_sc_hd__a21oi_1 _18559_ (.A1(net3807),
    .A2(_06244_),
    .B1(_06050_),
    .Y(_02727_));
 sky130_fd_sc_hd__xnor2_1 _18560_ (.A(_06031_),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__mux2_1 _18561_ (.A0(net3469),
    .A1(_02728_),
    .S(_02245_),
    .X(_02729_));
 sky130_fd_sc_hd__mux2_1 _18562_ (.A0(_02729_),
    .A1(net7575),
    .S(_06240_),
    .X(_02730_));
 sky130_fd_sc_hd__clkbuf_1 _18563_ (.A(net7577),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _18564_ (.A0(net3443),
    .A1(net3960),
    .S(_02245_),
    .X(_02731_));
 sky130_fd_sc_hd__mux2_1 _18565_ (.A0(net3961),
    .A1(_06104_),
    .S(_10260_),
    .X(_02732_));
 sky130_fd_sc_hd__clkbuf_1 _18566_ (.A(net3962),
    .X(_00618_));
 sky130_fd_sc_hd__nor2_1 _18567_ (.A(_06104_),
    .B(net7713),
    .Y(_02733_));
 sky130_fd_sc_hd__or3_1 _18568_ (.A(_08103_),
    .B(_09755_),
    .C(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__o21ai_1 _18569_ (.A1(net3991),
    .A2(_09788_),
    .B1(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__mux2_1 _18570_ (.A0(net7714),
    .A1(net4034),
    .S(net4648),
    .X(_02736_));
 sky130_fd_sc_hd__clkbuf_1 _18571_ (.A(net4035),
    .X(_00619_));
 sky130_fd_sc_hd__xnor2_1 _18572_ (.A(_09756_),
    .B(_09759_),
    .Y(_02737_));
 sky130_fd_sc_hd__mux2_1 _18573_ (.A0(net5916),
    .A1(_02737_),
    .S(_09788_),
    .X(_02738_));
 sky130_fd_sc_hd__nor2_1 _18574_ (.A(_09769_),
    .B(net5917),
    .Y(_02739_));
 sky130_fd_sc_hd__a21o_1 _18575_ (.A1(net3965),
    .A2(_09769_),
    .B1(net5918),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _18576_ (.A(_09761_),
    .B(_09753_),
    .Y(_02740_));
 sky130_fd_sc_hd__xnor2_1 _18577_ (.A(_09760_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__mux2_1 _18578_ (.A0(net7701),
    .A1(_02741_),
    .S(_02245_),
    .X(_02742_));
 sky130_fd_sc_hd__mux2_1 _18579_ (.A0(net7702),
    .A1(net3999),
    .S(net4648),
    .X(_02743_));
 sky130_fd_sc_hd__clkbuf_1 _18580_ (.A(net4000),
    .X(_00621_));
 sky130_fd_sc_hd__xor2_1 _18581_ (.A(_09752_),
    .B(_09762_),
    .X(_02744_));
 sky130_fd_sc_hd__mux2_1 _18582_ (.A0(net7705),
    .A1(_02744_),
    .S(net91),
    .X(_02745_));
 sky130_fd_sc_hd__mux2_1 _18583_ (.A0(net7706),
    .A1(net4049),
    .S(net4648),
    .X(_02746_));
 sky130_fd_sc_hd__clkbuf_1 _18584_ (.A(net4050),
    .X(_00622_));
 sky130_fd_sc_hd__a21oi_1 _18585_ (.A1(_06060_),
    .A2(_09103_),
    .B1(_09774_),
    .Y(_02747_));
 sky130_fd_sc_hd__xnor2_1 _18586_ (.A(_09751_),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__mux2_1 _18587_ (.A0(net4019),
    .A1(_02748_),
    .S(net89),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _18588_ (.A0(_02749_),
    .A1(net7631),
    .S(net4648),
    .X(_02750_));
 sky130_fd_sc_hd__clkbuf_1 _18589_ (.A(net7633),
    .X(_00623_));
 sky130_fd_sc_hd__nor2_1 _18590_ (.A(net4528),
    .B(net4848),
    .Y(_02751_));
 sky130_fd_sc_hd__nor2_1 _18591_ (.A(net4635),
    .B(net4879),
    .Y(_02752_));
 sky130_fd_sc_hd__nand2_1 _18592_ (.A(_05164_),
    .B(net681),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _18593_ (.A(net4423),
    .B(net652),
    .Y(_02754_));
 sky130_fd_sc_hd__or2_1 _18594_ (.A(net4598),
    .B(net681),
    .X(_02755_));
 sky130_fd_sc_hd__nand3b_1 _18595_ (.A_N(net4424),
    .B(net4599),
    .C(_02753_),
    .Y(_02756_));
 sky130_fd_sc_hd__and2_1 _18596_ (.A(_02753_),
    .B(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__nand2_1 _18597_ (.A(net4635),
    .B(net4879),
    .Y(_02758_));
 sky130_fd_sc_hd__o21a_1 _18598_ (.A1(_02752_),
    .A2(_02757_),
    .B1(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__nand2_1 _18599_ (.A(net4528),
    .B(net4848),
    .Y(_02760_));
 sky130_fd_sc_hd__o21a_1 _18600_ (.A1(_02751_),
    .A2(_02759_),
    .B1(net4529),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_1 _18601_ (.A(net3618),
    .X(_02762_));
 sky130_fd_sc_hd__nor2_1 _18602_ (.A(net3619),
    .B(net1002),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_1 _18603_ (.A(net3619),
    .B(net1002),
    .Y(_02764_));
 sky130_fd_sc_hd__or2b_1 _18604_ (.A(_02763_),
    .B_N(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__xor2_1 _18605_ (.A(net4530),
    .B(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__inv_2 _18606_ (.A(net4423),
    .Y(_02767_));
 sky130_fd_sc_hd__nor2_1 _18607_ (.A(_02767_),
    .B(_08038_),
    .Y(_02768_));
 sky130_fd_sc_hd__a221o_1 _18608_ (.A1(net8129),
    .A2(_02508_),
    .B1(_09739_),
    .B2(net4531),
    .C1(_02768_),
    .X(_00624_));
 sky130_fd_sc_hd__nand2_1 _18609_ (.A(_05164_),
    .B(net4423),
    .Y(_02769_));
 sky130_fd_sc_hd__or2_1 _18610_ (.A(_05164_),
    .B(net4423),
    .X(_02770_));
 sky130_fd_sc_hd__o21a_1 _18611_ (.A1(net4530),
    .A2(_02763_),
    .B1(_02764_),
    .X(_02771_));
 sky130_fd_sc_hd__nor2_1 _18612_ (.A(net3575),
    .B(net5925),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2_1 _18613_ (.A(net3575),
    .B(net5925),
    .Y(_02773_));
 sky130_fd_sc_hd__or2b_1 _18614_ (.A(_02772_),
    .B_N(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__or2_1 _18615_ (.A(_02771_),
    .B(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__a21oi_1 _18616_ (.A1(_02771_),
    .A2(_02774_),
    .B1(_04489_),
    .Y(_02776_));
 sky130_fd_sc_hd__a32o_1 _18617_ (.A1(_02526_),
    .A2(_02769_),
    .A3(_02770_),
    .B1(_02775_),
    .B2(_02776_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _18618_ (.A0(net5925),
    .A1(_02777_),
    .S(_02664_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_1 _18619_ (.A(net5927),
    .X(_00625_));
 sky130_fd_sc_hd__nand2_1 _18620_ (.A(net4635),
    .B(_02770_),
    .Y(_02779_));
 sky130_fd_sc_hd__or2_1 _18621_ (.A(net4635),
    .B(_02770_),
    .X(_02780_));
 sky130_fd_sc_hd__o21a_1 _18622_ (.A1(_02771_),
    .A2(_02772_),
    .B1(_02773_),
    .X(_02781_));
 sky130_fd_sc_hd__nor2_1 _18623_ (.A(net4686),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2_1 _18624_ (.A(net4686),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02783_));
 sky130_fd_sc_hd__or2b_1 _18625_ (.A(_02782_),
    .B_N(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__or2_1 _18626_ (.A(_02781_),
    .B(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__a21oi_1 _18627_ (.A1(_02781_),
    .A2(_02784_),
    .B1(_04489_),
    .Y(_02786_));
 sky130_fd_sc_hd__a32o_1 _18628_ (.A1(_02526_),
    .A2(_02779_),
    .A3(_02780_),
    .B1(_02785_),
    .B2(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _18629_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(_02787_),
    .S(_02664_),
    .X(_02788_));
 sky130_fd_sc_hd__clkbuf_1 _18630_ (.A(net5809),
    .X(_00626_));
 sky130_fd_sc_hd__or4_2 _18631_ (.A(net4528),
    .B(net4635),
    .C(_05164_),
    .D(net4423),
    .X(_02789_));
 sky130_fd_sc_hd__a21oi_1 _18632_ (.A1(net4528),
    .A2(_02780_),
    .B1(_04480_),
    .Y(_02790_));
 sky130_fd_sc_hd__o21ai_1 _18633_ (.A1(_02781_),
    .A2(_02782_),
    .B1(_02783_),
    .Y(_02791_));
 sky130_fd_sc_hd__clkbuf_1 _18634_ (.A(net3677),
    .X(_02792_));
 sky130_fd_sc_hd__nor2_1 _18635_ (.A(net3678),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_02793_));
 sky130_fd_sc_hd__and2_1 _18636_ (.A(net3677),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_02794_));
 sky130_fd_sc_hd__or2_1 _18637_ (.A(_02793_),
    .B(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__xnor2_1 _18638_ (.A(_02791_),
    .B(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__a22o_1 _18639_ (.A1(_02789_),
    .A2(_02790_),
    .B1(_02796_),
    .B2(_04481_),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _18640_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(_02797_),
    .S(_02664_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_1 _18641_ (.A(net5805),
    .X(_00627_));
 sky130_fd_sc_hd__o21a_1 _18642_ (.A1(net3678),
    .A2(\rbzero.wall_tracer.rayAddendY[-2] ),
    .B1(_02791_),
    .X(_02799_));
 sky130_fd_sc_hd__nand2_1 _18643_ (.A(net4560),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_02800_));
 sky130_fd_sc_hd__or2_1 _18644_ (.A(net4560),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02801_));
 sky130_fd_sc_hd__o211a_1 _18645_ (.A1(_02794_),
    .A2(net4771),
    .B1(net8025),
    .C1(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__inv_2 _18646_ (.A(net8026),
    .Y(_02803_));
 sky130_fd_sc_hd__a211o_1 _18647_ (.A1(_02801_),
    .A2(net8025),
    .B1(net4771),
    .C1(_02794_),
    .X(_02804_));
 sky130_fd_sc_hd__o31a_1 _18648_ (.A1(net4528),
    .A2(net4635),
    .A3(_05164_),
    .B1(_02767_),
    .X(_02805_));
 sky130_fd_sc_hd__or2_1 _18649_ (.A(net3619),
    .B(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__nand2_1 _18650_ (.A(net3619),
    .B(_02805_),
    .Y(_02807_));
 sky130_fd_sc_hd__a32o_1 _18651_ (.A1(_04490_),
    .A2(_02806_),
    .A3(_02807_),
    .B1(_09736_),
    .B2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02808_));
 sky130_fd_sc_hd__a31o_1 _18652_ (.A1(_02559_),
    .A2(net8027),
    .A3(net4772),
    .B1(net3534),
    .X(_00628_));
 sky130_fd_sc_hd__xor2_1 _18653_ (.A(net3575),
    .B(_05164_),
    .X(_02809_));
 sky130_fd_sc_hd__nand2_1 _18654_ (.A(net3619),
    .B(net4423),
    .Y(_02810_));
 sky130_fd_sc_hd__o21ai_1 _18655_ (.A1(net3619),
    .A2(_02789_),
    .B1(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__xnor2_1 _18656_ (.A(_02809_),
    .B(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__nand2_1 _18657_ (.A(net8025),
    .B(_02803_),
    .Y(_02813_));
 sky130_fd_sc_hd__or2_1 _18658_ (.A(net4709),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_02814_));
 sky130_fd_sc_hd__nand2_1 _18659_ (.A(net4709),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_02815_));
 sky130_fd_sc_hd__nand2_1 _18660_ (.A(_02814_),
    .B(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__xnor2_1 _18661_ (.A(_02813_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__mux2_1 _18662_ (.A0(_02812_),
    .A1(_02817_),
    .S(_04480_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _18663_ (.A0(\rbzero.wall_tracer.rayAddendY[0] ),
    .A1(_02818_),
    .S(_02664_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _18664_ (.A(net5796),
    .X(_00629_));
 sky130_fd_sc_hd__nand2_1 _18665_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_02820_));
 sky130_fd_sc_hd__or2_1 _18666_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_02821_));
 sky130_fd_sc_hd__a21bo_1 _18667_ (.A1(_02813_),
    .A2(_02814_),
    .B1_N(_02815_),
    .X(_02822_));
 sky130_fd_sc_hd__a21o_1 _18668_ (.A1(net4764),
    .A2(net8092),
    .B1(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__and3_1 _18669_ (.A(net4764),
    .B(net8092),
    .C(_02822_),
    .X(_02824_));
 sky130_fd_sc_hd__inv_2 _18670_ (.A(net8093),
    .Y(_02825_));
 sky130_fd_sc_hd__nor2_2 _18671_ (.A(net4686),
    .B(net4635),
    .Y(_02826_));
 sky130_fd_sc_hd__and2_1 _18672_ (.A(net4686),
    .B(net4635),
    .X(_02827_));
 sky130_fd_sc_hd__nor4_2 _18673_ (.A(net3575),
    .B(_05164_),
    .C(_02826_),
    .D(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__o22a_1 _18674_ (.A1(net3575),
    .A2(_05164_),
    .B1(_02826_),
    .B2(_02827_),
    .X(_02829_));
 sky130_fd_sc_hd__or2_1 _18675_ (.A(_02828_),
    .B(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__o2bb2a_1 _18676_ (.A1_N(_02809_),
    .A2_N(_02810_),
    .B1(net3619),
    .B2(_02789_),
    .X(_02831_));
 sky130_fd_sc_hd__nor2_1 _18677_ (.A(_02830_),
    .B(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21o_1 _18678_ (.A1(_02830_),
    .A2(_02831_),
    .B1(_04481_),
    .X(_02833_));
 sky130_fd_sc_hd__a2bb2o_1 _18679_ (.A1_N(_02832_),
    .A2_N(_02833_),
    .B1(\rbzero.wall_tracer.rayAddendY[1] ),
    .B2(_09735_),
    .X(_02834_));
 sky130_fd_sc_hd__a31o_1 _18680_ (.A1(_02559_),
    .A2(net4765),
    .A3(net8094),
    .B1(net3915),
    .X(_00630_));
 sky130_fd_sc_hd__xor2_1 _18681_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_02835_));
 sky130_fd_sc_hd__and2_1 _18682_ (.A(net4764),
    .B(_02825_),
    .X(_02836_));
 sky130_fd_sc_hd__xnor2_1 _18683_ (.A(_02835_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__xor2_2 _18684_ (.A(net3678),
    .B(net4528),
    .X(_02838_));
 sky130_fd_sc_hd__or3_1 _18685_ (.A(_02828_),
    .B(_02832_),
    .C(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__o21ai_2 _18686_ (.A1(_02828_),
    .A2(_02832_),
    .B1(_02838_),
    .Y(_02840_));
 sky130_fd_sc_hd__nand2_1 _18687_ (.A(_02839_),
    .B(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__xnor2_1 _18688_ (.A(_02826_),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__mux2_1 _18689_ (.A0(_02837_),
    .A1(_02842_),
    .S(_02526_),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _18690_ (.A0(\rbzero.wall_tracer.rayAddendY[2] ),
    .A1(_02843_),
    .S(_02664_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _18691_ (.A(net5856),
    .X(_00631_));
 sky130_fd_sc_hd__inv_2 _18692_ (.A(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02845_));
 sky130_fd_sc_hd__or2_1 _18693_ (.A(net4560),
    .B(net3619),
    .X(_02846_));
 sky130_fd_sc_hd__nand2_1 _18694_ (.A(net4560),
    .B(net3619),
    .Y(_02847_));
 sky130_fd_sc_hd__nand2_1 _18695_ (.A(_02846_),
    .B(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hd__or3_1 _18696_ (.A(net3678),
    .B(net4528),
    .C(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__o21ai_1 _18697_ (.A1(net3678),
    .A2(net4528),
    .B1(_02848_),
    .Y(_02850_));
 sky130_fd_sc_hd__nand2_1 _18698_ (.A(_02849_),
    .B(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__o21ai_1 _18699_ (.A1(_02832_),
    .A2(_02838_),
    .B1(_02826_),
    .Y(_02852_));
 sky130_fd_sc_hd__a21o_1 _18700_ (.A1(_02840_),
    .A2(_02852_),
    .B1(_02851_),
    .X(_02853_));
 sky130_fd_sc_hd__nand2_1 _18701_ (.A(_04490_),
    .B(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__a31o_1 _18702_ (.A1(_02840_),
    .A2(_02851_),
    .A3(_02852_),
    .B1(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_4 _18703_ (.A(net8241),
    .X(_02856_));
 sky130_fd_sc_hd__nand2_1 _18704_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02857_));
 sky130_fd_sc_hd__or2_1 _18705_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02858_));
 sky130_fd_sc_hd__o21a_1 _18706_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_02859_));
 sky130_fd_sc_hd__a21o_1 _18707_ (.A1(_02824_),
    .A2(_02835_),
    .B1(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__a21oi_1 _18708_ (.A1(net4797),
    .A2(_02858_),
    .B1(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__and3_1 _18709_ (.A(net4797),
    .B(_02858_),
    .C(_02860_),
    .X(_02862_));
 sky130_fd_sc_hd__or3_1 _18710_ (.A(_09747_),
    .B(net4798),
    .C(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__o211ai_1 _18711_ (.A1(net8113),
    .A2(_02537_),
    .B1(_02855_),
    .C1(net4799),
    .Y(_00632_));
 sky130_fd_sc_hd__xor2_1 _18712_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_02864_));
 sky130_fd_sc_hd__buf_2 _18713_ (.A(_02856_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_4 _18714_ (.A(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__a21oi_1 _18715_ (.A1(_02866_),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02862_),
    .Y(_02867_));
 sky130_fd_sc_hd__xnor2_1 _18716_ (.A(_02864_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__nor2_1 _18717_ (.A(net4709),
    .B(net3575),
    .Y(_02869_));
 sky130_fd_sc_hd__and2_1 _18718_ (.A(net4709),
    .B(net3575),
    .X(_02870_));
 sky130_fd_sc_hd__or2_1 _18719_ (.A(_02869_),
    .B(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__nand3_1 _18720_ (.A(_02849_),
    .B(_02853_),
    .C(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__a21o_1 _18721_ (.A1(_02849_),
    .A2(_02853_),
    .B1(_02871_),
    .X(_02873_));
 sky130_fd_sc_hd__a21oi_1 _18722_ (.A1(_02872_),
    .A2(_02873_),
    .B1(_02846_),
    .Y(_02874_));
 sky130_fd_sc_hd__and3_1 _18723_ (.A(_02846_),
    .B(_02872_),
    .C(_02873_),
    .X(_02875_));
 sky130_fd_sc_hd__or2_1 _18724_ (.A(_02874_),
    .B(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _18725_ (.A0(_02868_),
    .A1(_02876_),
    .S(_02526_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _18726_ (.A0(\rbzero.wall_tracer.rayAddendY[4] ),
    .A1(_02877_),
    .S(_02664_),
    .X(_02878_));
 sky130_fd_sc_hd__clkbuf_1 _18727_ (.A(net5777),
    .X(_00633_));
 sky130_fd_sc_hd__nand2_1 _18728_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_02879_));
 sky130_fd_sc_hd__or2_1 _18729_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_02880_));
 sky130_fd_sc_hd__and2_1 _18730_ (.A(net8060),
    .B(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__and2_1 _18731_ (.A(_02862_),
    .B(_02864_),
    .X(_02882_));
 sky130_fd_sc_hd__o21a_1 _18732_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02856_),
    .X(_02883_));
 sky130_fd_sc_hd__or3_1 _18733_ (.A(net8061),
    .B(_02882_),
    .C(net4807),
    .X(_02884_));
 sky130_fd_sc_hd__o21ai_1 _18734_ (.A1(_02882_),
    .A2(net4807),
    .B1(net8061),
    .Y(_02885_));
 sky130_fd_sc_hd__a21o_1 _18735_ (.A1(_02853_),
    .A2(_02871_),
    .B1(_02846_),
    .X(_02886_));
 sky130_fd_sc_hd__xor2_1 _18736_ (.A(_02856_),
    .B(net4686),
    .X(_02887_));
 sky130_fd_sc_hd__xnor2_1 _18737_ (.A(_02869_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__a21oi_1 _18738_ (.A1(_02873_),
    .A2(_02886_),
    .B1(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__a31o_1 _18739_ (.A1(_02873_),
    .A2(_02888_),
    .A3(_02886_),
    .B1(_04481_),
    .X(_02890_));
 sky130_fd_sc_hd__a2bb2o_1 _18740_ (.A1_N(_02889_),
    .A2_N(_02890_),
    .B1(\rbzero.wall_tracer.rayAddendY[5] ),
    .B2(_09735_),
    .X(_02891_));
 sky130_fd_sc_hd__a31o_1 _18741_ (.A1(_09739_),
    .A2(net4808),
    .A3(net8062),
    .B1(net3759),
    .X(_00634_));
 sky130_fd_sc_hd__xnor2_2 _18742_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_02892_));
 sky130_fd_sc_hd__a21oi_1 _18743_ (.A1(_02879_),
    .A2(_02885_),
    .B1(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__a31o_1 _18744_ (.A1(_02879_),
    .A2(_02885_),
    .A3(_02892_),
    .B1(_04478_),
    .X(_02894_));
 sky130_fd_sc_hd__or2_1 _18745_ (.A(_02856_),
    .B(net3678),
    .X(_02895_));
 sky130_fd_sc_hd__nand2_1 _18746_ (.A(_02865_),
    .B(net3678),
    .Y(_02896_));
 sky130_fd_sc_hd__a2bb2o_1 _18747_ (.A1_N(_02865_),
    .A2_N(net4686),
    .B1(_02895_),
    .B2(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__or3b_1 _18748_ (.A(_02865_),
    .B(net4686),
    .C_N(net3678),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_1 _18749_ (.A(_02897_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__a21o_1 _18750_ (.A1(_02869_),
    .A2(_02887_),
    .B1(_02889_),
    .X(_02900_));
 sky130_fd_sc_hd__xnor2_1 _18751_ (.A(_02899_),
    .B(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__a2bb2o_1 _18752_ (.A1_N(_02893_),
    .A2_N(_02894_),
    .B1(_02901_),
    .B2(_02526_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _18753_ (.A0(\rbzero.wall_tracer.rayAddendY[6] ),
    .A1(_02902_),
    .S(_02664_),
    .X(_02903_));
 sky130_fd_sc_hd__clkbuf_1 _18754_ (.A(net5842),
    .X(_00635_));
 sky130_fd_sc_hd__nand2_1 _18755_ (.A(_02865_),
    .B(net3761),
    .Y(_02904_));
 sky130_fd_sc_hd__or2_1 _18756_ (.A(_02865_),
    .B(net3761),
    .X(_02905_));
 sky130_fd_sc_hd__inv_2 _18757_ (.A(_02892_),
    .Y(_02906_));
 sky130_fd_sc_hd__o21a_1 _18758_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .B1(_02856_),
    .X(_02907_));
 sky130_fd_sc_hd__a311o_1 _18759_ (.A1(_02881_),
    .A2(_02882_),
    .A3(_02906_),
    .B1(net4856),
    .C1(net4807),
    .X(_02908_));
 sky130_fd_sc_hd__a21o_1 _18760_ (.A1(_02904_),
    .A2(_02905_),
    .B1(net4857),
    .X(_02909_));
 sky130_fd_sc_hd__nand3_1 _18761_ (.A(net8242),
    .B(_02905_),
    .C(net4857),
    .Y(_02910_));
 sky130_fd_sc_hd__or2_1 _18762_ (.A(_02865_),
    .B(net4560),
    .X(_02911_));
 sky130_fd_sc_hd__nand2_1 _18763_ (.A(_02865_),
    .B(net4560),
    .Y(_02912_));
 sky130_fd_sc_hd__a21bo_1 _18764_ (.A1(_02911_),
    .A2(_02912_),
    .B1_N(_02895_),
    .X(_02913_));
 sky130_fd_sc_hd__or3b_2 _18765_ (.A(_02865_),
    .B(net3678),
    .C_N(net4560),
    .X(_02914_));
 sky130_fd_sc_hd__nand2_1 _18766_ (.A(_02913_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__a21bo_1 _18767_ (.A1(_02897_),
    .A2(_02900_),
    .B1_N(_02898_),
    .X(_02916_));
 sky130_fd_sc_hd__xnor2_1 _18768_ (.A(_02915_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__a22o_1 _18769_ (.A1(net3761),
    .A2(_09736_),
    .B1(_02917_),
    .B2(_04490_),
    .X(_02918_));
 sky130_fd_sc_hd__a31o_1 _18770_ (.A1(_09739_),
    .A2(net4858),
    .A3(net8243),
    .B1(net3762),
    .X(_00636_));
 sky130_fd_sc_hd__nand2_1 _18771_ (.A(_02866_),
    .B(net6046),
    .Y(_02919_));
 sky130_fd_sc_hd__or2_1 _18772_ (.A(_02865_),
    .B(net6046),
    .X(_02920_));
 sky130_fd_sc_hd__nand2_1 _18773_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__a21oi_1 _18774_ (.A1(_02904_),
    .A2(_02910_),
    .B1(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__a31o_1 _18775_ (.A1(_02904_),
    .A2(_02910_),
    .A3(_02921_),
    .B1(_04489_),
    .X(_02923_));
 sky130_fd_sc_hd__or2b_1 _18776_ (.A(_02915_),
    .B_N(_02916_),
    .X(_02924_));
 sky130_fd_sc_hd__or2_1 _18777_ (.A(_02866_),
    .B(net4709),
    .X(_02925_));
 sky130_fd_sc_hd__nand2_1 _18778_ (.A(_02866_),
    .B(net4709),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_1 _18779_ (.A(_02925_),
    .B(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__xnor2_1 _18780_ (.A(_02911_),
    .B(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__a21oi_2 _18781_ (.A1(_02914_),
    .A2(_02924_),
    .B1(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__a31o_1 _18782_ (.A1(_02914_),
    .A2(_02924_),
    .A3(_02928_),
    .B1(_04480_),
    .X(_02930_));
 sky130_fd_sc_hd__o22ai_1 _18783_ (.A1(_02922_),
    .A2(_02923_),
    .B1(_02929_),
    .B2(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__mux2_1 _18784_ (.A0(net6046),
    .A1(_02931_),
    .S(_02536_),
    .X(_02932_));
 sky130_fd_sc_hd__clkbuf_1 _18785_ (.A(net6048),
    .X(_00637_));
 sky130_fd_sc_hd__or2_1 _18786_ (.A(_02866_),
    .B(net4838),
    .X(_02933_));
 sky130_fd_sc_hd__nand2_1 _18787_ (.A(_02866_),
    .B(net4838),
    .Y(_02934_));
 sky130_fd_sc_hd__nand2_1 _18788_ (.A(_02933_),
    .B(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__o211a_1 _18789_ (.A1(net8243),
    .A2(_02921_),
    .B1(_02919_),
    .C1(net8242),
    .X(_02936_));
 sky130_fd_sc_hd__xor2_1 _18790_ (.A(_02935_),
    .B(_02936_),
    .X(_02937_));
 sky130_fd_sc_hd__a211oi_1 _18791_ (.A1(net4709),
    .A2(net4560),
    .B1(_02929_),
    .C1(_02866_),
    .Y(_02938_));
 sky130_fd_sc_hd__a211o_1 _18792_ (.A1(_02925_),
    .A2(_02929_),
    .B1(net8246),
    .C1(_04482_),
    .X(_02939_));
 sky130_fd_sc_hd__o221a_1 _18793_ (.A1(net4838),
    .A2(_02537_),
    .B1(_09747_),
    .B2(_02937_),
    .C1(net8247),
    .X(_00638_));
 sky130_fd_sc_hd__o21ai_1 _18794_ (.A1(_02935_),
    .A2(_02936_),
    .B1(_02934_),
    .Y(_02940_));
 sky130_fd_sc_hd__xor2_1 _18795_ (.A(_02866_),
    .B(net5955),
    .X(_02941_));
 sky130_fd_sc_hd__xnor2_1 _18796_ (.A(_02940_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__inv_2 _18797_ (.A(net4709),
    .Y(_02943_));
 sky130_fd_sc_hd__a211o_1 _18798_ (.A1(_02943_),
    .A2(_02929_),
    .B1(_04480_),
    .C1(_02866_),
    .X(_02944_));
 sky130_fd_sc_hd__o21ai_1 _18799_ (.A1(_04490_),
    .A2(_02942_),
    .B1(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__mux2_1 _18800_ (.A0(net5955),
    .A1(_02945_),
    .S(_02536_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _18801_ (.A(net5957),
    .X(_00639_));
 sky130_fd_sc_hd__and2b_2 _18802_ (.A_N(net5863),
    .B(net7496),
    .X(_02947_));
 sky130_fd_sc_hd__and2b_1 _18803_ (.A_N(net4814),
    .B(net3940),
    .X(_02948_));
 sky130_fd_sc_hd__nand2_1 _18804_ (.A(net1878),
    .B(net3083),
    .Y(_02949_));
 sky130_fd_sc_hd__and3b_1 _18805_ (.A_N(net3940),
    .B(net4814),
    .C(net3084),
    .X(_02950_));
 sky130_fd_sc_hd__a21oi_2 _18806_ (.A1(net4832),
    .A2(_02948_),
    .B1(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__nor2_1 _18807_ (.A(net3485),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__or3_1 _18808_ (.A(net3695),
    .B(net5799),
    .C(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__or2_2 _18809_ (.A(net3770),
    .B(net4832),
    .X(_02954_));
 sky130_fd_sc_hd__a21oi_2 _18810_ (.A1(net3940),
    .A2(_02954_),
    .B1(net4814),
    .Y(_02955_));
 sky130_fd_sc_hd__nor2_1 _18811_ (.A(net1547),
    .B(net3909),
    .Y(_02956_));
 sky130_fd_sc_hd__o21a_1 _18812_ (.A1(net3851),
    .A2(net4814),
    .B1(net1547),
    .X(_02957_));
 sky130_fd_sc_hd__a21oi_1 _18813_ (.A1(net3084),
    .A2(_02955_),
    .B1(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__o311a_1 _18814_ (.A1(net1547),
    .A2(net3851),
    .A3(net4814),
    .B1(_02958_),
    .C1(net3909),
    .X(_02959_));
 sky130_fd_sc_hd__a31o_1 _18815_ (.A1(net3084),
    .A2(_02955_),
    .A3(_02956_),
    .B1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__or2b_1 _18816_ (.A(_02955_),
    .B_N(_02951_),
    .X(_02961_));
 sky130_fd_sc_hd__nor3_1 _18817_ (.A(net3909),
    .B(net5845),
    .C(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__a32o_1 _18818_ (.A1(net5845),
    .A2(_02960_),
    .A3(_02961_),
    .B1(_02962_),
    .B2(net1547),
    .X(_02963_));
 sky130_fd_sc_hd__a311o_1 _18819_ (.A1(net3770),
    .A2(_02472_),
    .A3(_02948_),
    .B1(_02955_),
    .C1(_02950_),
    .X(_02964_));
 sky130_fd_sc_hd__xnor2_1 _18820_ (.A(net3935),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_1 _18821_ (.A(_02963_),
    .B(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__a211o_1 _18822_ (.A1(net3485),
    .A2(_02951_),
    .B1(_02953_),
    .C1(net7695),
    .X(_02967_));
 sky130_fd_sc_hd__and2_1 _18823_ (.A(_02947_),
    .B(net3486),
    .X(_02968_));
 sky130_fd_sc_hd__nor2_2 _18824_ (.A(net4062),
    .B(_04102_),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2_1 _18825_ (.A(net5845),
    .B(_02947_),
    .Y(_02970_));
 sky130_fd_sc_hd__o211a_1 _18826_ (.A1(net5845),
    .A2(_02968_),
    .B1(net4063),
    .C1(net2199),
    .X(_00640_));
 sky130_fd_sc_hd__nand2_1 _18827_ (.A(net5877),
    .B(net5845),
    .Y(_02971_));
 sky130_fd_sc_hd__or2b_1 _18828_ (.A(net5863),
    .B_N(net2182),
    .X(_02972_));
 sky130_fd_sc_hd__a21o_1 _18829_ (.A1(net3486),
    .A2(_02971_),
    .B1(net5864),
    .X(_02973_));
 sky130_fd_sc_hd__a21o_1 _18830_ (.A1(net2198),
    .A2(_02947_),
    .B1(net3909),
    .X(_02974_));
 sky130_fd_sc_hd__and3_1 _18831_ (.A(_02969_),
    .B(_02973_),
    .C(net3910),
    .X(_02975_));
 sky130_fd_sc_hd__clkbuf_1 _18832_ (.A(net3911),
    .X(_00641_));
 sky130_fd_sc_hd__or3b_1 _18833_ (.A(net5878),
    .B(net1547),
    .C_N(_02968_),
    .X(_02976_));
 sky130_fd_sc_hd__nand2_1 _18834_ (.A(net1547),
    .B(_02973_),
    .Y(_02977_));
 sky130_fd_sc_hd__a21boi_1 _18835_ (.A1(net5879),
    .A2(net1548),
    .B1_N(net4063),
    .Y(_00642_));
 sky130_fd_sc_hd__a31o_1 _18836_ (.A1(net1547),
    .A2(net3909),
    .A3(net2198),
    .B1(net3935),
    .X(_02978_));
 sky130_fd_sc_hd__and4_1 _18837_ (.A(net3935),
    .B(net1547),
    .C(net3909),
    .D(net5845),
    .X(_02979_));
 sky130_fd_sc_hd__inv_2 _18838_ (.A(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__a32o_1 _18839_ (.A1(_02968_),
    .A2(_02978_),
    .A3(_02980_),
    .B1(net5864),
    .B2(net3935),
    .X(_02981_));
 sky130_fd_sc_hd__and2_1 _18840_ (.A(_02969_),
    .B(net3936),
    .X(_02982_));
 sky130_fd_sc_hd__clkbuf_1 _18841_ (.A(net3937),
    .X(_00643_));
 sky130_fd_sc_hd__and3_1 _18842_ (.A(net3485),
    .B(_02947_),
    .C(_02979_),
    .X(_02983_));
 sky130_fd_sc_hd__a21o_1 _18843_ (.A1(_02947_),
    .A2(_02979_),
    .B1(net3485),
    .X(_02984_));
 sky130_fd_sc_hd__and3b_1 _18844_ (.A_N(_02983_),
    .B(net4063),
    .C(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__o21a_1 _18845_ (.A1(net5864),
    .A2(net3486),
    .B1(_02985_),
    .X(_00644_));
 sky130_fd_sc_hd__and2_1 _18846_ (.A(net5799),
    .B(_02983_),
    .X(_02986_));
 sky130_fd_sc_hd__o21ai_1 _18847_ (.A1(net5799),
    .A2(_02983_),
    .B1(_02969_),
    .Y(_02987_));
 sky130_fd_sc_hd__nor2_1 _18848_ (.A(net5800),
    .B(net1251),
    .Y(_00645_));
 sky130_fd_sc_hd__nand2_1 _18849_ (.A(net3695),
    .B(_02986_),
    .Y(_02988_));
 sky130_fd_sc_hd__or2_1 _18850_ (.A(net3695),
    .B(net5800),
    .X(_02989_));
 sky130_fd_sc_hd__and3_1 _18851_ (.A(_02969_),
    .B(net3696),
    .C(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__clkbuf_1 _18852_ (.A(net3697),
    .X(_00646_));
 sky130_fd_sc_hd__nand2_1 _18853_ (.A(net3950),
    .B(net92),
    .Y(_02991_));
 sky130_fd_sc_hd__buf_4 _18854_ (.A(net2873),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_4 _18855_ (.A(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _18856_ (.A0(net3329),
    .A1(net4591),
    .S(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_1 _18857_ (.A(net3330),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18858_ (.A0(net3351),
    .A1(net4825),
    .S(_02993_),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_1 _18859_ (.A(net3352),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _18860_ (.A0(net2764),
    .A1(net7419),
    .S(_02993_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_1 _18861_ (.A(net7421),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18862_ (.A0(net3045),
    .A1(net6681),
    .S(_02993_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_1 _18863_ (.A(net1863),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _18864_ (.A0(net6413),
    .A1(net6560),
    .S(_02993_),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_1 _18865_ (.A(net1574),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _18866_ (.A0(net6661),
    .A1(net7003),
    .S(_02993_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _18867_ (.A(net1971),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _18868_ (.A0(net1682),
    .A1(net6693),
    .S(_02993_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_1 _18869_ (.A(net6695),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18870_ (.A0(net3026),
    .A1(net7538),
    .S(_02993_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_1 _18871_ (.A(net2469),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _18872_ (.A0(net3019),
    .A1(net7490),
    .S(_02993_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_1 _18873_ (.A(net3020),
    .X(_00655_));
 sky130_fd_sc_hd__clkbuf_4 _18874_ (.A(_02992_),
    .X(_03003_));
 sky130_fd_sc_hd__mux2_1 _18875_ (.A0(net3145),
    .A1(net7508),
    .S(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_1 _18876_ (.A(net2957),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _18877_ (.A0(net3111),
    .A1(net5045),
    .S(_03003_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_1 _18878_ (.A(net3112),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _18879_ (.A0(net2869),
    .A1(net7409),
    .S(_03003_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_1 _18880_ (.A(net7411),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _18881_ (.A0(net2771),
    .A1(net4803),
    .S(_03003_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _18882_ (.A(net1195),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _18883_ (.A0(net6231),
    .A1(net638),
    .S(_03003_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _18884_ (.A(net6233),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _18885_ (.A0(net6247),
    .A1(net2079),
    .S(_03003_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _18886_ (.A(net2080),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _18887_ (.A0(net3077),
    .A1(net7021),
    .S(_03003_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_1 _18888_ (.A(net2162),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _18889_ (.A0(net3063),
    .A1(net7045),
    .S(_03003_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_1 _18890_ (.A(net7047),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _18891_ (.A0(net1752),
    .A1(net7155),
    .S(_03003_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _18892_ (.A(net1753),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _18893_ (.A0(net3155),
    .A1(net6707),
    .S(_03003_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _18894_ (.A(net6709),
    .X(_00665_));
 sky130_fd_sc_hd__clkbuf_4 _18895_ (.A(_02992_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _18896_ (.A0(net6125),
    .A1(net2364),
    .S(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_1 _18897_ (.A(net2365),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _18898_ (.A0(net3186),
    .A1(net7188),
    .S(_03014_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_1 _18899_ (.A(net1947),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _18900_ (.A0(net3056),
    .A1(net5476),
    .S(_03014_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_1 _18901_ (.A(net3057),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _18902_ (.A0(net7443),
    .A1(net3182),
    .S(_03014_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _18903_ (.A(net7445),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _18904_ (.A0(net6512),
    .A1(net1057),
    .S(_03014_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _18905_ (.A(net6514),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _18906_ (.A0(net3173),
    .A1(net7548),
    .S(_03014_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_1 _18907_ (.A(net3290),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _18908_ (.A0(net6649),
    .A1(net6954),
    .S(_03014_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_1 _18909_ (.A(net2486),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _18910_ (.A0(net6357),
    .A1(net7143),
    .S(_03014_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_1 _18911_ (.A(net1916),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _18912_ (.A0(net3195),
    .A1(net7552),
    .S(_03014_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_1 _18913_ (.A(net3196),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _18914_ (.A0(net3179),
    .A1(net7544),
    .S(_03014_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _18915_ (.A(net7546),
    .X(_00675_));
 sky130_fd_sc_hd__clkbuf_4 _18916_ (.A(_02992_),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_1 _18917_ (.A0(net3342),
    .A1(net7583),
    .S(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_1 _18918_ (.A(net3293),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _18919_ (.A0(net3302),
    .A1(net7565),
    .S(_03025_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_1 _18920_ (.A(net3208),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _18921_ (.A0(net7516),
    .A1(net7550),
    .S(_03025_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _18922_ (.A(net3277),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _18923_ (.A0(net3256),
    .A1(net7613),
    .S(_03025_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _18924_ (.A(net3081),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _18925_ (.A0(net6436),
    .A1(net3407),
    .S(_03025_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _18926_ (.A(net6438),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _18927_ (.A0(net3273),
    .A1(net7595),
    .S(_03025_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _18928_ (.A(net3274),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _18929_ (.A0(net3298),
    .A1(net7593),
    .S(_03025_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _18930_ (.A(net1647),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _18931_ (.A0(net3125),
    .A1(net3362),
    .S(_03025_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _18932_ (.A(net3363),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _18933_ (.A0(net6731),
    .A1(net3435),
    .S(_03025_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _18934_ (.A(net6733),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _18935_ (.A0(net2934),
    .A1(net7481),
    .S(_03025_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _18936_ (.A(net1103),
    .X(_00685_));
 sky130_fd_sc_hd__clkbuf_4 _18937_ (.A(_02992_),
    .X(_03036_));
 sky130_fd_sc_hd__mux2_1 _18938_ (.A0(net3320),
    .A1(net6878),
    .S(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_1 _18939_ (.A(net1933),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _18940_ (.A0(net3214),
    .A1(net7334),
    .S(_03036_),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_1 _18941_ (.A(net2585),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _18942_ (.A0(net3166),
    .A1(net7461),
    .S(_03036_),
    .X(_03039_));
 sky130_fd_sc_hd__clkbuf_1 _18943_ (.A(net7463),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _18944_ (.A0(net3260),
    .A1(net7093),
    .S(_03036_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _18945_ (.A(net2331),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _18946_ (.A0(net2974),
    .A1(net7083),
    .S(_03036_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _18947_ (.A(net2089),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _18948_ (.A0(net7178),
    .A1(net3440),
    .S(_03036_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _18949_ (.A(net2759),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _18950_ (.A0(net3138),
    .A1(net5704),
    .S(_03036_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _18951_ (.A(net2839),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _18952_ (.A0(net7453),
    .A1(net7471),
    .S(_03036_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_1 _18953_ (.A(net3253),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _18954_ (.A0(net6744),
    .A1(net5750),
    .S(_03036_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _18955_ (.A(net1907),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _18956_ (.A0(net2801),
    .A1(net7573),
    .S(_03036_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _18957_ (.A(net1146),
    .X(_00695_));
 sky130_fd_sc_hd__clkbuf_1 _18958_ (.A(net2873),
    .X(_03047_));
 sky130_fd_sc_hd__mux2_1 _18959_ (.A0(net3227),
    .A1(net5743),
    .S(net2874),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _18960_ (.A(net1789),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _18961_ (.A0(net5710),
    .A1(net4327),
    .S(net2874),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _18962_ (.A(net5712),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _18963_ (.A0(net7367),
    .A1(net5771),
    .S(net2874),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_1 _18964_ (.A(net3324),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _18965_ (.A0(net3052),
    .A1(net7567),
    .S(net2874),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _18966_ (.A(net2875),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _18967_ (.A0(net6201),
    .A1(net4901),
    .S(net2874),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _18968_ (.A(net2427),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _18969_ (.A0(net3121),
    .A1(net6687),
    .S(net2874),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _18970_ (.A(net1559),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _18971_ (.A0(net2829),
    .A1(net7465),
    .S(net2874),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _18972_ (.A(net7467),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _18973_ (.A0(net3312),
    .A1(net5737),
    .S(net2874),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _18974_ (.A(net3224),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _18975_ (.A0(net3283),
    .A1(net6061),
    .S(net2874),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _18976_ (.A(net3039),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _18977_ (.A0(net3060),
    .A1(net5733),
    .S(net2874),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _18978_ (.A(net5735),
    .X(_00705_));
 sky130_fd_sc_hd__clkbuf_4 _18979_ (.A(net2873),
    .X(_03058_));
 sky130_fd_sc_hd__mux2_1 _18980_ (.A0(net7455),
    .A1(net5745),
    .S(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_1 _18981_ (.A(net3099),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _18982_ (.A0(net6239),
    .A1(net5816),
    .S(_03058_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_1 _18983_ (.A(net1536),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _18984_ (.A0(net7520),
    .A1(net5835),
    .S(_03058_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_1 _18985_ (.A(net3412),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _18986_ (.A0(net7449),
    .A1(net7536),
    .S(_03058_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_1 _18987_ (.A(net3270),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _18988_ (.A0(net3159),
    .A1(net7587),
    .S(_03058_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _18989_ (.A(net1472),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _18990_ (.A0(net2927),
    .A1(net5783),
    .S(_03058_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _18991_ (.A(net2864),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _18992_ (.A0(net7175),
    .A1(net5849),
    .S(_03058_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _18993_ (.A(net3267),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _18994_ (.A0(net5812),
    .A1(net4490),
    .S(_03058_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _18995_ (.A(net5814),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _18996_ (.A0(net3009),
    .A1(net5826),
    .S(_03058_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _18997_ (.A(net1704),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _18998_ (.A0(net5988),
    .A1(net5868),
    .S(_03058_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _18999_ (.A(net3280),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _19000_ (.A0(net3237),
    .A1(net5791),
    .S(_02992_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _19001_ (.A(net5793),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _19002_ (.A0(net5764),
    .A1(net4454),
    .S(_02992_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _19003_ (.A(net5766),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _19004_ (.A0(net6327),
    .A1(net5898),
    .S(_02992_),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_1 _19005_ (.A(net3016),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _19006_ (.A0(net7510),
    .A1(net3345),
    .S(_02992_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _19007_ (.A(net7512),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _19008_ (.A0(net1613),
    .A1(net5784),
    .S(_02992_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _19009_ (.A(net5786),
    .X(_00720_));
 sky130_fd_sc_hd__or3_1 _19010_ (.A(net3485),
    .B(net3935),
    .C(net1547),
    .X(_03074_));
 sky130_fd_sc_hd__nor3_1 _19011_ (.A(net3695),
    .B(net1250),
    .C(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__or3b_1 _19012_ (.A(_02972_),
    .B(net3395),
    .C_N(_02969_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _19013_ (.A(net3396),
    .X(_03077_));
 sky130_fd_sc_hd__buf_4 _19014_ (.A(net3397),
    .X(_03078_));
 sky130_fd_sc_hd__mux2_1 _19015_ (.A0(net3793),
    .A1(net3899),
    .S(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _19016_ (.A(net3900),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _19017_ (.A0(net3899),
    .A1(net4030),
    .S(_03078_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _19018_ (.A(_03080_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _19019_ (.A0(net4030),
    .A1(net1493),
    .S(_03078_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _19020_ (.A(net4031),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _19021_ (.A0(net1493),
    .A1(net4076),
    .S(_03078_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _19022_ (.A(net4077),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _19023_ (.A0(net1426),
    .A1(net4016),
    .S(_03078_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _19024_ (.A(net4017),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _19025_ (.A0(net4040),
    .A1(net2205),
    .S(_03078_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_1 _19026_ (.A(net4041),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _19027_ (.A0(net2205),
    .A1(net3863),
    .S(_03078_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _19028_ (.A(net3864),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _19029_ (.A0(net3863),
    .A1(net3816),
    .S(_03078_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _19030_ (.A(net3878),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _19031_ (.A0(net3816),
    .A1(net3402),
    .S(_03078_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _19032_ (.A(net3817),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _19033_ (.A0(net3402),
    .A1(net7698),
    .S(_03078_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_1 _19034_ (.A(net3403),
    .X(_00730_));
 sky130_fd_sc_hd__buf_1 _19035_ (.A(net3397),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _19036_ (.A0(net7698),
    .A1(net3838),
    .S(net3398),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _19037_ (.A(net3839),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _19038_ (.A0(net3838),
    .A1(net3745),
    .S(net3398),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _19039_ (.A(net3746),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _19040_ (.A0(net3745),
    .A1(net3596),
    .S(net3398),
    .X(_03092_));
 sky130_fd_sc_hd__clkbuf_1 _19041_ (.A(net3399),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _19042_ (.A0(net3596),
    .A1(net3562),
    .S(net3398),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _19043_ (.A(net3597),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _19044_ (.A0(net3562),
    .A1(net3738),
    .S(net3398),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_1 _19045_ (.A(net3563),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _19046_ (.A0(net3738),
    .A1(net7621),
    .S(net3398),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_1 _19047_ (.A(net3739),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _19048_ (.A0(net7621),
    .A1(net7589),
    .S(net3398),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _19049_ (.A(net3593),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _19050_ (.A0(net7589),
    .A1(net3674),
    .S(net3398),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _19051_ (.A(net7591),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _19052_ (.A0(net7615),
    .A1(net3866),
    .S(net3398),
    .X(_03098_));
 sky130_fd_sc_hd__clkbuf_1 _19053_ (.A(net7617),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _19054_ (.A0(net7629),
    .A1(net7585),
    .S(net3398),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _19055_ (.A(net3867),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _19056_ (.A0(net7585),
    .A1(net7579),
    .S(net3397),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _19057_ (.A(net3479),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _19058_ (.A0(net7579),
    .A1(net3481),
    .S(net3397),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_1 _19059_ (.A(net7581),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _19060_ (.A0(net7597),
    .A1(net3583),
    .S(net3397),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _19061_ (.A(net7599),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _19062_ (.A0(net7601),
    .A1(net3631),
    .S(net3397),
    .X(_03103_));
 sky130_fd_sc_hd__clkbuf_1 _19063_ (.A(net7603),
    .X(_00744_));
 sky130_fd_sc_hd__and3_2 _19064_ (.A(_02947_),
    .B(_02969_),
    .C(net3395),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _19065_ (.A0(net3770),
    .A1(net3793),
    .S(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _19066_ (.A(net3794),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _19067_ (.A0(_02472_),
    .A1(net3770),
    .S(_03104_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _19068_ (.A(net3771),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _19069_ (.A0(net3940),
    .A1(_02472_),
    .S(_03104_),
    .X(_03107_));
 sky130_fd_sc_hd__clkbuf_1 _19070_ (.A(net3941),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _19071_ (.A0(net5895),
    .A1(net3940),
    .S(_03104_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _19072_ (.A(net3852),
    .X(_00748_));
 sky130_fd_sc_hd__buf_4 _19073_ (.A(_04458_),
    .X(_03109_));
 sky130_fd_sc_hd__mux2_1 _19074_ (.A0(net44),
    .A1(net6611),
    .S(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _19075_ (.A(net1728),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _19076_ (.A0(net3793),
    .A1(net6611),
    .S(_09725_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _19077_ (.A(net2047),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _19078_ (.A0(net43),
    .A1(net7277),
    .S(_03109_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _19079_ (.A(net2436),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _19080_ (.A0(net4062),
    .A1(net7277),
    .S(_09725_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_1 _19081_ (.A(net3033),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _19082_ (.A0(net46),
    .A1(net6792),
    .S(_03109_),
    .X(_03114_));
 sky130_fd_sc_hd__clkbuf_1 _19083_ (.A(net2056),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _19084_ (.A0(net2182),
    .A1(net6792),
    .S(_09725_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _19085_ (.A(net6794),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _19086_ (.A0(net7496),
    .A1(net5863),
    .S(_03109_),
    .X(_03116_));
 sky130_fd_sc_hd__clkbuf_1 _19087_ (.A(net3042),
    .X(_00755_));
 sky130_fd_sc_hd__and3_1 _19088_ (.A(net7681),
    .B(net5981),
    .C(net4102),
    .X(_03117_));
 sky130_fd_sc_hd__nand2_1 _19089_ (.A(net4095),
    .B(net3970),
    .Y(_03118_));
 sky130_fd_sc_hd__nor2_1 _19090_ (.A(_09733_),
    .B(net4096),
    .Y(_03119_));
 sky130_fd_sc_hd__and4_1 _19091_ (.A(net4092),
    .B(net4138),
    .C(_04657_),
    .D(net4127),
    .X(_03120_));
 sky130_fd_sc_hd__and4b_1 _19092_ (.A_N(net3996),
    .B(_05730_),
    .C(net4097),
    .D(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__buf_4 _19093_ (.A(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__buf_6 _19094_ (.A(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__and2_1 _19095_ (.A(net3623),
    .B(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_4 _19096_ (.A(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__nand2_4 _19097_ (.A(net3623),
    .B(_03123_),
    .Y(_03126_));
 sky130_fd_sc_hd__or2_1 _19098_ (.A(net3367),
    .B(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_4 _19099_ (.A(_09721_),
    .X(_03128_));
 sky130_fd_sc_hd__o211a_1 _19100_ (.A1(net5755),
    .A2(_03125_),
    .B1(net2629),
    .C1(_03128_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _19101_ (.A(net3333),
    .B(_03126_),
    .X(_03129_));
 sky130_fd_sc_hd__o211a_1 _19102_ (.A1(net4309),
    .A2(_03125_),
    .B1(net3036),
    .C1(_03128_),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _19103_ (.A(net2709),
    .B(_03126_),
    .X(_03130_));
 sky130_fd_sc_hd__o211a_1 _19104_ (.A1(net4315),
    .A2(_03125_),
    .B1(net2710),
    .C1(_03128_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _19105_ (.A(net889),
    .B(_03126_),
    .X(_03131_));
 sky130_fd_sc_hd__o211a_1 _19106_ (.A1(net4347),
    .A2(_03125_),
    .B1(net890),
    .C1(_03128_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _19107_ (.A(net5570),
    .B(_03126_),
    .X(_03132_));
 sky130_fd_sc_hd__o211a_1 _19108_ (.A1(net2185),
    .A2(_03125_),
    .B1(net5571),
    .C1(_03128_),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _19109_ (.A(net5526),
    .B(_03126_),
    .X(_03133_));
 sky130_fd_sc_hd__o211a_1 _19110_ (.A1(net1817),
    .A2(_03125_),
    .B1(net5527),
    .C1(_03128_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _19111_ (.A(net5540),
    .B(_03126_),
    .X(_03134_));
 sky130_fd_sc_hd__o211a_1 _19112_ (.A1(net2038),
    .A2(_03125_),
    .B1(net5541),
    .C1(_03128_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _19113_ (.A(net1061),
    .B(_03126_),
    .X(_03135_));
 sky130_fd_sc_hd__o211a_1 _19114_ (.A1(net4324),
    .A2(_03125_),
    .B1(net1062),
    .C1(_03128_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _19115_ (.A(net1076),
    .B(_03126_),
    .X(_03136_));
 sky130_fd_sc_hd__o211a_1 _19116_ (.A1(net4306),
    .A2(_03125_),
    .B1(net1077),
    .C1(_03128_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _19117_ (.A(net5535),
    .B(_03126_),
    .X(_03137_));
 sky130_fd_sc_hd__o211a_1 _19118_ (.A1(net1803),
    .A2(_03125_),
    .B1(net5536),
    .C1(_03128_),
    .X(_00765_));
 sky130_fd_sc_hd__inv_2 _19119_ (.A(net3374),
    .Y(_03138_));
 sky130_fd_sc_hd__nand4b_4 _19120_ (.A_N(net3996),
    .B(_05730_),
    .C(net4097),
    .D(_03120_),
    .Y(_03139_));
 sky130_fd_sc_hd__buf_4 _19121_ (.A(_03122_),
    .X(_03140_));
 sky130_fd_sc_hd__clkbuf_4 _19122_ (.A(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__a21o_1 _19123_ (.A1(net3374),
    .A2(_03141_),
    .B1(net4450),
    .X(_03142_));
 sky130_fd_sc_hd__o311a_1 _19124_ (.A1(net6816),
    .A2(net3375),
    .A3(_03139_),
    .B1(net4451),
    .C1(_08093_),
    .X(_00766_));
 sky130_fd_sc_hd__and2_1 _19125_ (.A(net886),
    .B(_03140_),
    .X(_03143_));
 sky130_fd_sc_hd__clkbuf_2 _19126_ (.A(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_4 _19127_ (.A(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__nand2_2 _19128_ (.A(net886),
    .B(_03140_),
    .Y(_03146_));
 sky130_fd_sc_hd__buf_2 _19129_ (.A(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__or2_1 _19130_ (.A(net1289),
    .B(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__clkbuf_4 _19131_ (.A(_09721_),
    .X(_03149_));
 sky130_fd_sc_hd__o211a_1 _19132_ (.A1(net4354),
    .A2(_03145_),
    .B1(net1290),
    .C1(_03149_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _19133_ (.A(net1176),
    .B(_03147_),
    .X(_03150_));
 sky130_fd_sc_hd__o211a_1 _19134_ (.A1(net4369),
    .A2(_03145_),
    .B1(net1177),
    .C1(_03149_),
    .X(_00768_));
 sky130_fd_sc_hd__or2_1 _19135_ (.A(net1203),
    .B(_03147_),
    .X(_03151_));
 sky130_fd_sc_hd__o211a_1 _19136_ (.A1(net4420),
    .A2(_03145_),
    .B1(net1204),
    .C1(_03149_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _19137_ (.A(net1238),
    .B(_03147_),
    .X(_03152_));
 sky130_fd_sc_hd__o211a_1 _19138_ (.A1(net4431),
    .A2(_03145_),
    .B1(net1239),
    .C1(_03149_),
    .X(_00770_));
 sky130_fd_sc_hd__or2_1 _19139_ (.A(net1133),
    .B(_03147_),
    .X(_03153_));
 sky130_fd_sc_hd__o211a_1 _19140_ (.A1(net5505),
    .A2(_03145_),
    .B1(net1134),
    .C1(_03149_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _19141_ (.A(net1637),
    .B(_03147_),
    .X(_03154_));
 sky130_fd_sc_hd__o211a_1 _19142_ (.A1(net5432),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03149_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _19143_ (.A(net5613),
    .B(_03147_),
    .X(_03155_));
 sky130_fd_sc_hd__o211a_1 _19144_ (.A1(net2587),
    .A2(_03145_),
    .B1(net5614),
    .C1(_03149_),
    .X(_00773_));
 sky130_fd_sc_hd__or2_1 _19145_ (.A(net957),
    .B(_03147_),
    .X(_03156_));
 sky130_fd_sc_hd__o211a_1 _19146_ (.A1(net4366),
    .A2(_03145_),
    .B1(net958),
    .C1(_03149_),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _19147_ (.A(net1830),
    .B(_03147_),
    .X(_03157_));
 sky130_fd_sc_hd__o211a_1 _19148_ (.A1(net4393),
    .A2(_03145_),
    .B1(net1831),
    .C1(_03149_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _19149_ (.A(net2066),
    .B(_03147_),
    .X(_03158_));
 sky130_fd_sc_hd__o211a_1 _19150_ (.A1(net4384),
    .A2(_03145_),
    .B1(net2067),
    .C1(_03149_),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _19151_ (.A(net836),
    .B(_03146_),
    .X(_03159_));
 sky130_fd_sc_hd__clkbuf_4 _19152_ (.A(_09721_),
    .X(_03160_));
 sky130_fd_sc_hd__o211a_1 _19153_ (.A1(net4357),
    .A2(_03144_),
    .B1(net837),
    .C1(_03160_),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _19154_ (.A(net1292),
    .B(_03146_),
    .X(_03161_));
 sky130_fd_sc_hd__o211a_1 _19155_ (.A1(net5468),
    .A2(_03144_),
    .B1(_03161_),
    .C1(_03160_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _19156_ (.A(net1319),
    .B(_03146_),
    .X(_03162_));
 sky130_fd_sc_hd__o211a_1 _19157_ (.A1(net5157),
    .A2(_03144_),
    .B1(_03162_),
    .C1(_03160_),
    .X(_00779_));
 sky130_fd_sc_hd__or2_1 _19158_ (.A(net3002),
    .B(_03146_),
    .X(_03163_));
 sky130_fd_sc_hd__o211a_1 _19159_ (.A1(net5416),
    .A2(_03144_),
    .B1(_03163_),
    .C1(_03160_),
    .X(_00780_));
 sky130_fd_sc_hd__or2_1 _19160_ (.A(net1429),
    .B(_03146_),
    .X(_03164_));
 sky130_fd_sc_hd__o211a_1 _19161_ (.A1(net5420),
    .A2(_03144_),
    .B1(_03164_),
    .C1(_03160_),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _19162_ (.A(net1997),
    .B(_03146_),
    .X(_03165_));
 sky130_fd_sc_hd__o211a_1 _19163_ (.A1(net5392),
    .A2(_03144_),
    .B1(_03165_),
    .C1(_03160_),
    .X(_00782_));
 sky130_fd_sc_hd__and2_1 _19164_ (.A(net3842),
    .B(_03140_),
    .X(_03166_));
 sky130_fd_sc_hd__buf_2 _19165_ (.A(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__buf_4 _19166_ (.A(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__nand2_2 _19167_ (.A(net3842),
    .B(_03123_),
    .Y(_03169_));
 sky130_fd_sc_hd__clkbuf_4 _19168_ (.A(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__or2_1 _19169_ (.A(net6305),
    .B(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__o211a_1 _19170_ (.A1(net5093),
    .A2(_03168_),
    .B1(_03171_),
    .C1(_03160_),
    .X(_00783_));
 sky130_fd_sc_hd__or2_1 _19171_ (.A(net6285),
    .B(_03170_),
    .X(_03172_));
 sky130_fd_sc_hd__o211a_1 _19172_ (.A1(net5053),
    .A2(_03168_),
    .B1(_03172_),
    .C1(_03160_),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _19173_ (.A(net6253),
    .B(_03170_),
    .X(_03173_));
 sky130_fd_sc_hd__o211a_1 _19174_ (.A1(net5236),
    .A2(_03168_),
    .B1(_03173_),
    .C1(_03160_),
    .X(_00785_));
 sky130_fd_sc_hd__or2_1 _19175_ (.A(net6263),
    .B(_03170_),
    .X(_03174_));
 sky130_fd_sc_hd__o211a_1 _19176_ (.A1(net5005),
    .A2(_03168_),
    .B1(_03174_),
    .C1(_03160_),
    .X(_00786_));
 sky130_fd_sc_hd__or2_1 _19177_ (.A(net6448),
    .B(_03170_),
    .X(_03175_));
 sky130_fd_sc_hd__buf_4 _19178_ (.A(_09721_),
    .X(_03176_));
 sky130_fd_sc_hd__o211a_1 _19179_ (.A1(net5081),
    .A2(_03168_),
    .B1(_03175_),
    .C1(_03176_),
    .X(_00787_));
 sky130_fd_sc_hd__or2_1 _19180_ (.A(net6367),
    .B(_03170_),
    .X(_03177_));
 sky130_fd_sc_hd__o211a_1 _19181_ (.A1(net5185),
    .A2(_03168_),
    .B1(_03177_),
    .C1(_03176_),
    .X(_00788_));
 sky130_fd_sc_hd__or2_1 _19182_ (.A(net6297),
    .B(_03170_),
    .X(_03178_));
 sky130_fd_sc_hd__o211a_1 _19183_ (.A1(net5364),
    .A2(_03168_),
    .B1(_03178_),
    .C1(_03176_),
    .X(_00789_));
 sky130_fd_sc_hd__or2_1 _19184_ (.A(net6542),
    .B(_03170_),
    .X(_03179_));
 sky130_fd_sc_hd__o211a_1 _19185_ (.A1(net5256),
    .A2(_03168_),
    .B1(_03179_),
    .C1(_03176_),
    .X(_00790_));
 sky130_fd_sc_hd__or2_1 _19186_ (.A(net6281),
    .B(_03170_),
    .X(_03180_));
 sky130_fd_sc_hd__o211a_1 _19187_ (.A1(net5240),
    .A2(_03168_),
    .B1(_03180_),
    .C1(_03176_),
    .X(_00791_));
 sky130_fd_sc_hd__or2_1 _19188_ (.A(net6566),
    .B(_03170_),
    .X(_03181_));
 sky130_fd_sc_hd__o211a_1 _19189_ (.A1(net5324),
    .A2(_03168_),
    .B1(_03181_),
    .C1(_03176_),
    .X(_00792_));
 sky130_fd_sc_hd__buf_4 _19190_ (.A(_03167_),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_4 _19191_ (.A(_03169_),
    .X(_03183_));
 sky130_fd_sc_hd__or2_1 _19192_ (.A(net6315),
    .B(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__o211a_1 _19193_ (.A1(net5212),
    .A2(_03182_),
    .B1(_03184_),
    .C1(_03176_),
    .X(_00793_));
 sky130_fd_sc_hd__or2_1 _19194_ (.A(net1923),
    .B(_03183_),
    .X(_03185_));
 sky130_fd_sc_hd__o211a_1 _19195_ (.A1(net5292),
    .A2(_03182_),
    .B1(_03185_),
    .C1(_03176_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _19196_ (.A(net6434),
    .B(_03183_),
    .X(_03186_));
 sky130_fd_sc_hd__o211a_1 _19197_ (.A1(net5244),
    .A2(_03182_),
    .B1(_03186_),
    .C1(_03176_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _19198_ (.A(net6388),
    .B(_03183_),
    .X(_03187_));
 sky130_fd_sc_hd__o211a_1 _19199_ (.A1(net5372),
    .A2(_03182_),
    .B1(_03187_),
    .C1(_03176_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _19200_ (.A(net6697),
    .B(_03183_),
    .X(_03188_));
 sky130_fd_sc_hd__buf_4 _19201_ (.A(_09721_),
    .X(_03189_));
 sky130_fd_sc_hd__o211a_1 _19202_ (.A1(net5121),
    .A2(_03182_),
    .B1(_03188_),
    .C1(_03189_),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _19203_ (.A(net6520),
    .B(_03183_),
    .X(_03190_));
 sky130_fd_sc_hd__o211a_1 _19204_ (.A1(net5232),
    .A2(_03182_),
    .B1(_03190_),
    .C1(_03189_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _19205_ (.A(net6301),
    .B(_03183_),
    .X(_03191_));
 sky130_fd_sc_hd__o211a_1 _19206_ (.A1(net5065),
    .A2(_03182_),
    .B1(_03191_),
    .C1(_03189_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _19207_ (.A(net6862),
    .B(_03183_),
    .X(_03192_));
 sky130_fd_sc_hd__o211a_1 _19208_ (.A1(net5149),
    .A2(_03182_),
    .B1(_03192_),
    .C1(_03189_),
    .X(_00800_));
 sky130_fd_sc_hd__or2_1 _19209_ (.A(net6727),
    .B(_03183_),
    .X(_03193_));
 sky130_fd_sc_hd__o211a_1 _19210_ (.A1(net5165),
    .A2(_03182_),
    .B1(_03193_),
    .C1(_03189_),
    .X(_00801_));
 sky130_fd_sc_hd__or2_1 _19211_ (.A(net6516),
    .B(_03183_),
    .X(_03194_));
 sky130_fd_sc_hd__o211a_1 _19212_ (.A1(net5220),
    .A2(_03182_),
    .B1(_03194_),
    .C1(_03189_),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _19213_ (.A(net1331),
    .B(_03169_),
    .X(_03195_));
 sky130_fd_sc_hd__o211a_1 _19214_ (.A1(net5336),
    .A2(_03167_),
    .B1(_03195_),
    .C1(_03189_),
    .X(_00803_));
 sky130_fd_sc_hd__or2_1 _19215_ (.A(net1649),
    .B(_03169_),
    .X(_03196_));
 sky130_fd_sc_hd__o211a_1 _19216_ (.A1(net5348),
    .A2(_03167_),
    .B1(_03196_),
    .C1(_03189_),
    .X(_00804_));
 sky130_fd_sc_hd__or2_1 _19217_ (.A(net1432),
    .B(_03169_),
    .X(_03197_));
 sky130_fd_sc_hd__o211a_1 _19218_ (.A1(net5436),
    .A2(_03167_),
    .B1(_03197_),
    .C1(_03189_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _19219_ (.A(net6321),
    .B(_03169_),
    .X(_03198_));
 sky130_fd_sc_hd__o211a_1 _19220_ (.A1(net5444),
    .A2(_03167_),
    .B1(_03198_),
    .C1(_03189_),
    .X(_00806_));
 sky130_fd_sc_hd__and2_1 _19221_ (.A(net1030),
    .B(_03140_),
    .X(_03199_));
 sky130_fd_sc_hd__buf_2 _19222_ (.A(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_4 _19223_ (.A(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__nand2_2 _19224_ (.A(net1030),
    .B(_03123_),
    .Y(_03202_));
 sky130_fd_sc_hd__buf_2 _19225_ (.A(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__or2_1 _19226_ (.A(net6474),
    .B(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__clkbuf_4 _19227_ (.A(_08092_),
    .X(_03205_));
 sky130_fd_sc_hd__clkbuf_4 _19228_ (.A(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__o211a_1 _19229_ (.A1(net5264),
    .A2(_03201_),
    .B1(_03204_),
    .C1(_03206_),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _19230_ (.A(net6313),
    .B(_03203_),
    .X(_03207_));
 sky130_fd_sc_hd__o211a_1 _19231_ (.A1(net5332),
    .A2(_03201_),
    .B1(_03207_),
    .C1(_03206_),
    .X(_00808_));
 sky130_fd_sc_hd__or2_1 _19232_ (.A(net6341),
    .B(_03203_),
    .X(_03208_));
 sky130_fd_sc_hd__o211a_1 _19233_ (.A1(net5125),
    .A2(_03201_),
    .B1(_03208_),
    .C1(_03206_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _19234_ (.A(net6504),
    .B(_03203_),
    .X(_03209_));
 sky130_fd_sc_hd__o211a_1 _19235_ (.A1(net5352),
    .A2(_03201_),
    .B1(_03209_),
    .C1(_03206_),
    .X(_00810_));
 sky130_fd_sc_hd__or2_1 _19236_ (.A(net6440),
    .B(_03203_),
    .X(_03210_));
 sky130_fd_sc_hd__o211a_1 _19237_ (.A1(net5097),
    .A2(_03201_),
    .B1(_03210_),
    .C1(_03206_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _19238_ (.A(net6419),
    .B(_03203_),
    .X(_03211_));
 sky130_fd_sc_hd__o211a_1 _19239_ (.A1(net5141),
    .A2(_03201_),
    .B1(_03211_),
    .C1(_03206_),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _19240_ (.A(net6599),
    .B(_03203_),
    .X(_03212_));
 sky130_fd_sc_hd__o211a_1 _19241_ (.A1(net5228),
    .A2(_03201_),
    .B1(_03212_),
    .C1(_03206_),
    .X(_00813_));
 sky130_fd_sc_hd__or2_1 _19242_ (.A(net6532),
    .B(_03203_),
    .X(_03213_));
 sky130_fd_sc_hd__o211a_1 _19243_ (.A1(net5029),
    .A2(_03201_),
    .B1(_03213_),
    .C1(_03206_),
    .X(_00814_));
 sky130_fd_sc_hd__or2_1 _19244_ (.A(net1552),
    .B(_03203_),
    .X(_03214_));
 sky130_fd_sc_hd__o211a_1 _19245_ (.A1(net5077),
    .A2(_03201_),
    .B1(_03214_),
    .C1(_03206_),
    .X(_00815_));
 sky130_fd_sc_hd__or2_1 _19246_ (.A(net6351),
    .B(_03203_),
    .X(_03215_));
 sky130_fd_sc_hd__o211a_1 _19247_ (.A1(net5061),
    .A2(_03201_),
    .B1(_03215_),
    .C1(_03206_),
    .X(_00816_));
 sky130_fd_sc_hd__clkbuf_4 _19248_ (.A(_03200_),
    .X(_03216_));
 sky130_fd_sc_hd__buf_2 _19249_ (.A(_03202_),
    .X(_03217_));
 sky130_fd_sc_hd__or2_1 _19250_ (.A(net6417),
    .B(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_4 _19251_ (.A(_03205_),
    .X(_03219_));
 sky130_fd_sc_hd__o211a_1 _19252_ (.A1(net5388),
    .A2(_03216_),
    .B1(_03218_),
    .C1(_03219_),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _19253_ (.A(net6325),
    .B(_03217_),
    .X(_03220_));
 sky130_fd_sc_hd__o211a_1 _19254_ (.A1(net5424),
    .A2(_03216_),
    .B1(_03220_),
    .C1(_03219_),
    .X(_00818_));
 sky130_fd_sc_hd__or2_1 _19255_ (.A(net6370),
    .B(_03217_),
    .X(_03221_));
 sky130_fd_sc_hd__o211a_1 _19256_ (.A1(net5145),
    .A2(_03216_),
    .B1(_03221_),
    .C1(_03219_),
    .X(_00819_));
 sky130_fd_sc_hd__or2_1 _19257_ (.A(net6484),
    .B(_03217_),
    .X(_03222_));
 sky130_fd_sc_hd__o211a_1 _19258_ (.A1(net5169),
    .A2(_03216_),
    .B1(_03222_),
    .C1(_03219_),
    .X(_00820_));
 sky130_fd_sc_hd__or2_1 _19259_ (.A(net986),
    .B(_03217_),
    .X(_03223_));
 sky130_fd_sc_hd__o211a_1 _19260_ (.A1(net8135),
    .A2(_03216_),
    .B1(net987),
    .C1(_03219_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _19261_ (.A(net6422),
    .B(_03217_),
    .X(_03224_));
 sky130_fd_sc_hd__o211a_1 _19262_ (.A1(net5320),
    .A2(_03216_),
    .B1(_03224_),
    .C1(_03219_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _19263_ (.A(net6347),
    .B(_03217_),
    .X(_03225_));
 sky130_fd_sc_hd__o211a_1 _19264_ (.A1(net5284),
    .A2(_03216_),
    .B1(_03225_),
    .C1(_03219_),
    .X(_00823_));
 sky130_fd_sc_hd__or2_1 _19265_ (.A(net6623),
    .B(_03217_),
    .X(_03226_));
 sky130_fd_sc_hd__o211a_1 _19266_ (.A1(net5109),
    .A2(_03216_),
    .B1(_03226_),
    .C1(_03219_),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _19267_ (.A(net6629),
    .B(_03217_),
    .X(_03227_));
 sky130_fd_sc_hd__o211a_1 _19268_ (.A1(net5308),
    .A2(_03216_),
    .B1(_03227_),
    .C1(_03219_),
    .X(_00825_));
 sky130_fd_sc_hd__or2_1 _19269_ (.A(net6562),
    .B(_03217_),
    .X(_03228_));
 sky130_fd_sc_hd__o211a_1 _19270_ (.A1(net5412),
    .A2(_03216_),
    .B1(_03228_),
    .C1(_03219_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _19271_ (.A(net2075),
    .B(_03202_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_4 _19272_ (.A(_03205_),
    .X(_03230_));
 sky130_fd_sc_hd__o211a_1 _19273_ (.A1(net5057),
    .A2(_03200_),
    .B1(_03229_),
    .C1(_03230_),
    .X(_00827_));
 sky130_fd_sc_hd__or2_1 _19274_ (.A(net2414),
    .B(_03202_),
    .X(_03231_));
 sky130_fd_sc_hd__o211a_1 _19275_ (.A1(net5037),
    .A2(_03200_),
    .B1(_03231_),
    .C1(_03230_),
    .X(_00828_));
 sky130_fd_sc_hd__or2_1 _19276_ (.A(net6132),
    .B(_03202_),
    .X(_03232_));
 sky130_fd_sc_hd__o211a_1 _19277_ (.A1(net5368),
    .A2(_03200_),
    .B1(_03232_),
    .C1(_03230_),
    .X(_00829_));
 sky130_fd_sc_hd__or2_1 _19278_ (.A(net1523),
    .B(_03202_),
    .X(_03233_));
 sky130_fd_sc_hd__o211a_1 _19279_ (.A1(net5089),
    .A2(_03200_),
    .B1(_03233_),
    .C1(_03230_),
    .X(_00830_));
 sky130_fd_sc_hd__and2_1 _19280_ (.A(net4842),
    .B(_03140_),
    .X(_03234_));
 sky130_fd_sc_hd__buf_2 _19281_ (.A(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_4 _19282_ (.A(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__nand2_4 _19283_ (.A(net4842),
    .B(_03123_),
    .Y(_03237_));
 sky130_fd_sc_hd__buf_2 _19284_ (.A(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__or2_1 _19285_ (.A(net1286),
    .B(_03238_),
    .X(_03239_));
 sky130_fd_sc_hd__o211a_1 _19286_ (.A1(net5129),
    .A2(_03236_),
    .B1(_03239_),
    .C1(_03230_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _19287_ (.A(net597),
    .B(_03238_),
    .X(_03240_));
 sky130_fd_sc_hd__o211a_1 _19288_ (.A1(net8118),
    .A2(_03236_),
    .B1(net598),
    .C1(_03230_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _19289_ (.A(net1422),
    .B(_03238_),
    .X(_03241_));
 sky130_fd_sc_hd__o211a_1 _19290_ (.A1(net5161),
    .A2(_03236_),
    .B1(_03241_),
    .C1(_03230_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_1 _19291_ (.A(net1281),
    .B(_03238_),
    .X(_03242_));
 sky130_fd_sc_hd__o211a_1 _19292_ (.A1(net5268),
    .A2(_03236_),
    .B1(_03242_),
    .C1(_03230_),
    .X(_00834_));
 sky130_fd_sc_hd__or2_1 _19293_ (.A(net6299),
    .B(_03238_),
    .X(_03243_));
 sky130_fd_sc_hd__o211a_1 _19294_ (.A1(net5201),
    .A2(_03236_),
    .B1(_03243_),
    .C1(_03230_),
    .X(_00835_));
 sky130_fd_sc_hd__or2_1 _19295_ (.A(net6390),
    .B(_03238_),
    .X(_03244_));
 sky130_fd_sc_hd__o211a_1 _19296_ (.A1(net5216),
    .A2(_03236_),
    .B1(_03244_),
    .C1(_03230_),
    .X(_00836_));
 sky130_fd_sc_hd__or2_1 _19297_ (.A(net1538),
    .B(_03238_),
    .X(_03245_));
 sky130_fd_sc_hd__buf_4 _19298_ (.A(_03205_),
    .X(_03246_));
 sky130_fd_sc_hd__o211a_1 _19299_ (.A1(net5117),
    .A2(_03236_),
    .B1(_03245_),
    .C1(_03246_),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _19300_ (.A(net1631),
    .B(_03238_),
    .X(_03247_));
 sky130_fd_sc_hd__o211a_1 _19301_ (.A1(net5296),
    .A2(_03236_),
    .B1(_03247_),
    .C1(_03246_),
    .X(_00838_));
 sky130_fd_sc_hd__or2_1 _19302_ (.A(net1508),
    .B(_03238_),
    .X(_03248_));
 sky130_fd_sc_hd__o211a_1 _19303_ (.A1(net5073),
    .A2(_03236_),
    .B1(_03248_),
    .C1(_03246_),
    .X(_00839_));
 sky130_fd_sc_hd__or2_1 _19304_ (.A(net1514),
    .B(_03238_),
    .X(_03249_));
 sky130_fd_sc_hd__o211a_1 _19305_ (.A1(net5137),
    .A2(_03236_),
    .B1(_03249_),
    .C1(_03246_),
    .X(_00840_));
 sky130_fd_sc_hd__buf_4 _19306_ (.A(_03235_),
    .X(_03250_));
 sky130_fd_sc_hd__clkbuf_4 _19307_ (.A(_03237_),
    .X(_03251_));
 sky130_fd_sc_hd__or2_1 _19308_ (.A(net1435),
    .B(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__o211a_1 _19309_ (.A1(net5260),
    .A2(_03250_),
    .B1(_03252_),
    .C1(_03246_),
    .X(_00841_));
 sky130_fd_sc_hd__or2_1 _19310_ (.A(net1859),
    .B(_03251_),
    .X(_03253_));
 sky130_fd_sc_hd__o211a_1 _19311_ (.A1(net5085),
    .A2(_03250_),
    .B1(_03253_),
    .C1(_03246_),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _19312_ (.A(net1456),
    .B(_03251_),
    .X(_03254_));
 sky130_fd_sc_hd__o211a_1 _19313_ (.A1(net5300),
    .A2(_03250_),
    .B1(_03254_),
    .C1(_03246_),
    .X(_00843_));
 sky130_fd_sc_hd__or2_1 _19314_ (.A(net1677),
    .B(_03251_),
    .X(_03255_));
 sky130_fd_sc_hd__o211a_1 _19315_ (.A1(net5316),
    .A2(_03250_),
    .B1(_03255_),
    .C1(_03246_),
    .X(_00844_));
 sky130_fd_sc_hd__or2_1 _19316_ (.A(net1380),
    .B(_03251_),
    .X(_03256_));
 sky130_fd_sc_hd__o211a_1 _19317_ (.A1(net5456),
    .A2(_03250_),
    .B1(_03256_),
    .C1(_03246_),
    .X(_00845_));
 sky130_fd_sc_hd__or2_1 _19318_ (.A(net1444),
    .B(_03251_),
    .X(_03257_));
 sky130_fd_sc_hd__o211a_1 _19319_ (.A1(net5177),
    .A2(_03250_),
    .B1(_03257_),
    .C1(_03246_),
    .X(_00846_));
 sky130_fd_sc_hd__or2_1 _19320_ (.A(net1371),
    .B(_03251_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_4 _19321_ (.A(_03205_),
    .X(_03259_));
 sky130_fd_sc_hd__o211a_1 _19322_ (.A1(net5181),
    .A2(_03250_),
    .B1(_03258_),
    .C1(_03259_),
    .X(_00847_));
 sky130_fd_sc_hd__or2_1 _19323_ (.A(net1718),
    .B(_03251_),
    .X(_03260_));
 sky130_fd_sc_hd__o211a_1 _19324_ (.A1(net5276),
    .A2(_03250_),
    .B1(_03260_),
    .C1(_03259_),
    .X(_00848_));
 sky130_fd_sc_hd__or2_1 _19325_ (.A(net1602),
    .B(_03251_),
    .X(_03261_));
 sky130_fd_sc_hd__o211a_1 _19326_ (.A1(net5133),
    .A2(_03250_),
    .B1(_03261_),
    .C1(_03259_),
    .X(_00849_));
 sky130_fd_sc_hd__or2_1 _19327_ (.A(net839),
    .B(_03251_),
    .X(_03262_));
 sky130_fd_sc_hd__o211a_1 _19328_ (.A1(net8116),
    .A2(_03250_),
    .B1(net840),
    .C1(_03259_),
    .X(_00850_));
 sky130_fd_sc_hd__or2_1 _19329_ (.A(net1343),
    .B(_03237_),
    .X(_03263_));
 sky130_fd_sc_hd__o211a_1 _19330_ (.A1(net5013),
    .A2(_03235_),
    .B1(_03263_),
    .C1(_03259_),
    .X(_00851_));
 sky130_fd_sc_hd__or2_1 _19331_ (.A(net1505),
    .B(_03237_),
    .X(_03264_));
 sky130_fd_sc_hd__o211a_1 _19332_ (.A1(net5069),
    .A2(_03235_),
    .B1(_03264_),
    .C1(_03259_),
    .X(_00852_));
 sky130_fd_sc_hd__or2_1 _19333_ (.A(net1599),
    .B(_03237_),
    .X(_03265_));
 sky130_fd_sc_hd__o211a_1 _19334_ (.A1(net5304),
    .A2(_03235_),
    .B1(_03265_),
    .C1(_03259_),
    .X(_00853_));
 sky130_fd_sc_hd__or2_1 _19335_ (.A(net6331),
    .B(_03237_),
    .X(_03266_));
 sky130_fd_sc_hd__o211a_1 _19336_ (.A1(net5344),
    .A2(_03235_),
    .B1(_03266_),
    .C1(_03259_),
    .X(_00854_));
 sky130_fd_sc_hd__and2_1 _19337_ (.A(net1020),
    .B(_03140_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_2 _19338_ (.A(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__clkbuf_4 _19339_ (.A(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__nand2_2 _19340_ (.A(net1020),
    .B(_03140_),
    .Y(_03270_));
 sky130_fd_sc_hd__clkbuf_4 _19341_ (.A(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__or2_1 _19342_ (.A(net6275),
    .B(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__o211a_1 _19343_ (.A1(net5017),
    .A2(_03269_),
    .B1(_03272_),
    .C1(_03259_),
    .X(_00855_));
 sky130_fd_sc_hd__or2_1 _19344_ (.A(net6552),
    .B(_03271_),
    .X(_03273_));
 sky130_fd_sc_hd__o211a_1 _19345_ (.A1(net5041),
    .A2(_03269_),
    .B1(_03273_),
    .C1(_03259_),
    .X(_00856_));
 sky130_fd_sc_hd__or2_1 _19346_ (.A(net6374),
    .B(_03271_),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_4 _19347_ (.A(_03205_),
    .X(_03275_));
 sky130_fd_sc_hd__o211a_1 _19348_ (.A1(net5193),
    .A2(_03269_),
    .B1(_03274_),
    .C1(_03275_),
    .X(_00857_));
 sky130_fd_sc_hd__or2_1 _19349_ (.A(net6409),
    .B(_03271_),
    .X(_03276_));
 sky130_fd_sc_hd__o211a_1 _19350_ (.A1(net4992),
    .A2(_03269_),
    .B1(_03276_),
    .C1(_03275_),
    .X(_00858_));
 sky130_fd_sc_hd__or2_1 _19351_ (.A(net6510),
    .B(_03271_),
    .X(_03277_));
 sky130_fd_sc_hd__o211a_1 _19352_ (.A1(net5113),
    .A2(_03269_),
    .B1(_03277_),
    .C1(_03275_),
    .X(_00859_));
 sky130_fd_sc_hd__or2_1 _19353_ (.A(net6450),
    .B(_03271_),
    .X(_03278_));
 sky130_fd_sc_hd__o211a_1 _19354_ (.A1(net5360),
    .A2(_03269_),
    .B1(_03278_),
    .C1(_03275_),
    .X(_00860_));
 sky130_fd_sc_hd__or2_1 _19355_ (.A(net6283),
    .B(_03271_),
    .X(_03279_));
 sky130_fd_sc_hd__o211a_1 _19356_ (.A1(net5396),
    .A2(_03269_),
    .B1(_03279_),
    .C1(_03275_),
    .X(_00861_));
 sky130_fd_sc_hd__or2_1 _19357_ (.A(net6378),
    .B(_03271_),
    .X(_03280_));
 sky130_fd_sc_hd__o211a_1 _19358_ (.A1(net5312),
    .A2(_03269_),
    .B1(_03280_),
    .C1(_03275_),
    .X(_00862_));
 sky130_fd_sc_hd__or2_1 _19359_ (.A(net6265),
    .B(_03271_),
    .X(_03281_));
 sky130_fd_sc_hd__o211a_1 _19360_ (.A1(net5105),
    .A2(_03269_),
    .B1(_03281_),
    .C1(_03275_),
    .X(_00863_));
 sky130_fd_sc_hd__or2_1 _19361_ (.A(net6309),
    .B(_03271_),
    .X(_03282_));
 sky130_fd_sc_hd__o211a_1 _19362_ (.A1(net5288),
    .A2(_03269_),
    .B1(_03282_),
    .C1(_03275_),
    .X(_00864_));
 sky130_fd_sc_hd__buf_4 _19363_ (.A(_03268_),
    .X(_03283_));
 sky130_fd_sc_hd__clkbuf_4 _19364_ (.A(_03270_),
    .X(_03284_));
 sky130_fd_sc_hd__or2_1 _19365_ (.A(net1474),
    .B(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_1 _19366_ (.A1(net5021),
    .A2(_03283_),
    .B1(_03285_),
    .C1(_03275_),
    .X(_00865_));
 sky130_fd_sc_hd__or2_1 _19367_ (.A(net1785),
    .B(_03284_),
    .X(_03286_));
 sky130_fd_sc_hd__o211a_1 _19368_ (.A1(net5009),
    .A2(_03283_),
    .B1(_03286_),
    .C1(_03275_),
    .X(_00866_));
 sky130_fd_sc_hd__or2_1 _19369_ (.A(net6257),
    .B(_03284_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_4 _19370_ (.A(_03205_),
    .X(_03288_));
 sky130_fd_sc_hd__o211a_1 _19371_ (.A1(net5025),
    .A2(_03283_),
    .B1(_03287_),
    .C1(_03288_),
    .X(_00867_));
 sky130_fd_sc_hd__or2_1 _19372_ (.A(net6470),
    .B(_03284_),
    .X(_03289_));
 sky130_fd_sc_hd__o211a_1 _19373_ (.A1(net5001),
    .A2(_03283_),
    .B1(_03289_),
    .C1(_03288_),
    .X(_00868_));
 sky130_fd_sc_hd__or2_1 _19374_ (.A(net6372),
    .B(_03284_),
    .X(_03290_));
 sky130_fd_sc_hd__o211a_1 _19375_ (.A1(net5101),
    .A2(_03283_),
    .B1(_03290_),
    .C1(_03288_),
    .X(_00869_));
 sky130_fd_sc_hd__or2_1 _19376_ (.A(net6570),
    .B(_03284_),
    .X(_03291_));
 sky130_fd_sc_hd__o211a_1 _19377_ (.A1(net5224),
    .A2(_03283_),
    .B1(_03291_),
    .C1(_03288_),
    .X(_00870_));
 sky130_fd_sc_hd__or2_1 _19378_ (.A(net6496),
    .B(_03284_),
    .X(_03292_));
 sky130_fd_sc_hd__o211a_1 _19379_ (.A1(net5153),
    .A2(_03283_),
    .B1(_03292_),
    .C1(_03288_),
    .X(_00871_));
 sky130_fd_sc_hd__or2_1 _19380_ (.A(net6677),
    .B(_03284_),
    .X(_03293_));
 sky130_fd_sc_hd__o211a_1 _19381_ (.A1(net5173),
    .A2(_03283_),
    .B1(_03293_),
    .C1(_03288_),
    .X(_00872_));
 sky130_fd_sc_hd__or2_1 _19382_ (.A(net6317),
    .B(_03284_),
    .X(_03294_));
 sky130_fd_sc_hd__o211a_1 _19383_ (.A1(net5189),
    .A2(_03283_),
    .B1(_03294_),
    .C1(_03288_),
    .X(_00873_));
 sky130_fd_sc_hd__or2_1 _19384_ (.A(net6683),
    .B(_03284_),
    .X(_03295_));
 sky130_fd_sc_hd__o211a_1 _19385_ (.A1(net5197),
    .A2(_03283_),
    .B1(_03295_),
    .C1(_03288_),
    .X(_00874_));
 sky130_fd_sc_hd__or2_1 _19386_ (.A(net6136),
    .B(_03270_),
    .X(_03296_));
 sky130_fd_sc_hd__o211a_1 _19387_ (.A1(net4988),
    .A2(_03268_),
    .B1(_03296_),
    .C1(_03288_),
    .X(_00875_));
 sky130_fd_sc_hd__or2_1 _19388_ (.A(net6080),
    .B(_03270_),
    .X(_03297_));
 sky130_fd_sc_hd__o211a_1 _19389_ (.A1(net5248),
    .A2(_03268_),
    .B1(_03297_),
    .C1(_03288_),
    .X(_00876_));
 sky130_fd_sc_hd__or2_1 _19390_ (.A(net6180),
    .B(_03270_),
    .X(_03298_));
 sky130_fd_sc_hd__buf_4 _19391_ (.A(_03205_),
    .X(_03299_));
 sky130_fd_sc_hd__o211a_1 _19392_ (.A1(net5272),
    .A2(_03268_),
    .B1(_03298_),
    .C1(_03299_),
    .X(_00877_));
 sky130_fd_sc_hd__or2_1 _19393_ (.A(net1386),
    .B(_03270_),
    .X(_03300_));
 sky130_fd_sc_hd__o211a_1 _19394_ (.A1(net4976),
    .A2(_03268_),
    .B1(_03300_),
    .C1(_03299_),
    .X(_00878_));
 sky130_fd_sc_hd__and2_1 _19395_ (.A(net3217),
    .B(_03123_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_2 _19396_ (.A(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__nand2_2 _19397_ (.A(net3217),
    .B(_03141_),
    .Y(_03303_));
 sky130_fd_sc_hd__or2_1 _19398_ (.A(net2447),
    .B(_03303_),
    .X(_03304_));
 sky130_fd_sc_hd__o211a_1 _19399_ (.A1(net5440),
    .A2(_03302_),
    .B1(_03304_),
    .C1(_03299_),
    .X(_00879_));
 sky130_fd_sc_hd__or2_1 _19400_ (.A(net1643),
    .B(_03303_),
    .X(_03305_));
 sky130_fd_sc_hd__o211a_1 _19401_ (.A1(net5460),
    .A2(_03302_),
    .B1(_03305_),
    .C1(_03299_),
    .X(_00880_));
 sky130_fd_sc_hd__or2_1 _19402_ (.A(net2256),
    .B(_03303_),
    .X(_03306_));
 sky130_fd_sc_hd__o211a_1 _19403_ (.A1(net5484),
    .A2(_03302_),
    .B1(_03306_),
    .C1(_03299_),
    .X(_00881_));
 sky130_fd_sc_hd__or2_1 _19404_ (.A(net5500),
    .B(_03303_),
    .X(_03307_));
 sky130_fd_sc_hd__o211a_1 _19405_ (.A1(net1255),
    .A2(_03302_),
    .B1(net5501),
    .C1(_03299_),
    .X(_00882_));
 sky130_fd_sc_hd__or2_1 _19406_ (.A(net1671),
    .B(_03303_),
    .X(_03308_));
 sky130_fd_sc_hd__o211a_1 _19407_ (.A1(net5518),
    .A2(_03302_),
    .B1(_03308_),
    .C1(_03299_),
    .X(_00883_));
 sky130_fd_sc_hd__or2_1 _19408_ (.A(net2146),
    .B(_03303_),
    .X(_03309_));
 sky130_fd_sc_hd__o211a_1 _19409_ (.A1(net5509),
    .A2(_03302_),
    .B1(_03309_),
    .C1(_03299_),
    .X(_00884_));
 sky130_fd_sc_hd__nand2_2 _19410_ (.A(net3902),
    .B(_03140_),
    .Y(_03310_));
 sky130_fd_sc_hd__and3_1 _19411_ (.A(net1733),
    .B(net3902),
    .C(_03141_),
    .X(_03311_));
 sky130_fd_sc_hd__buf_6 _19412_ (.A(_04459_),
    .X(_03312_));
 sky130_fd_sc_hd__a211o_1 _19413_ (.A1(net5356),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03312_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _19414_ (.A0(net1532),
    .A1(net3569),
    .S(_03310_),
    .X(_03313_));
 sky130_fd_sc_hd__and2_1 _19415_ (.A(_08093_),
    .B(net3570),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_1 _19416_ (.A(net3571),
    .X(_00886_));
 sky130_fd_sc_hd__and3_1 _19417_ (.A(net2321),
    .B(net3902),
    .C(_03141_),
    .X(_03315_));
 sky130_fd_sc_hd__buf_4 _19418_ (.A(_04459_),
    .X(_03316_));
 sky130_fd_sc_hd__a211o_1 _19419_ (.A1(net4964),
    .A2(_03310_),
    .B1(_03315_),
    .C1(_03316_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _19420_ (.A0(net1724),
    .A1(net3670),
    .S(_03310_),
    .X(_03317_));
 sky130_fd_sc_hd__and2_1 _19421_ (.A(_08093_),
    .B(net3671),
    .X(_03318_));
 sky130_fd_sc_hd__clkbuf_1 _19422_ (.A(net3672),
    .X(_00888_));
 sky130_fd_sc_hd__and3_1 _19423_ (.A(net2441),
    .B(net3902),
    .C(_03141_),
    .X(_03319_));
 sky130_fd_sc_hd__a211o_1 _19424_ (.A1(net5049),
    .A2(_03310_),
    .B1(_03319_),
    .C1(_03316_),
    .X(_00889_));
 sky130_fd_sc_hd__clkbuf_4 _19425_ (.A(_08092_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _19426_ (.A0(net2060),
    .A1(net3651),
    .S(_03310_),
    .X(_03321_));
 sky130_fd_sc_hd__and2_1 _19427_ (.A(_03320_),
    .B(net3652),
    .X(_03322_));
 sky130_fd_sc_hd__clkbuf_1 _19428_ (.A(net3653),
    .X(_00890_));
 sky130_fd_sc_hd__nand2_2 _19429_ (.A(net3519),
    .B(_03122_),
    .Y(_03323_));
 sky130_fd_sc_hd__mux2_1 _19430_ (.A0(net1480),
    .A1(net3656),
    .S(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__and2_1 _19431_ (.A(_03320_),
    .B(net3657),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _19432_ (.A(net3658),
    .X(_00891_));
 sky130_fd_sc_hd__and3_1 _19433_ (.A(net1593),
    .B(net3519),
    .C(_03141_),
    .X(_03326_));
 sky130_fd_sc_hd__a211o_1 _19434_ (.A1(net4960),
    .A2(_03323_),
    .B1(_03326_),
    .C1(_03316_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _19435_ (.A0(net1564),
    .A1(net3547),
    .S(_03323_),
    .X(_03327_));
 sky130_fd_sc_hd__and2_1 _19436_ (.A(_03320_),
    .B(net3548),
    .X(_03328_));
 sky130_fd_sc_hd__clkbuf_1 _19437_ (.A(net3549),
    .X(_00893_));
 sky130_fd_sc_hd__and3_1 _19438_ (.A(net1625),
    .B(net3519),
    .C(_03141_),
    .X(_03329_));
 sky130_fd_sc_hd__a211o_1 _19439_ (.A1(net4952),
    .A2(_03323_),
    .B1(_03329_),
    .C1(_03316_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _19440_ (.A0(net2232),
    .A1(net3644),
    .S(_03323_),
    .X(_03330_));
 sky130_fd_sc_hd__and2_1 _19441_ (.A(_03320_),
    .B(net3645),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _19442_ (.A(net3646),
    .X(_00895_));
 sky130_fd_sc_hd__and3_1 _19443_ (.A(net1561),
    .B(net3519),
    .C(_03141_),
    .X(_03332_));
 sky130_fd_sc_hd__a211o_1 _19444_ (.A1(net4956),
    .A2(_03323_),
    .B1(_03332_),
    .C1(_03316_),
    .X(_00896_));
 sky130_fd_sc_hd__and2_1 _19445_ (.A(net3978),
    .B(_03123_),
    .X(_03333_));
 sky130_fd_sc_hd__clkbuf_2 _19446_ (.A(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__nand2_2 _19447_ (.A(net3978),
    .B(_03123_),
    .Y(_03335_));
 sky130_fd_sc_hd__or2_1 _19448_ (.A(net1033),
    .B(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__o211a_1 _19449_ (.A1(net4312),
    .A2(_03334_),
    .B1(net1034),
    .C1(_03299_),
    .X(_00897_));
 sky130_fd_sc_hd__or2_1 _19450_ (.A(net5513),
    .B(_03335_),
    .X(_03337_));
 sky130_fd_sc_hd__o211a_1 _19451_ (.A1(net1658),
    .A2(_03334_),
    .B1(net5514),
    .C1(_03299_),
    .X(_00898_));
 sky130_fd_sc_hd__or2_1 _19452_ (.A(net5562),
    .B(_03335_),
    .X(_03338_));
 sky130_fd_sc_hd__buf_4 _19453_ (.A(_03205_),
    .X(_03339_));
 sky130_fd_sc_hd__o211a_1 _19454_ (.A1(net1851),
    .A2(_03334_),
    .B1(net5563),
    .C1(_03339_),
    .X(_00899_));
 sky130_fd_sc_hd__or2_1 _19455_ (.A(net2098),
    .B(_03335_),
    .X(_03340_));
 sky130_fd_sc_hd__o211a_1 _19456_ (.A1(net4230),
    .A2(_03334_),
    .B1(net1366),
    .C1(_03339_),
    .X(_00900_));
 sky130_fd_sc_hd__or2_1 _19457_ (.A(net1742),
    .B(_03335_),
    .X(_03341_));
 sky130_fd_sc_hd__o211a_1 _19458_ (.A1(net5464),
    .A2(_03334_),
    .B1(_03341_),
    .C1(_03339_),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _19459_ (.A(net2223),
    .B(_03335_),
    .X(_03342_));
 sky130_fd_sc_hd__o211a_1 _19460_ (.A1(net5452),
    .A2(_03334_),
    .B1(_03342_),
    .C1(_03339_),
    .X(_00902_));
 sky130_fd_sc_hd__and4bb_1 _19461_ (.A_N(net3486),
    .B_N(net3906),
    .C(_02947_),
    .D(_02969_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _19462_ (.A(net3907),
    .X(_00903_));
 sky130_fd_sc_hd__or3b_4 _19463_ (.A(net3940),
    .B(net5895),
    .C_N(net3906),
    .X(_03344_));
 sky130_fd_sc_hd__or3_4 _19464_ (.A(_04458_),
    .B(_02954_),
    .C(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _19465_ (.A0(net1622),
    .A1(net5994),
    .S(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__clkbuf_1 _19466_ (.A(net1734),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _19467_ (.A0(net1396),
    .A1(net6014),
    .S(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__clkbuf_1 _19468_ (.A(net1533),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _19469_ (.A0(net1493),
    .A1(net5996),
    .S(_03345_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _19470_ (.A(net5998),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _19471_ (.A0(net1426),
    .A1(net6003),
    .S(_03345_),
    .X(_03349_));
 sky130_fd_sc_hd__clkbuf_1 _19472_ (.A(net1725),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _19473_ (.A0(net4016),
    .A1(net6005),
    .S(_03345_),
    .X(_03350_));
 sky130_fd_sc_hd__clkbuf_1 _19474_ (.A(net2442),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _19475_ (.A0(net2205),
    .A1(net6007),
    .S(_03345_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_1 _19476_ (.A(net2061),
    .X(_00909_));
 sky130_fd_sc_hd__clkbuf_8 _19477_ (.A(_04459_),
    .X(_03352_));
 sky130_fd_sc_hd__o2bb2a_1 _19478_ (.A1_N(net5940),
    .A2_N(_03139_),
    .B1(_03344_),
    .B2(_02954_),
    .X(_03353_));
 sky130_fd_sc_hd__nor2_1 _19479_ (.A(_03352_),
    .B(net3903),
    .Y(_00910_));
 sky130_fd_sc_hd__or4_4 _19480_ (.A(net1879),
    .B(_02472_),
    .C(_04458_),
    .D(_03344_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _19481_ (.A0(net1622),
    .A1(net6019),
    .S(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__clkbuf_1 _19482_ (.A(net1481),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _19483_ (.A0(net1396),
    .A1(net6050),
    .S(_03354_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _19484_ (.A(net1594),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _19485_ (.A0(net1493),
    .A1(net6010),
    .S(_03354_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _19486_ (.A(net6012),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _19487_ (.A0(net1426),
    .A1(net6056),
    .S(_03354_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_1 _19488_ (.A(net1626),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _19489_ (.A0(net4016),
    .A1(net6024),
    .S(_03354_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_1 _19490_ (.A(net2233),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _19491_ (.A0(net2205),
    .A1(net6021),
    .S(_03354_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_1 _19492_ (.A(net1562),
    .X(_00916_));
 sky130_fd_sc_hd__inv_2 _19493_ (.A(net3519),
    .Y(_03361_));
 sky130_fd_sc_hd__o32a_1 _19494_ (.A1(net1879),
    .A2(_02472_),
    .A3(_03344_),
    .B1(_03141_),
    .B2(net3520),
    .X(_03362_));
 sky130_fd_sc_hd__nor2_1 _19495_ (.A(_03352_),
    .B(net3521),
    .Y(_00917_));
 sky130_fd_sc_hd__and2_1 _19496_ (.A(net1879),
    .B(_02472_),
    .X(_03363_));
 sky130_fd_sc_hd__and2b_1 _19497_ (.A_N(_03344_),
    .B(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__nand2_4 _19498_ (.A(_08092_),
    .B(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__mux2_1 _19499_ (.A0(net1622),
    .A1(net6938),
    .S(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__clkbuf_1 _19500_ (.A(net2448),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _19501_ (.A0(net1396),
    .A1(net6546),
    .S(_03365_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_1 _19502_ (.A(net1644),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _19503_ (.A0(net1493),
    .A1(net6844),
    .S(_03365_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_1 _19504_ (.A(net2257),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _19505_ (.A0(net1426),
    .A1(net5500),
    .S(_03365_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_1 _19506_ (.A(net1635),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _19507_ (.A0(net4016),
    .A1(net6578),
    .S(_03365_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _19508_ (.A(net1672),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _19509_ (.A0(net2205),
    .A1(net6739),
    .S(_03365_),
    .X(_03371_));
 sky130_fd_sc_hd__clkbuf_1 _19510_ (.A(net2147),
    .X(_00923_));
 sky130_fd_sc_hd__a21oi_1 _19511_ (.A1(net5978),
    .A2(_03139_),
    .B1(_03364_),
    .Y(_03372_));
 sky130_fd_sc_hd__nor2_1 _19512_ (.A(_03352_),
    .B(net3218),
    .Y(_00924_));
 sky130_fd_sc_hd__or3_1 _19513_ (.A(_04102_),
    .B(net3084),
    .C(_03344_),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_1 _19514_ (.A(net3085),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _19515_ (.A0(net1622),
    .A1(net5526),
    .S(net3086),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _19516_ (.A(net1641),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _19517_ (.A0(net1396),
    .A1(net5540),
    .S(net3086),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_1 _19518_ (.A(net1737),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _19519_ (.A0(net1493),
    .A1(net6494),
    .S(net3086),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_1 _19520_ (.A(net1494),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19521_ (.A0(net1426),
    .A1(net6486),
    .S(net3086),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _19522_ (.A(net1427),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _19523_ (.A0(net4016),
    .A1(net5535),
    .S(net3086),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _19524_ (.A(net1701),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19525_ (.A0(net3863),
    .A1(net3367),
    .S(net3086),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_1 _19526_ (.A(net3368),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _19527_ (.A0(net3816),
    .A1(net3333),
    .S(net3086),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_1 _19528_ (.A(net3334),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _19529_ (.A0(net3402),
    .A1(net7558),
    .S(net3086),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_1 _19530_ (.A(net3087),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _19531_ (.A0(net2953),
    .A1(net7524),
    .S(net3086),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_1 _19532_ (.A(net7526),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _19533_ (.A0(net3838),
    .A1(net5570),
    .S(net3086),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_1 _19534_ (.A(net1765),
    .X(_00934_));
 sky130_fd_sc_hd__o2bb2a_1 _19535_ (.A1_N(net5943),
    .A2_N(_03139_),
    .B1(_03344_),
    .B2(net3084),
    .X(_03385_));
 sky130_fd_sc_hd__nor2_1 _19536_ (.A(_03352_),
    .B(net3624),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_1 _19537_ (.A(net3770),
    .B(net4833),
    .Y(_03386_));
 sky130_fd_sc_hd__and2_1 _19538_ (.A(net3906),
    .B(_02948_),
    .X(_03387_));
 sky130_fd_sc_hd__and3_2 _19539_ (.A(_08092_),
    .B(_03386_),
    .C(net1777),
    .X(_03388_));
 sky130_fd_sc_hd__mux2_1 _19540_ (.A0(net6613),
    .A1(net1622),
    .S(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_1 _19541_ (.A(net1623),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _19542_ (.A0(net5513),
    .A1(net1396),
    .S(_03388_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _19543_ (.A(net1583),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _19544_ (.A0(net5562),
    .A1(net1493),
    .S(_03388_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _19545_ (.A(net1403),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _19546_ (.A0(net2098),
    .A1(net1426),
    .S(_03388_),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_1 _19547_ (.A(net2099),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _19548_ (.A0(net6544),
    .A1(net4016),
    .S(_03388_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _19549_ (.A(net1743),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _19550_ (.A0(net6960),
    .A1(net2205),
    .S(_03388_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_1 _19551_ (.A(net2224),
    .X(_00941_));
 sky130_fd_sc_hd__a22o_1 _19552_ (.A1(net3978),
    .A2(_03139_),
    .B1(net1777),
    .B2(_03386_),
    .X(_03395_));
 sky130_fd_sc_hd__and2_1 _19553_ (.A(_03320_),
    .B(net3979),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _19554_ (.A(net3980),
    .X(_00942_));
 sky130_fd_sc_hd__nand2_1 _19555_ (.A(net1880),
    .B(net1777),
    .Y(_03397_));
 sky130_fd_sc_hd__nor2_1 _19556_ (.A(_04458_),
    .B(net1881),
    .Y(_03398_));
 sky130_fd_sc_hd__mux2_1 _19557_ (.A0(net6816),
    .A1(net1622),
    .S(net1882),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _19558_ (.A(net1883),
    .X(_00943_));
 sky130_fd_sc_hd__o21a_1 _19559_ (.A1(net3375),
    .A2(_03141_),
    .B1(net1881),
    .X(_03400_));
 sky130_fd_sc_hd__nor2_1 _19560_ (.A(_03352_),
    .B(net3376),
    .Y(_00944_));
 sky130_fd_sc_hd__nand2_1 _19561_ (.A(_03363_),
    .B(net1777),
    .Y(_03401_));
 sky130_fd_sc_hd__nor2_1 _19562_ (.A(_04102_),
    .B(net1778),
    .Y(_03402_));
 sky130_fd_sc_hd__clkbuf_4 _19563_ (.A(net1779),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _19564_ (.A0(net6411),
    .A1(net1622),
    .S(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _19565_ (.A(net1430),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _19566_ (.A0(net6800),
    .A1(net1396),
    .S(_03403_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _19567_ (.A(net1998),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _19568_ (.A0(net6395),
    .A1(net1493),
    .S(_03403_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _19569_ (.A(net6397),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _19570_ (.A0(net7395),
    .A1(net1426),
    .S(_03403_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_1 _19571_ (.A(net3003),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _19572_ (.A0(net5613),
    .A1(net4016),
    .S(_03403_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _19573_ (.A(net2105),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _19574_ (.A0(net7303),
    .A1(net2205),
    .S(_03403_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _19575_ (.A(net2206),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _19576_ (.A0(net7522),
    .A1(net3863),
    .S(_03403_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _19577_ (.A(net2645),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _19578_ (.A0(net7475),
    .A1(net3816),
    .S(_03403_),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _19579_ (.A(net2599),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _19580_ (.A0(net7085),
    .A1(net3402),
    .S(_03403_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _19581_ (.A(net2004),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _19582_ (.A0(net6287),
    .A1(net2953),
    .S(_03403_),
    .X(_03413_));
 sky130_fd_sc_hd__clkbuf_1 _19583_ (.A(net6289),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _19584_ (.A0(net6482),
    .A1(net3838),
    .S(net1779),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _19585_ (.A(net1478),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _19586_ (.A0(net6464),
    .A1(net3745),
    .S(net1779),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _19587_ (.A(net1393),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _19588_ (.A0(net6597),
    .A1(net3596),
    .S(net1779),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _19589_ (.A(net1542),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _19590_ (.A0(net6742),
    .A1(net3562),
    .S(net1779),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _19591_ (.A(net1656),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _19592_ (.A0(net6858),
    .A1(net3738),
    .S(net1779),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _19593_ (.A(net1780),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _19594_ (.A0(net6574),
    .A1(net3592),
    .S(net1779),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _19595_ (.A(net6576),
    .X(_00960_));
 sky130_fd_sc_hd__nand2_1 _19596_ (.A(net6065),
    .B(_03139_),
    .Y(_03420_));
 sky130_fd_sc_hd__a21oi_1 _19597_ (.A1(net1778),
    .A2(net887),
    .B1(_03312_),
    .Y(_00961_));
 sky130_fd_sc_hd__a32o_1 _19598_ (.A1(net3770),
    .A2(_02472_),
    .A3(net1777),
    .B1(_03139_),
    .B2(net3842),
    .X(_03421_));
 sky130_fd_sc_hd__and2_1 _19599_ (.A(_03320_),
    .B(net3843),
    .X(_03422_));
 sky130_fd_sc_hd__clkbuf_1 _19600_ (.A(net3844),
    .X(_00962_));
 sky130_fd_sc_hd__nand2_1 _19601_ (.A(net1030),
    .B(_03139_),
    .Y(_03423_));
 sky130_fd_sc_hd__nand2_1 _19602_ (.A(net4815),
    .B(net4834),
    .Y(_03424_));
 sky130_fd_sc_hd__a21oi_1 _19603_ (.A1(net1031),
    .A2(net4835),
    .B1(_03312_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _19604_ (.A(net4842),
    .B(_03139_),
    .Y(_03425_));
 sky130_fd_sc_hd__a21oi_1 _19605_ (.A1(_02475_),
    .A2(net4844),
    .B1(_03312_),
    .Y(_00964_));
 sky130_fd_sc_hd__nand2_1 _19606_ (.A(net1020),
    .B(_03139_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _19607_ (.A(net4815),
    .B(_03363_),
    .Y(_03427_));
 sky130_fd_sc_hd__a21oi_1 _19608_ (.A1(net1021),
    .A2(net4816),
    .B1(_03312_),
    .Y(_00965_));
 sky130_fd_sc_hd__and4_1 _19609_ (.A(net3770),
    .B(_02472_),
    .C(net92),
    .D(net1777),
    .X(_03428_));
 sky130_fd_sc_hd__buf_2 _19610_ (.A(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__buf_4 _19611_ (.A(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_1 _19612_ (.A0(net6305),
    .A1(net3897),
    .S(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__clkbuf_1 _19613_ (.A(net1302),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _19614_ (.A0(net6285),
    .A1(net1396),
    .S(_03430_),
    .X(_03432_));
 sky130_fd_sc_hd__clkbuf_1 _19615_ (.A(net1378),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _19616_ (.A0(net6253),
    .A1(net1493),
    .S(_03430_),
    .X(_03433_));
 sky130_fd_sc_hd__clkbuf_1 _19617_ (.A(net6255),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _19618_ (.A0(net6263),
    .A1(net1426),
    .S(_03430_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_1 _19619_ (.A(net1248),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _19620_ (.A0(net6448),
    .A1(net4016),
    .S(_03430_),
    .X(_03435_));
 sky130_fd_sc_hd__clkbuf_1 _19621_ (.A(net1545),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _19622_ (.A0(net6367),
    .A1(net2205),
    .S(_03430_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_1 _19623_ (.A(net1375),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _19624_ (.A0(net6297),
    .A1(net3863),
    .S(_03430_),
    .X(_03437_));
 sky130_fd_sc_hd__clkbuf_1 _19625_ (.A(net1296),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _19626_ (.A0(net6542),
    .A1(net3816),
    .S(_03430_),
    .X(_03438_));
 sky130_fd_sc_hd__clkbuf_1 _19627_ (.A(net1669),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _19628_ (.A0(net6281),
    .A1(net3402),
    .S(_03430_),
    .X(_03439_));
 sky130_fd_sc_hd__clkbuf_1 _19629_ (.A(net1279),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _19630_ (.A0(net6566),
    .A1(net2953),
    .S(_03430_),
    .X(_03440_));
 sky130_fd_sc_hd__clkbuf_1 _19631_ (.A(net6568),
    .X(_00975_));
 sky130_fd_sc_hd__buf_4 _19632_ (.A(_03429_),
    .X(_03441_));
 sky130_fd_sc_hd__mux2_1 _19633_ (.A0(net6315),
    .A1(net3838),
    .S(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_1 _19634_ (.A(net1469),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _19635_ (.A0(net6647),
    .A1(net3745),
    .S(_03441_),
    .X(_03443_));
 sky130_fd_sc_hd__clkbuf_1 _19636_ (.A(net1924),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _19637_ (.A0(net6434),
    .A1(net3596),
    .S(_03441_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_1 _19638_ (.A(net1484),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _19639_ (.A0(net6388),
    .A1(net3562),
    .S(_03441_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_1 _19640_ (.A(net1406),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _19641_ (.A0(net6697),
    .A1(net3738),
    .S(_03441_),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_1 _19642_ (.A(net1771),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _19643_ (.A0(net6520),
    .A1(net3592),
    .S(_03441_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _19644_ (.A(net6522),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _19645_ (.A0(net6301),
    .A1(net3556),
    .S(_03441_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_1 _19646_ (.A(net6303),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _19647_ (.A0(net6862),
    .A1(net3674),
    .S(_03441_),
    .X(_03449_));
 sky130_fd_sc_hd__clkbuf_1 _19648_ (.A(net6864),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _19649_ (.A0(net6727),
    .A1(net3866),
    .S(_03441_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _19650_ (.A(net6729),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _19651_ (.A0(net6516),
    .A1(net1447),
    .S(_03441_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_1 _19652_ (.A(net6518),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _19653_ (.A0(net6401),
    .A1(net3478),
    .S(_03429_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_1 _19654_ (.A(net6403),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _19655_ (.A0(net6619),
    .A1(net3481),
    .S(_03429_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _19656_ (.A(net6621),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _19657_ (.A0(net6430),
    .A1(net3583),
    .S(_03429_),
    .X(_03454_));
 sky130_fd_sc_hd__clkbuf_1 _19658_ (.A(net6432),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _19659_ (.A0(net6321),
    .A1(net3631),
    .S(_03429_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_1 _19660_ (.A(net6323),
    .X(_00989_));
 sky130_fd_sc_hd__nor2_4 _19661_ (.A(_04102_),
    .B(net4835),
    .Y(_03456_));
 sky130_fd_sc_hd__buf_4 _19662_ (.A(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__mux2_1 _19663_ (.A0(net6474),
    .A1(net3897),
    .S(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_1 _19664_ (.A(net1308),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _19665_ (.A0(net6313),
    .A1(net4028),
    .S(_03457_),
    .X(_03459_));
 sky130_fd_sc_hd__clkbuf_1 _19666_ (.A(net1311),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _19667_ (.A0(net6341),
    .A1(net1492),
    .S(_03457_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _19668_ (.A(net6343),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _19669_ (.A0(net6504),
    .A1(net4074),
    .S(_03457_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_1 _19670_ (.A(net1695),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _19671_ (.A0(net6440),
    .A1(net4038),
    .S(_03457_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_1 _19672_ (.A(net1347),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _19673_ (.A0(net6419),
    .A1(net2205),
    .S(_03457_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_1 _19674_ (.A(net1417),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _19675_ (.A0(net6599),
    .A1(net3863),
    .S(_03457_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_1 _19676_ (.A(net1692),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _19677_ (.A0(net6532),
    .A1(net3816),
    .S(_03457_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_1 _19678_ (.A(net1801),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _19679_ (.A0(net6399),
    .A1(net3402),
    .S(_03457_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _19680_ (.A(net1553),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _19681_ (.A0(net6351),
    .A1(net2953),
    .S(_03457_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_1 _19682_ (.A(net6353),
    .X(_00999_));
 sky130_fd_sc_hd__buf_4 _19683_ (.A(_03456_),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_1 _19684_ (.A0(net6417),
    .A1(net3838),
    .S(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _19685_ (.A(net1490),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _19686_ (.A0(net6325),
    .A1(net3745),
    .S(_03468_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_1 _19687_ (.A(net1350),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _19688_ (.A0(net6370),
    .A1(net3596),
    .S(_03468_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_1 _19689_ (.A(net1454),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _19690_ (.A0(net6484),
    .A1(net3562),
    .S(_03468_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _19691_ (.A(net1463),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _19692_ (.A0(net6472),
    .A1(net3738),
    .S(_03468_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_1 _19693_ (.A(net1335),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _19694_ (.A0(net6422),
    .A1(net3592),
    .S(_03468_),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_1 _19695_ (.A(net6424),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _19696_ (.A0(net6347),
    .A1(net3556),
    .S(_03468_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _19697_ (.A(net6349),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _19698_ (.A0(net6623),
    .A1(net3674),
    .S(_03468_),
    .X(_03476_));
 sky130_fd_sc_hd__clkbuf_1 _19699_ (.A(net6625),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _19700_ (.A0(net6629),
    .A1(net3866),
    .S(_03468_),
    .X(_03477_));
 sky130_fd_sc_hd__clkbuf_1 _19701_ (.A(net6631),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _19702_ (.A0(net6562),
    .A1(net1447),
    .S(_03468_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_1 _19703_ (.A(net6564),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _19704_ (.A0(net6068),
    .A1(net3478),
    .S(_03456_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_1 _19705_ (.A(net6070),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _19706_ (.A0(net6076),
    .A1(net3481),
    .S(_03456_),
    .X(_03480_));
 sky130_fd_sc_hd__clkbuf_1 _19707_ (.A(net6078),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _19708_ (.A0(net6132),
    .A1(net3583),
    .S(_03456_),
    .X(_03481_));
 sky130_fd_sc_hd__clkbuf_1 _19709_ (.A(net6134),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _19710_ (.A0(net6207),
    .A1(net3631),
    .S(_03456_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_1 _19711_ (.A(net6209),
    .X(_01013_));
 sky130_fd_sc_hd__or2_2 _19712_ (.A(net41),
    .B(net40),
    .X(_03483_));
 sky130_fd_sc_hd__nand2_2 _19713_ (.A(_03122_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__clkbuf_4 _19714_ (.A(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__o211a_1 _19715_ (.A1(net3950),
    .A2(net4997),
    .B1(_08093_),
    .C1(_03485_),
    .X(_01014_));
 sky130_fd_sc_hd__nor2b_1 _19716_ (.A(net7272),
    .B_N(net3220),
    .Y(_03486_));
 sky130_fd_sc_hd__nor2_1 _19717_ (.A(net2309),
    .B(_04102_),
    .Y(_03487_));
 sky130_fd_sc_hd__o21ai_1 _19718_ (.A1(net5280),
    .A2(net7273),
    .B1(net2310),
    .Y(_03488_));
 sky130_fd_sc_hd__a21oi_1 _19719_ (.A1(net5280),
    .A2(net7273),
    .B1(_03488_),
    .Y(_01015_));
 sky130_fd_sc_hd__and3_1 _19720_ (.A(net7685),
    .B(net5280),
    .C(net7273),
    .X(_03489_));
 sky130_fd_sc_hd__a21o_1 _19721_ (.A1(net973),
    .A2(net7273),
    .B1(net3703),
    .X(_03490_));
 sky130_fd_sc_hd__and4bb_1 _19722_ (.A_N(net7655),
    .B_N(net7648),
    .C(net7673),
    .D(net4944),
    .X(_03491_));
 sky130_fd_sc_hd__and4bb_1 _19723_ (.A_N(net5496),
    .B_N(net7685),
    .C(net5280),
    .D(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__a21boi_2 _19724_ (.A1(net7273),
    .A2(_03492_),
    .B1_N(net2310),
    .Y(_03493_));
 sky130_fd_sc_hd__and3b_1 _19725_ (.A_N(_03489_),
    .B(net3704),
    .C(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _19726_ (.A(net3705),
    .X(_01016_));
 sky130_fd_sc_hd__a21boi_1 _19727_ (.A1(net5496),
    .A2(_03489_),
    .B1_N(net2310),
    .Y(_03495_));
 sky130_fd_sc_hd__o21a_1 _19728_ (.A1(net5496),
    .A2(_03489_),
    .B1(_03495_),
    .X(_01017_));
 sky130_fd_sc_hd__and3_1 _19729_ (.A(net7673),
    .B(net5496),
    .C(_03489_),
    .X(_03496_));
 sky130_fd_sc_hd__a21o_1 _19730_ (.A1(net1253),
    .A2(_03489_),
    .B1(net3707),
    .X(_03497_));
 sky130_fd_sc_hd__and3b_1 _19731_ (.A_N(net7674),
    .B(_03493_),
    .C(net3708),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_1 _19732_ (.A(net7676),
    .X(_01018_));
 sky130_fd_sc_hd__and2_1 _19733_ (.A(net7648),
    .B(_03496_),
    .X(_03499_));
 sky130_fd_sc_hd__or2_1 _19734_ (.A(net3921),
    .B(_03496_),
    .X(_03500_));
 sky130_fd_sc_hd__and3b_1 _19735_ (.A_N(net7649),
    .B(net2310),
    .C(net3922),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_1 _19736_ (.A(net3923),
    .X(_01019_));
 sky130_fd_sc_hd__and3_1 _19737_ (.A(net7655),
    .B(net7648),
    .C(_03496_),
    .X(_03502_));
 sky130_fd_sc_hd__or2_1 _19738_ (.A(net3823),
    .B(net7649),
    .X(_03503_));
 sky130_fd_sc_hd__and3b_1 _19739_ (.A_N(net7656),
    .B(net2310),
    .C(net3824),
    .X(_03504_));
 sky130_fd_sc_hd__clkbuf_1 _19740_ (.A(net3825),
    .X(_01020_));
 sky130_fd_sc_hd__o21ai_1 _19741_ (.A1(net4944),
    .A2(net7656),
    .B1(_03493_),
    .Y(_03505_));
 sky130_fd_sc_hd__a21oi_1 _19742_ (.A1(net4944),
    .A2(net7656),
    .B1(_03505_),
    .Y(_01021_));
 sky130_fd_sc_hd__buf_1 _19743_ (.A(clknet_1_0__leaf__05645_),
    .X(_03506_));
 sky130_fd_sc_hd__buf_1 _19744_ (.A(clknet_1_0__leaf__03506_),
    .X(_03507_));
 sky130_fd_sc_hd__inv_2 _19745__27 (.A(clknet_1_1__leaf__03507_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _19746__28 (.A(clknet_1_1__leaf__03507_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _19747__29 (.A(clknet_1_1__leaf__03507_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _19748__30 (.A(clknet_1_1__leaf__03507_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _19749__31 (.A(clknet_1_0__leaf__03507_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _19750__32 (.A(clknet_1_0__leaf__03507_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _19751__33 (.A(clknet_1_0__leaf__03507_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _19752__34 (.A(clknet_1_0__leaf__03507_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _19753__35 (.A(clknet_1_0__leaf__03507_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _19754__36 (.A(clknet_1_0__leaf__03507_),
    .Y(net178));
 sky130_fd_sc_hd__buf_1 _19755_ (.A(clknet_1_0__leaf__03506_),
    .X(_03508_));
 sky130_fd_sc_hd__inv_2 _19756__37 (.A(clknet_1_0__leaf__03508_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _19757__38 (.A(clknet_1_0__leaf__03508_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _19758__39 (.A(clknet_1_0__leaf__03508_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _19759__40 (.A(clknet_1_0__leaf__03508_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _19760__41 (.A(clknet_1_0__leaf__03508_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _19761__42 (.A(clknet_1_1__leaf__03508_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _19762__43 (.A(clknet_1_1__leaf__03508_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _19763__44 (.A(clknet_1_1__leaf__03508_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _19764__45 (.A(clknet_1_1__leaf__03508_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _19765__46 (.A(clknet_1_1__leaf__03508_),
    .Y(net188));
 sky130_fd_sc_hd__buf_1 _19766_ (.A(clknet_1_1__leaf__03506_),
    .X(_03509_));
 sky130_fd_sc_hd__inv_2 _19767__47 (.A(clknet_1_1__leaf__03509_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _19768__48 (.A(clknet_1_1__leaf__03509_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _19769__49 (.A(clknet_1_1__leaf__03509_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _19770__50 (.A(clknet_1_1__leaf__03509_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _19771__51 (.A(clknet_1_0__leaf__03509_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _19772__52 (.A(clknet_1_0__leaf__03509_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _19773__53 (.A(clknet_1_0__leaf__03509_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _19774__54 (.A(clknet_1_0__leaf__03509_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _19775__55 (.A(clknet_1_0__leaf__03509_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _19776__56 (.A(clknet_1_0__leaf__03509_),
    .Y(net198));
 sky130_fd_sc_hd__buf_1 _19777_ (.A(clknet_1_1__leaf__03506_),
    .X(_03510_));
 sky130_fd_sc_hd__inv_2 _19778__57 (.A(clknet_1_0__leaf__03510_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _19779__58 (.A(clknet_1_0__leaf__03510_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _19780__59 (.A(clknet_1_0__leaf__03510_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _19781__60 (.A(clknet_1_0__leaf__03510_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _19782__61 (.A(clknet_1_1__leaf__03510_),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _19783__62 (.A(clknet_1_1__leaf__03510_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _19784__63 (.A(clknet_1_1__leaf__03510_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _19785__64 (.A(clknet_1_1__leaf__03510_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _19786__65 (.A(clknet_1_1__leaf__03510_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _19787__66 (.A(clknet_1_1__leaf__03510_),
    .Y(net208));
 sky130_fd_sc_hd__buf_1 _19788_ (.A(clknet_1_1__leaf__03506_),
    .X(_03511_));
 sky130_fd_sc_hd__inv_2 _19789__67 (.A(clknet_1_1__leaf__03511_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _19790__68 (.A(clknet_1_1__leaf__03511_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _19791__69 (.A(clknet_1_1__leaf__03511_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _19792__70 (.A(clknet_1_1__leaf__03511_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _19793__71 (.A(clknet_1_1__leaf__03511_),
    .Y(net213));
 sky130_fd_sc_hd__inv_2 _19794__72 (.A(clknet_1_1__leaf__03511_),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _19795__73 (.A(clknet_1_0__leaf__03511_),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _19796__74 (.A(clknet_1_0__leaf__03511_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _19797__75 (.A(clknet_1_0__leaf__03511_),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _19798__76 (.A(clknet_1_0__leaf__03511_),
    .Y(net218));
 sky130_fd_sc_hd__buf_1 _19799_ (.A(clknet_1_1__leaf__03506_),
    .X(_03512_));
 sky130_fd_sc_hd__inv_2 _19800__77 (.A(clknet_1_1__leaf__03512_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _19801__78 (.A(clknet_1_1__leaf__03512_),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _19802__79 (.A(clknet_1_1__leaf__03512_),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _19803__80 (.A(clknet_1_1__leaf__03512_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _19804__81 (.A(clknet_1_1__leaf__03512_),
    .Y(net223));
 sky130_fd_sc_hd__inv_2 _19805__82 (.A(clknet_1_0__leaf__03512_),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _19806__83 (.A(clknet_1_0__leaf__03512_),
    .Y(net225));
 sky130_fd_sc_hd__inv_2 _19807__84 (.A(clknet_1_0__leaf__03512_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _19808__85 (.A(clknet_1_0__leaf__03512_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _19809__86 (.A(clknet_1_0__leaf__03512_),
    .Y(net228));
 sky130_fd_sc_hd__buf_1 _19810_ (.A(clknet_1_0__leaf__05645_),
    .X(_03513_));
 sky130_fd_sc_hd__buf_1 _19811_ (.A(clknet_1_1__leaf__03513_),
    .X(_03514_));
 sky130_fd_sc_hd__inv_2 _19812__87 (.A(clknet_1_1__leaf__03514_),
    .Y(net229));
 sky130_fd_sc_hd__inv_2 _19813__88 (.A(clknet_1_1__leaf__03514_),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _19814__89 (.A(clknet_1_1__leaf__03514_),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _19815__90 (.A(clknet_1_1__leaf__03514_),
    .Y(net232));
 sky130_fd_sc_hd__nand2_1 _19816_ (.A(net2310),
    .B(net7273),
    .Y(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _19817_ (.A(net2311),
    .X(_03516_));
 sky130_fd_sc_hd__clkbuf_4 _19818_ (.A(net2312),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_1 _19819_ (.A0(net7312),
    .A1(net3329),
    .S(_03517_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_1 _19820_ (.A(net1815),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _19821_ (.A0(net3329),
    .A1(net3351),
    .S(_03517_),
    .X(_03519_));
 sky130_fd_sc_hd__clkbuf_1 _19822_ (.A(net3211),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _19823_ (.A0(net3351),
    .A1(net7554),
    .S(_03517_),
    .X(_03520_));
 sky130_fd_sc_hd__clkbuf_1 _19824_ (.A(net3231),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _19825_ (.A0(net7554),
    .A1(net3045),
    .S(_03517_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_1 _19826_ (.A(net2507),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _19827_ (.A0(net3045),
    .A1(net6413),
    .S(_03517_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _19828_ (.A(net3046),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _19829_ (.A0(net6413),
    .A1(net1579),
    .S(_03517_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_1 _19830_ (.A(net6415),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _19831_ (.A0(net6661),
    .A1(net1682),
    .S(_03517_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _19832_ (.A(net6663),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _19833_ (.A0(net7310),
    .A1(net3026),
    .S(_03517_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_1 _19834_ (.A(net2263),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _19835_ (.A0(net3026),
    .A1(net3019),
    .S(_03517_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _19836_ (.A(net3027),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _19837_ (.A0(net3019),
    .A1(net3145),
    .S(_03517_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_1 _19838_ (.A(net1857),
    .X(_01095_));
 sky130_fd_sc_hd__clkbuf_4 _19839_ (.A(net2312),
    .X(_03528_));
 sky130_fd_sc_hd__mux2_1 _19840_ (.A0(net3145),
    .A1(net3111),
    .S(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _19841_ (.A(net3146),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _19842_ (.A0(net3111),
    .A1(net7542),
    .S(_03528_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _19843_ (.A(net3102),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _19844_ (.A0(net7542),
    .A1(net2771),
    .S(_03528_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_1 _19845_ (.A(net2870),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _19846_ (.A0(net2771),
    .A1(net6231),
    .S(_03528_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_1 _19847_ (.A(net2772),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _19848_ (.A0(net6231),
    .A1(net6247),
    .S(_03528_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_1 _19849_ (.A(net1183),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _19850_ (.A0(net6247),
    .A1(net3077),
    .S(_03528_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _19851_ (.A(net2808),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _19852_ (.A0(net3077),
    .A1(net7540),
    .S(_03528_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _19853_ (.A(net3078),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _19854_ (.A0(net7540),
    .A1(net1752),
    .S(_03528_),
    .X(_03536_));
 sky130_fd_sc_hd__clkbuf_1 _19855_ (.A(net3064),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _19856_ (.A0(net1752),
    .A1(net7498),
    .S(_03528_),
    .X(_03537_));
 sky130_fd_sc_hd__clkbuf_1 _19857_ (.A(net1707),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _19858_ (.A0(net7498),
    .A1(net6125),
    .S(_03528_),
    .X(_03538_));
 sky130_fd_sc_hd__clkbuf_1 _19859_ (.A(net3156),
    .X(_01105_));
 sky130_fd_sc_hd__clkbuf_4 _19860_ (.A(net2312),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_1 _19861_ (.A0(net6125),
    .A1(net3186),
    .S(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _19862_ (.A(net736),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _19863_ (.A0(net3186),
    .A1(net3056),
    .S(_03539_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_1 _19864_ (.A(net3187),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _19865_ (.A0(net3056),
    .A1(net7443),
    .S(_03539_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_1 _19866_ (.A(net2921),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _19867_ (.A0(net7443),
    .A1(net6512),
    .S(_03539_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _19868_ (.A(net3023),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _19869_ (.A0(net6512),
    .A1(net3173),
    .S(_03539_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _19870_ (.A(net2180),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _19871_ (.A0(net3173),
    .A1(net6649),
    .S(_03539_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _19872_ (.A(net3174),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _19873_ (.A0(net6649),
    .A1(net6357),
    .S(_03539_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _19874_ (.A(net1689),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _19875_ (.A0(net6357),
    .A1(net3195),
    .S(_03539_),
    .X(_03547_));
 sky130_fd_sc_hd__clkbuf_1 _19876_ (.A(net1231),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _19877_ (.A0(net3195),
    .A1(net7556),
    .S(_03539_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_1 _19878_ (.A(net3149),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _19879_ (.A0(net7556),
    .A1(net3342),
    .S(_03539_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _19880_ (.A(net3343),
    .X(_01115_));
 sky130_fd_sc_hd__clkbuf_4 _19881_ (.A(net2312),
    .X(_03550_));
 sky130_fd_sc_hd__mux2_1 _19882_ (.A0(net3342),
    .A1(net3302),
    .S(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _19883_ (.A(net3303),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _19884_ (.A0(net3302),
    .A1(net7516),
    .S(_03550_),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_1 _19885_ (.A(net3234),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _19886_ (.A0(net7516),
    .A1(net3256),
    .S(_03550_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _19887_ (.A(net3257),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _19888_ (.A0(net3256),
    .A1(net6436),
    .S(_03550_),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _19889_ (.A(net3074),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _19890_ (.A0(net6436),
    .A1(net3273),
    .S(_03550_),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_1 _19891_ (.A(net1359),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _19892_ (.A0(net3273),
    .A1(net3298),
    .S(_03550_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _19893_ (.A(net3299),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _19894_ (.A0(net3298),
    .A1(net3125),
    .S(_03550_),
    .X(_03557_));
 sky130_fd_sc_hd__clkbuf_1 _19895_ (.A(net3096),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _19896_ (.A0(net3125),
    .A1(net6731),
    .S(_03550_),
    .X(_03558_));
 sky130_fd_sc_hd__clkbuf_1 _19897_ (.A(net3126),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _19898_ (.A0(net6731),
    .A1(net2934),
    .S(_03550_),
    .X(_03559_));
 sky130_fd_sc_hd__clkbuf_1 _19899_ (.A(net2935),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _19900_ (.A0(net2934),
    .A1(net3320),
    .S(_03550_),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _19901_ (.A(net1152),
    .X(_01125_));
 sky130_fd_sc_hd__clkbuf_4 _19902_ (.A(net2312),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _19903_ (.A0(net3320),
    .A1(net3214),
    .S(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_1 _19904_ (.A(net3321),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _19905_ (.A0(net3214),
    .A1(net7534),
    .S(_03561_),
    .X(_03563_));
 sky130_fd_sc_hd__clkbuf_1 _19906_ (.A(net3215),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _19907_ (.A0(net7534),
    .A1(net3260),
    .S(_03561_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _19908_ (.A(net3167),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _19909_ (.A0(net3260),
    .A1(net2974),
    .S(_03561_),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _19910_ (.A(net3261),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _19911_ (.A0(net2974),
    .A1(net7178),
    .S(_03561_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _19912_ (.A(net2975),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _19913_ (.A0(net7178),
    .A1(net3138),
    .S(_03561_),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _19914_ (.A(net2070),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(net3138),
    .A1(net7453),
    .S(_03561_),
    .X(_03568_));
 sky130_fd_sc_hd__clkbuf_1 _19916_ (.A(net3139),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _19917_ (.A0(net7453),
    .A1(net6744),
    .S(_03561_),
    .X(_03569_));
 sky130_fd_sc_hd__clkbuf_1 _19918_ (.A(net3135),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _19919_ (.A0(net6744),
    .A1(net2801),
    .S(_03561_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _19920_ (.A(net1886),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _19921_ (.A0(net2801),
    .A1(net3227),
    .S(_03561_),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_1 _19922_ (.A(net2802),
    .X(_01135_));
 sky130_fd_sc_hd__clkbuf_4 _19923_ (.A(net2312),
    .X(_03572_));
 sky130_fd_sc_hd__mux2_1 _19924_ (.A0(net3227),
    .A1(net5710),
    .S(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__clkbuf_1 _19925_ (.A(net3228),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _19926_ (.A0(net5710),
    .A1(net7367),
    .S(_03572_),
    .X(_03574_));
 sky130_fd_sc_hd__clkbuf_1 _19927_ (.A(net2412),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _19928_ (.A0(net7367),
    .A1(net3052),
    .S(_03572_),
    .X(_03575_));
 sky130_fd_sc_hd__clkbuf_1 _19929_ (.A(net3053),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _19930_ (.A0(net3052),
    .A1(net6201),
    .S(_03572_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _19931_ (.A(net2543),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _19932_ (.A0(net6201),
    .A1(net3121),
    .S(_03572_),
    .X(_03577_));
 sky130_fd_sc_hd__clkbuf_1 _19933_ (.A(net1111),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _19934_ (.A0(net3121),
    .A1(net7560),
    .S(_03572_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_1 _19935_ (.A(net3122),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _19936_ (.A0(net7560),
    .A1(net3312),
    .S(_03572_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_1 _19937_ (.A(net3313),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _19938_ (.A0(net3312),
    .A1(net3283),
    .S(_03572_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_1 _19939_ (.A(net3284),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _19940_ (.A0(net3283),
    .A1(net3060),
    .S(_03572_),
    .X(_03581_));
 sky130_fd_sc_hd__clkbuf_1 _19941_ (.A(net2861),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _19942_ (.A0(net3060),
    .A1(net7455),
    .S(_03572_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _19943_ (.A(net3061),
    .X(_01145_));
 sky130_fd_sc_hd__buf_4 _19944_ (.A(net2311),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _19945_ (.A0(net7455),
    .A1(net6239),
    .S(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _19946_ (.A(net2904),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _19947_ (.A0(net6239),
    .A1(net3286),
    .S(_03583_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_1 _19948_ (.A(net6241),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _19949_ (.A0(net7520),
    .A1(net7449),
    .S(_03583_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _19950_ (.A(net3287),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _19951_ (.A0(net7449),
    .A1(net3159),
    .S(_03583_),
    .X(_03587_));
 sky130_fd_sc_hd__clkbuf_1 _19952_ (.A(net2713),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _19953_ (.A0(net3159),
    .A1(net2927),
    .S(_03583_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _19954_ (.A(net3160),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _19955_ (.A0(net2927),
    .A1(net7175),
    .S(_03583_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _19956_ (.A(net2928),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _19957_ (.A0(net7175),
    .A1(net5812),
    .S(_03583_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _19958_ (.A(net2191),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _19959_ (.A0(net5812),
    .A1(net3009),
    .S(_03583_),
    .X(_03591_));
 sky130_fd_sc_hd__clkbuf_1 _19960_ (.A(net3010),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _19961_ (.A0(net3009),
    .A1(net5988),
    .S(_03583_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _19962_ (.A(net1568),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _19963_ (.A0(net5988),
    .A1(net3237),
    .S(_03583_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _19964_ (.A(net588),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _19965_ (.A0(net3237),
    .A1(net5764),
    .S(net2312),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_1 _19966_ (.A(net3238),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _19967_ (.A0(net5764),
    .A1(net6327),
    .S(net2312),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_1 _19968_ (.A(net2313),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _19969_ (.A0(net6327),
    .A1(net1869),
    .S(net2312),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_1 _19970_ (.A(net6329),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _19971_ (.A0(net1869),
    .A1(net6665),
    .S(net2312),
    .X(_03597_));
 sky130_fd_sc_hd__clkbuf_1 _19972_ (.A(net6667),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _19973_ (.A0(net54),
    .A1(net1866),
    .S(_03109_),
    .X(_03598_));
 sky130_fd_sc_hd__clkbuf_1 _19974_ (.A(net1867),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _19975_ (.A0(net7312),
    .A1(net1866),
    .S(_09725_),
    .X(_03599_));
 sky130_fd_sc_hd__clkbuf_1 _19976_ (.A(net1809),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _19977_ (.A0(net53),
    .A1(net3199),
    .S(_03109_),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _19978_ (.A(net3200),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _19979_ (.A0(net7506),
    .A1(net3199),
    .S(_08092_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _19980_ (.A(net3049),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _19981_ (.A0(net55),
    .A1(net7425),
    .S(_03109_),
    .X(_03602_));
 sky130_fd_sc_hd__clkbuf_1 _19982_ (.A(net2890),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _19983_ (.A0(net7502),
    .A1(net7425),
    .S(_08092_),
    .X(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _19984_ (.A(net3221),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _19985_ (.A0(net7272),
    .A1(net7502),
    .S(_08092_),
    .X(_03604_));
 sky130_fd_sc_hd__clkbuf_1 _19986_ (.A(net3306),
    .X(_01166_));
 sky130_fd_sc_hd__and2_2 _19987_ (.A(net4997),
    .B(_03484_),
    .X(_03605_));
 sky130_fd_sc_hd__o21a_2 _19988_ (.A1(net40),
    .A2(_03605_),
    .B1(_03122_),
    .X(_03606_));
 sky130_fd_sc_hd__clkbuf_4 _19989_ (.A(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__o21ai_2 _19990_ (.A1(net40),
    .A2(_03605_),
    .B1(_03122_),
    .Y(_03608_));
 sky130_fd_sc_hd__buf_2 _19991_ (.A(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__clkbuf_4 _19992_ (.A(_03484_),
    .X(_03610_));
 sky130_fd_sc_hd__nor2_1 _19993_ (.A(net4168),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__a211o_1 _19994_ (.A1(net5745),
    .A2(_03485_),
    .B1(_03609_),
    .C1(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__o211a_1 _19995_ (.A1(net4168),
    .A2(_03607_),
    .B1(net5746),
    .C1(_03339_),
    .X(_01167_));
 sky130_fd_sc_hd__and2_1 _19996_ (.A(_03122_),
    .B(_03483_),
    .X(_03613_));
 sky130_fd_sc_hd__buf_2 _19997_ (.A(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_4 _19998_ (.A(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__mux2_1 _19999_ (.A0(net5816),
    .A1(_08158_),
    .S(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__or2_1 _20000_ (.A(_03609_),
    .B(net5817),
    .X(_03617_));
 sky130_fd_sc_hd__o211a_1 _20001_ (.A1(net3536),
    .A2(_03607_),
    .B1(net5818),
    .C1(_03339_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _20002_ (.A0(net5835),
    .A1(_08171_),
    .S(_03615_),
    .X(_03618_));
 sky130_fd_sc_hd__or2_1 _20003_ (.A(_03609_),
    .B(net5836),
    .X(_03619_));
 sky130_fd_sc_hd__o211a_1 _20004_ (.A1(net3348),
    .A2(_03607_),
    .B1(net5837),
    .C1(_03339_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _20005_ (.A0(net3269),
    .A1(_08198_),
    .S(_03615_),
    .X(_03620_));
 sky130_fd_sc_hd__or2_1 _20006_ (.A(_03609_),
    .B(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__o211a_1 _20007_ (.A1(net5887),
    .A2(_03607_),
    .B1(_03621_),
    .C1(_03339_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _20008_ (.A0(net3543),
    .A1(_08218_),
    .S(_03614_),
    .X(_03622_));
 sky130_fd_sc_hd__or2_1 _20009_ (.A(_03609_),
    .B(net3544),
    .X(_03623_));
 sky130_fd_sc_hd__o211a_1 _20010_ (.A1(net5904),
    .A2(_03607_),
    .B1(net3545),
    .C1(_03339_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _20011_ (.A0(net4441),
    .A1(_08238_),
    .S(_03614_),
    .X(_03624_));
 sky130_fd_sc_hd__or2_1 _20012_ (.A(_03609_),
    .B(net4442),
    .X(_03625_));
 sky130_fd_sc_hd__o211a_1 _20013_ (.A1(net3339),
    .A2(_03607_),
    .B1(net4443),
    .C1(_03339_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _20014_ (.A0(net5849),
    .A1(_08263_),
    .S(_03614_),
    .X(_03626_));
 sky130_fd_sc_hd__or2_1 _20015_ (.A(_03608_),
    .B(net5850),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_4 _20016_ (.A(_03205_),
    .X(_03628_));
 sky130_fd_sc_hd__o211a_1 _20017_ (.A1(net3457),
    .A2(_03607_),
    .B1(net5851),
    .C1(_03628_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _20018_ (.A0(net4490),
    .A1(_08292_),
    .S(_03614_),
    .X(_03629_));
 sky130_fd_sc_hd__or2_1 _20019_ (.A(_03608_),
    .B(net4491),
    .X(_03630_));
 sky130_fd_sc_hd__o211a_1 _20020_ (.A1(net3461),
    .A2(_03607_),
    .B1(net4492),
    .C1(_03628_),
    .X(_01174_));
 sky130_fd_sc_hd__clkbuf_4 _20021_ (.A(_03615_),
    .X(_03631_));
 sky130_fd_sc_hd__nand2_1 _20022_ (.A(_08297_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__o211a_1 _20023_ (.A1(net5826),
    .A2(_03631_),
    .B1(_03606_),
    .C1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__a211o_1 _20024_ (.A1(net2898),
    .A2(_03609_),
    .B1(net5827),
    .C1(_03316_),
    .X(_01175_));
 sky130_fd_sc_hd__or2_1 _20025_ (.A(net3443),
    .B(_08295_),
    .X(_03634_));
 sky130_fd_sc_hd__nand2_1 _20026_ (.A(_03615_),
    .B(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__a21o_1 _20027_ (.A1(net3443),
    .A2(_08295_),
    .B1(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__o211a_1 _20028_ (.A1(net5868),
    .A2(_03631_),
    .B1(_03606_),
    .C1(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__a211o_1 _20029_ (.A1(net3443),
    .A2(_03609_),
    .B1(net5869),
    .C1(_03316_),
    .X(_01176_));
 sky130_fd_sc_hd__o21ai_1 _20030_ (.A1(net3990),
    .A2(_03634_),
    .B1(_03615_),
    .Y(_03638_));
 sky130_fd_sc_hd__o211a_1 _20031_ (.A1(net5907),
    .A2(_03615_),
    .B1(_03606_),
    .C1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a21oi_1 _20032_ (.A1(_03606_),
    .A2(_03635_),
    .B1(net3991),
    .Y(_03640_));
 sky130_fd_sc_hd__or3_1 _20033_ (.A(_03109_),
    .B(net5908),
    .C(net3992),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _20034_ (.A(net3993),
    .X(_01177_));
 sky130_fd_sc_hd__or3_1 _20035_ (.A(net5915),
    .B(net3990),
    .C(_03634_),
    .X(_03642_));
 sky130_fd_sc_hd__o21ai_1 _20036_ (.A1(net3990),
    .A2(_03634_),
    .B1(net3389),
    .Y(_03643_));
 sky130_fd_sc_hd__a21oi_1 _20037_ (.A1(_03642_),
    .A2(_03643_),
    .B1(_03610_),
    .Y(_03644_));
 sky130_fd_sc_hd__a211o_1 _20038_ (.A1(net4454),
    .A2(_03485_),
    .B1(_03609_),
    .C1(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__o211a_1 _20039_ (.A1(net3389),
    .A2(_03607_),
    .B1(net4455),
    .C1(_03628_),
    .X(_01178_));
 sky130_fd_sc_hd__or2_1 _20040_ (.A(net3431),
    .B(_03642_),
    .X(_03646_));
 sky130_fd_sc_hd__inv_2 _20041_ (.A(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__a21o_1 _20042_ (.A1(net3431),
    .A2(_03642_),
    .B1(_03484_),
    .X(_03648_));
 sky130_fd_sc_hd__o221a_1 _20043_ (.A1(net5898),
    .A2(_03631_),
    .B1(_03647_),
    .B2(_03648_),
    .C1(_03607_),
    .X(_03649_));
 sky130_fd_sc_hd__a211o_1 _20044_ (.A1(net3431),
    .A2(_03609_),
    .B1(net5899),
    .C1(_03316_),
    .X(_01179_));
 sky130_fd_sc_hd__or2_1 _20045_ (.A(net3682),
    .B(_03646_),
    .X(_03650_));
 sky130_fd_sc_hd__a21o_1 _20046_ (.A1(_03483_),
    .A2(_03650_),
    .B1(_03608_),
    .X(_03651_));
 sky130_fd_sc_hd__nor2_1 _20047_ (.A(net7605),
    .B(_03631_),
    .Y(_03652_));
 sky130_fd_sc_hd__a21oi_1 _20048_ (.A1(_03483_),
    .A2(_03646_),
    .B1(_03608_),
    .Y(_03653_));
 sky130_fd_sc_hd__o22a_1 _20049_ (.A1(_03651_),
    .A2(_03652_),
    .B1(_03653_),
    .B2(net3683),
    .X(_03654_));
 sky130_fd_sc_hd__nor2_1 _20050_ (.A(_03352_),
    .B(net7607),
    .Y(_01180_));
 sky130_fd_sc_hd__or2_1 _20051_ (.A(net4019),
    .B(_03484_),
    .X(_03655_));
 sky130_fd_sc_hd__a2bb2o_1 _20052_ (.A1_N(_03650_),
    .A2_N(_03655_),
    .B1(net5784),
    .B2(_03484_),
    .X(_03656_));
 sky130_fd_sc_hd__a22o_1 _20053_ (.A1(net4019),
    .A2(_03651_),
    .B1(_03656_),
    .B2(_03606_),
    .X(_03657_));
 sky130_fd_sc_hd__and2_1 _20054_ (.A(_03320_),
    .B(net4020),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_1 _20055_ (.A(net4021),
    .X(_01181_));
 sky130_fd_sc_hd__o21a_1 _20056_ (.A1(net41),
    .A2(_03605_),
    .B1(_03123_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_4 _20057_ (.A(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__o21ai_4 _20058_ (.A1(net41),
    .A2(_03605_),
    .B1(_03140_),
    .Y(_03661_));
 sky130_fd_sc_hd__clkbuf_4 _20059_ (.A(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__nor2_1 _20060_ (.A(net5929),
    .B(_03610_),
    .Y(_03663_));
 sky130_fd_sc_hd__a211o_1 _20061_ (.A1(net3440),
    .A2(_03485_),
    .B1(_03662_),
    .C1(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__o211a_1 _20062_ (.A1(net5929),
    .A2(_03660_),
    .B1(net3441),
    .C1(_03628_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _20063_ (.A0(net4616),
    .A1(_08145_),
    .S(_03614_),
    .X(_03665_));
 sky130_fd_sc_hd__or2_1 _20064_ (.A(_03661_),
    .B(net4617),
    .X(_03666_));
 sky130_fd_sc_hd__o211a_1 _20065_ (.A1(net3489),
    .A2(_03660_),
    .B1(net4618),
    .C1(_03628_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _20066_ (.A0(net3252),
    .A1(_08177_),
    .S(_03614_),
    .X(_03667_));
 sky130_fd_sc_hd__or2_1 _20067_ (.A(_03661_),
    .B(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__o211a_1 _20068_ (.A1(net5859),
    .A2(_03660_),
    .B1(_03668_),
    .C1(_03628_),
    .X(_01184_));
 sky130_fd_sc_hd__nor2_1 _20069_ (.A(_08190_),
    .B(_03610_),
    .Y(_03669_));
 sky130_fd_sc_hd__a211o_1 _20070_ (.A1(net5750),
    .A2(_03485_),
    .B1(_03662_),
    .C1(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__o211a_1 _20071_ (.A1(net3372),
    .A2(_03660_),
    .B1(net5751),
    .C1(_03628_),
    .X(_01185_));
 sky130_fd_sc_hd__nor2_1 _20072_ (.A(_08214_),
    .B(_03610_),
    .Y(_03671_));
 sky130_fd_sc_hd__a211o_1 _20073_ (.A1(net3414),
    .A2(_03485_),
    .B1(_03662_),
    .C1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__o211a_1 _20074_ (.A1(net4344),
    .A2(_03660_),
    .B1(net3415),
    .C1(_03628_),
    .X(_01186_));
 sky130_fd_sc_hd__nor2_1 _20075_ (.A(_08232_),
    .B(_03610_),
    .Y(_03673_));
 sky130_fd_sc_hd__a211o_1 _20076_ (.A1(net4362),
    .A2(_03485_),
    .B1(_03662_),
    .C1(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__o211a_1 _20077_ (.A1(net3317),
    .A2(_03660_),
    .B1(net4363),
    .C1(_03628_),
    .X(_01187_));
 sky130_fd_sc_hd__nor2_1 _20078_ (.A(_08258_),
    .B(_03610_),
    .Y(_03675_));
 sky130_fd_sc_hd__a211o_1 _20079_ (.A1(net4327),
    .A2(_03485_),
    .B1(_03662_),
    .C1(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__o211a_1 _20080_ (.A1(net3433),
    .A2(_03660_),
    .B1(net4328),
    .C1(_03628_),
    .X(_01188_));
 sky130_fd_sc_hd__nor2_1 _20081_ (.A(_08288_),
    .B(_03610_),
    .Y(_03677_));
 sky130_fd_sc_hd__a211o_1 _20082_ (.A1(net5771),
    .A2(_03485_),
    .B1(_03662_),
    .C1(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_4 _20083_ (.A(_09725_),
    .X(_03679_));
 sky130_fd_sc_hd__o211a_1 _20084_ (.A1(net3445),
    .A2(_03660_),
    .B1(net5772),
    .C1(_03679_),
    .X(_01189_));
 sky130_fd_sc_hd__nand2_1 _20085_ (.A(_08301_),
    .B(_03631_),
    .Y(_03680_));
 sky130_fd_sc_hd__o211a_1 _20086_ (.A1(net2396),
    .A2(_03631_),
    .B1(_03659_),
    .C1(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__a211o_1 _20087_ (.A1(net4284),
    .A2(_03662_),
    .B1(net2397),
    .C1(_03316_),
    .X(_01190_));
 sky130_fd_sc_hd__or2_2 _20088_ (.A(net3326),
    .B(_08299_),
    .X(_03682_));
 sky130_fd_sc_hd__nand2_1 _20089_ (.A(net3326),
    .B(_08299_),
    .Y(_03683_));
 sky130_fd_sc_hd__a21oi_1 _20090_ (.A1(_03682_),
    .A2(_03683_),
    .B1(_03610_),
    .Y(_03684_));
 sky130_fd_sc_hd__a211o_1 _20091_ (.A1(net4901),
    .A2(_03485_),
    .B1(_03662_),
    .C1(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__o211a_1 _20092_ (.A1(net3326),
    .A2(_03660_),
    .B1(net4902),
    .C1(_03679_),
    .X(_01191_));
 sky130_fd_sc_hd__or2_1 _20093_ (.A(net616),
    .B(_03631_),
    .X(_03686_));
 sky130_fd_sc_hd__o21ai_1 _20094_ (.A1(net4748),
    .A2(_03682_),
    .B1(_03615_),
    .Y(_03687_));
 sky130_fd_sc_hd__a22o_1 _20095_ (.A1(net4748),
    .A2(_03682_),
    .B1(_03687_),
    .B2(_03659_),
    .X(_03688_));
 sky130_fd_sc_hd__buf_4 _20096_ (.A(_04458_),
    .X(_03689_));
 sky130_fd_sc_hd__a221o_1 _20097_ (.A1(net4748),
    .A2(_03662_),
    .B1(net617),
    .B2(_03688_),
    .C1(_03689_),
    .X(_01192_));
 sky130_fd_sc_hd__or3_2 _20098_ (.A(net4436),
    .B(net4748),
    .C(_03682_),
    .X(_03690_));
 sky130_fd_sc_hd__o21ai_1 _20099_ (.A1(net4052),
    .A2(_03682_),
    .B1(net4436),
    .Y(_03691_));
 sky130_fd_sc_hd__a21oi_1 _20100_ (.A1(_03690_),
    .A2(_03691_),
    .B1(_03484_),
    .Y(_03692_));
 sky130_fd_sc_hd__a211o_1 _20101_ (.A1(net663),
    .A2(_03610_),
    .B1(_03661_),
    .C1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__o211a_1 _20102_ (.A1(net4436),
    .A2(_03660_),
    .B1(net664),
    .C1(_03679_),
    .X(_01193_));
 sky130_fd_sc_hd__or2_1 _20103_ (.A(net3473),
    .B(_03690_),
    .X(_03694_));
 sky130_fd_sc_hd__inv_2 _20104_ (.A(_03694_),
    .Y(_03695_));
 sky130_fd_sc_hd__a21o_1 _20105_ (.A1(net3473),
    .A2(_03690_),
    .B1(_03484_),
    .X(_03696_));
 sky130_fd_sc_hd__o221a_1 _20106_ (.A1(net4374),
    .A2(_03631_),
    .B1(_03695_),
    .B2(_03696_),
    .C1(_03659_),
    .X(_03697_));
 sky130_fd_sc_hd__a211o_1 _20107_ (.A1(net3473),
    .A2(_03662_),
    .B1(net4375),
    .C1(_03316_),
    .X(_01194_));
 sky130_fd_sc_hd__or2_1 _20108_ (.A(net3552),
    .B(_03694_),
    .X(_03698_));
 sky130_fd_sc_hd__a21o_1 _20109_ (.A1(_03483_),
    .A2(_03698_),
    .B1(_03661_),
    .X(_03699_));
 sky130_fd_sc_hd__nor2_1 _20110_ (.A(net6061),
    .B(_03631_),
    .Y(_03700_));
 sky130_fd_sc_hd__a21oi_1 _20111_ (.A1(_03483_),
    .A2(_03694_),
    .B1(_03661_),
    .Y(_03701_));
 sky130_fd_sc_hd__o22a_1 _20112_ (.A1(_03699_),
    .A2(_03700_),
    .B1(_03701_),
    .B2(net3553),
    .X(_03702_));
 sky130_fd_sc_hd__nor2_1 _20113_ (.A(_03352_),
    .B(net6063),
    .Y(_01195_));
 sky130_fd_sc_hd__o21ai_1 _20114_ (.A1(net3469),
    .A2(_03698_),
    .B1(_03615_),
    .Y(_03703_));
 sky130_fd_sc_hd__o211a_1 _20115_ (.A1(net5759),
    .A2(_03615_),
    .B1(_03659_),
    .C1(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__a21oi_1 _20116_ (.A1(net3469),
    .A2(_03699_),
    .B1(net5760),
    .Y(_03705_));
 sky130_fd_sc_hd__nor2_1 _20117_ (.A(_03352_),
    .B(net5762),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_4 _20118_ (.A(_03123_),
    .B(_03605_),
    .Y(_03706_));
 sky130_fd_sc_hd__clkbuf_4 _20119_ (.A(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__and3_1 _20120_ (.A(net4997),
    .B(_03122_),
    .C(_03484_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_4 _20121_ (.A(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_4 _20122_ (.A(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__buf_2 _20123_ (.A(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__or2_1 _20124_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__o211a_1 _20125_ (.A1(net3407),
    .A2(_03707_),
    .B1(net4626),
    .C1(_03679_),
    .X(_01197_));
 sky130_fd_sc_hd__or2_1 _20126_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(_03711_),
    .X(_03713_));
 sky130_fd_sc_hd__o211a_1 _20127_ (.A1(net7595),
    .A2(_03707_),
    .B1(net4477),
    .C1(_03679_),
    .X(_01198_));
 sky130_fd_sc_hd__or2_1 _20128_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(_03711_),
    .X(_03714_));
 sky130_fd_sc_hd__o211a_1 _20129_ (.A1(net7593),
    .A2(_03707_),
    .B1(net4473),
    .C1(_03679_),
    .X(_01199_));
 sky130_fd_sc_hd__or2_1 _20130_ (.A(net4462),
    .B(_03711_),
    .X(_03715_));
 sky130_fd_sc_hd__o211a_1 _20131_ (.A1(net3362),
    .A2(_03707_),
    .B1(net4463),
    .C1(_03679_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _20132_ (.A0(\rbzero.debug_overlay.facingX[-5] ),
    .A1(net3435),
    .S(_03710_),
    .X(_03716_));
 sky130_fd_sc_hd__or2_1 _20133_ (.A(_03689_),
    .B(net7660),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_1 _20134_ (.A(net3437),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _20135_ (.A0(\rbzero.debug_overlay.facingX[-4] ),
    .A1(net3690),
    .S(_03710_),
    .X(_03718_));
 sky130_fd_sc_hd__or2_1 _20136_ (.A(_03689_),
    .B(net7663),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_1 _20137_ (.A(net3692),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _20138_ (.A0(\rbzero.debug_overlay.facingX[-3] ),
    .A1(net1932),
    .S(_03710_),
    .X(_03720_));
 sky130_fd_sc_hd__or2_1 _20139_ (.A(_03689_),
    .B(net7653),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_1 _20140_ (.A(net3609),
    .X(_01203_));
 sky130_fd_sc_hd__or2_1 _20141_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(_03711_),
    .X(_03722_));
 sky130_fd_sc_hd__o211a_1 _20142_ (.A1(net7334),
    .A2(_03707_),
    .B1(net4595),
    .C1(_03679_),
    .X(_01204_));
 sky130_fd_sc_hd__buf_4 _20143_ (.A(_03709_),
    .X(_03723_));
 sky130_fd_sc_hd__mux2_1 _20144_ (.A0(net3719),
    .A1(net3131),
    .S(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__or2_1 _20145_ (.A(_03689_),
    .B(net3720),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_1 _20146_ (.A(net3721),
    .X(_01205_));
 sky130_fd_sc_hd__or2_1 _20147_ (.A(net4513),
    .B(_03711_),
    .X(_03726_));
 sky130_fd_sc_hd__o211a_1 _20148_ (.A1(net7093),
    .A2(_03707_),
    .B1(net4514),
    .C1(_03679_),
    .X(_01206_));
 sky130_fd_sc_hd__or2_1 _20149_ (.A(net4446),
    .B(_03711_),
    .X(_03727_));
 sky130_fd_sc_hd__o211a_1 _20150_ (.A1(net7083),
    .A2(_03707_),
    .B1(net4447),
    .C1(_03679_),
    .X(_01207_));
 sky130_fd_sc_hd__clkbuf_4 _20151_ (.A(_04458_),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_1 _20152_ (.A0(\rbzero.debug_overlay.facingY[-9] ),
    .A1(net3182),
    .S(_03723_),
    .X(_03729_));
 sky130_fd_sc_hd__or2_1 _20153_ (.A(_03728_),
    .B(net7640),
    .X(_03730_));
 sky130_fd_sc_hd__clkbuf_1 _20154_ (.A(net3688),
    .X(_01208_));
 sky130_fd_sc_hd__or2_1 _20155_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_03711_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_4 _20156_ (.A(_09725_),
    .X(_03732_));
 sky130_fd_sc_hd__o211a_1 _20157_ (.A1(net1057),
    .A2(_03707_),
    .B1(_03731_),
    .C1(_03732_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _20158_ (.A0(\rbzero.debug_overlay.facingY[-7] ),
    .A1(net3289),
    .S(_03723_),
    .X(_03733_));
 sky130_fd_sc_hd__or2_1 _20159_ (.A(_03728_),
    .B(net7627),
    .X(_03734_));
 sky130_fd_sc_hd__clkbuf_1 _20160_ (.A(net3505),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _20161_ (.A0(\rbzero.debug_overlay.facingY[-6] ),
    .A1(net2485),
    .S(_03723_),
    .X(_03735_));
 sky130_fd_sc_hd__or2_1 _20162_ (.A(_03728_),
    .B(net7643),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_1 _20163_ (.A(net3581),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _20164_ (.A0(\rbzero.debug_overlay.facingY[-5] ),
    .A1(net1915),
    .S(_03723_),
    .X(_03737_));
 sky130_fd_sc_hd__or2_1 _20165_ (.A(_03728_),
    .B(net7624),
    .X(_03738_));
 sky130_fd_sc_hd__clkbuf_1 _20166_ (.A(net3882),
    .X(_01212_));
 sky130_fd_sc_hd__or2_1 _20167_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(_03711_),
    .X(_03739_));
 sky130_fd_sc_hd__o211a_1 _20168_ (.A1(net7552),
    .A2(_03707_),
    .B1(net4467),
    .C1(_03732_),
    .X(_01213_));
 sky130_fd_sc_hd__or2_1 _20169_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(_03711_),
    .X(_03740_));
 sky130_fd_sc_hd__o211a_1 _20170_ (.A1(net7544),
    .A2(_03707_),
    .B1(net4487),
    .C1(_03732_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _20171_ (.A0(\rbzero.debug_overlay.facingY[-2] ),
    .A1(net3711),
    .S(_03723_),
    .X(_03741_));
 sky130_fd_sc_hd__or2_1 _20172_ (.A(_03728_),
    .B(net7646),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _20173_ (.A(net3713),
    .X(_01215_));
 sky130_fd_sc_hd__clkbuf_4 _20174_ (.A(_03706_),
    .X(_03743_));
 sky130_fd_sc_hd__buf_2 _20175_ (.A(_03710_),
    .X(_03744_));
 sky130_fd_sc_hd__or2_1 _20176_ (.A(net4416),
    .B(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__o211a_1 _20177_ (.A1(net7565),
    .A2(_03743_),
    .B1(net4417),
    .C1(_03732_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _20178_ (.A0(net7744),
    .A1(net3276),
    .S(_03723_),
    .X(_03746_));
 sky130_fd_sc_hd__or2_1 _20179_ (.A(_03728_),
    .B(net3928),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_1 _20180_ (.A(net3929),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _20181_ (.A0(net7746),
    .A1(net3080),
    .S(_03723_),
    .X(_03748_));
 sky130_fd_sc_hd__or2_1 _20182_ (.A(_03728_),
    .B(net4003),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_1 _20183_ (.A(net4004),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _20184_ (.A0(net3565),
    .A1(net2943),
    .S(_03723_),
    .X(_03750_));
 sky130_fd_sc_hd__or2_1 _20185_ (.A(_03728_),
    .B(net3566),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_1 _20186_ (.A(net3567),
    .X(_01219_));
 sky130_fd_sc_hd__or2_1 _20187_ (.A(_05155_),
    .B(_03744_),
    .X(_03752_));
 sky130_fd_sc_hd__o211a_1 _20188_ (.A1(net4803),
    .A2(_03743_),
    .B1(_03752_),
    .C1(_03732_),
    .X(_01220_));
 sky130_fd_sc_hd__or2_1 _20189_ (.A(net4733),
    .B(_03744_),
    .X(_03753_));
 sky130_fd_sc_hd__o211a_1 _20190_ (.A1(net8103),
    .A2(_03743_),
    .B1(net4734),
    .C1(_03732_),
    .X(_01221_));
 sky130_fd_sc_hd__or2_1 _20191_ (.A(net4501),
    .B(_03744_),
    .X(_03754_));
 sky130_fd_sc_hd__o211a_1 _20192_ (.A1(net2079),
    .A2(_03743_),
    .B1(net4502),
    .C1(_03732_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _20193_ (.A0(net3661),
    .A1(net2161),
    .S(_03723_),
    .X(_03755_));
 sky130_fd_sc_hd__or2_1 _20194_ (.A(_03728_),
    .B(net3662),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _20195_ (.A(net3663),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _20196_ (.A0(net3509),
    .A1(net2125),
    .S(_03709_),
    .X(_03757_));
 sky130_fd_sc_hd__or2_1 _20197_ (.A(_03728_),
    .B(net3510),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _20198_ (.A(net3511),
    .X(_01224_));
 sky130_fd_sc_hd__or2_1 _20199_ (.A(net4698),
    .B(_03744_),
    .X(_03759_));
 sky130_fd_sc_hd__o211a_1 _20200_ (.A1(net7155),
    .A2(_03743_),
    .B1(net4699),
    .C1(_03732_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _20201_ (.A0(net3494),
    .A1(net1875),
    .S(_03709_),
    .X(_03760_));
 sky130_fd_sc_hd__or2_1 _20202_ (.A(_04459_),
    .B(net3495),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _20203_ (.A(net3496),
    .X(_01226_));
 sky130_fd_sc_hd__or2_1 _20204_ (.A(net4554),
    .B(_03744_),
    .X(_03762_));
 sky130_fd_sc_hd__o211a_1 _20205_ (.A1(net2364),
    .A2(_03743_),
    .B1(net4555),
    .C1(_03732_),
    .X(_01227_));
 sky130_fd_sc_hd__or2_1 _20206_ (.A(net4603),
    .B(_03744_),
    .X(_03763_));
 sky130_fd_sc_hd__o211a_1 _20207_ (.A1(net7188),
    .A2(_03743_),
    .B1(net4604),
    .C1(_03732_),
    .X(_01228_));
 sky130_fd_sc_hd__or2_1 _20208_ (.A(_02627_),
    .B(_03744_),
    .X(_03764_));
 sky130_fd_sc_hd__buf_4 _20209_ (.A(_09725_),
    .X(_03765_));
 sky130_fd_sc_hd__o211a_1 _20210_ (.A1(net5476),
    .A2(_03743_),
    .B1(_03764_),
    .C1(_03765_),
    .X(_01229_));
 sky130_fd_sc_hd__or2_1 _20211_ (.A(net4423),
    .B(_03744_),
    .X(_03766_));
 sky130_fd_sc_hd__o211a_1 _20212_ (.A1(net4591),
    .A2(_03743_),
    .B1(_03766_),
    .C1(_03765_),
    .X(_01230_));
 sky130_fd_sc_hd__or2_1 _20213_ (.A(_05164_),
    .B(_03744_),
    .X(_03767_));
 sky130_fd_sc_hd__o211a_1 _20214_ (.A1(net4825),
    .A2(_03743_),
    .B1(_03767_),
    .C1(_03765_),
    .X(_01231_));
 sky130_fd_sc_hd__or2_1 _20215_ (.A(net4635),
    .B(_03710_),
    .X(_03768_));
 sky130_fd_sc_hd__o211a_1 _20216_ (.A1(net7419),
    .A2(_03706_),
    .B1(net4636),
    .C1(_03765_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _20217_ (.A0(net4528),
    .A1(net1862),
    .S(_03709_),
    .X(_03769_));
 sky130_fd_sc_hd__or2_1 _20218_ (.A(_04459_),
    .B(net3539),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _20219_ (.A(net3540),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _20220_ (.A0(net3619),
    .A1(net1573),
    .S(_03709_),
    .X(_03771_));
 sky130_fd_sc_hd__or2_1 _20221_ (.A(_04459_),
    .B(net3620),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _20222_ (.A(net3621),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _20223_ (.A0(net3575),
    .A1(net1970),
    .S(_03709_),
    .X(_03773_));
 sky130_fd_sc_hd__or2_1 _20224_ (.A(_04459_),
    .B(net3576),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_1 _20225_ (.A(net3577),
    .X(_01235_));
 sky130_fd_sc_hd__or2_1 _20226_ (.A(net4686),
    .B(_03710_),
    .X(_03775_));
 sky130_fd_sc_hd__o211a_1 _20227_ (.A1(net6693),
    .A2(_03706_),
    .B1(net4687),
    .C1(_03765_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _20228_ (.A0(net3678),
    .A1(net2468),
    .S(_03709_),
    .X(_03776_));
 sky130_fd_sc_hd__or2_1 _20229_ (.A(_04459_),
    .B(net3679),
    .X(_03777_));
 sky130_fd_sc_hd__clkbuf_1 _20230_ (.A(net3680),
    .X(_01237_));
 sky130_fd_sc_hd__or2_1 _20231_ (.A(net4560),
    .B(_03710_),
    .X(_03778_));
 sky130_fd_sc_hd__o211a_1 _20232_ (.A1(net7490),
    .A2(_03706_),
    .B1(net4561),
    .C1(_03765_),
    .X(_01238_));
 sky130_fd_sc_hd__or2_1 _20233_ (.A(net4709),
    .B(_03710_),
    .X(_03779_));
 sky130_fd_sc_hd__o211a_1 _20234_ (.A1(net7508),
    .A2(_03706_),
    .B1(net4710),
    .C1(_03765_),
    .X(_01239_));
 sky130_fd_sc_hd__or2_1 _20235_ (.A(_02866_),
    .B(_03710_),
    .X(_03780_));
 sky130_fd_sc_hd__o211a_1 _20236_ (.A1(net5045),
    .A2(_03706_),
    .B1(_03780_),
    .C1(_03765_),
    .X(_01240_));
 sky130_fd_sc_hd__a31o_1 _20237_ (.A1(net2310),
    .A2(net7273),
    .A3(_03492_),
    .B1(net3950),
    .X(_03781_));
 sky130_fd_sc_hd__and2_1 _20238_ (.A(_02993_),
    .B(net3951),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_1 _20239_ (.A(net3952),
    .X(_01241_));
 sky130_fd_sc_hd__and4bb_1 _20240_ (.A_N(net3996),
    .B_N(net4128),
    .C(_05050_),
    .D(_05730_),
    .X(_03783_));
 sky130_fd_sc_hd__nand2_1 _20241_ (.A(net4024),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__or4b_1 _20242_ (.A(net4111),
    .B(net4103),
    .C(net5983),
    .D_N(_05673_),
    .X(_03785_));
 sky130_fd_sc_hd__inv_2 _20243_ (.A(net4024),
    .Y(_03786_));
 sky130_fd_sc_hd__inv_2 _20244_ (.A(net4103),
    .Y(_03787_));
 sky130_fd_sc_hd__and4_1 _20245_ (.A(_05673_),
    .B(net4111),
    .C(net4025),
    .D(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__a221oi_1 _20246_ (.A1(net3337),
    .A2(net5984),
    .B1(_03788_),
    .B2(_03783_),
    .C1(_03689_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand3_1 _20247_ (.A(_04648_),
    .B(_04026_),
    .C(_05184_),
    .Y(_03789_));
 sky130_fd_sc_hd__and3_1 _20248_ (.A(net5206),
    .B(_04648_),
    .C(_04027_),
    .X(_03790_));
 sky130_fd_sc_hd__a41o_1 _20249_ (.A1(_04464_),
    .A2(_04684_),
    .A3(_04749_),
    .A4(net5207),
    .B1(net900),
    .X(_03791_));
 sky130_fd_sc_hd__o311a_1 _20250_ (.A1(_04500_),
    .A2(net3642),
    .A3(_03789_),
    .B1(net5208),
    .C1(_08093_),
    .X(_01243_));
 sky130_fd_sc_hd__or3b_1 _20251_ (.A(_05730_),
    .B(_05044_),
    .C_N(net3996),
    .X(_03792_));
 sky130_fd_sc_hd__or4b_1 _20252_ (.A(net4092),
    .B(_03792_),
    .C(net4071),
    .D_N(_03788_),
    .X(_03793_));
 sky130_fd_sc_hd__and2_1 _20253_ (.A(net4122),
    .B(net7619),
    .X(_03794_));
 sky130_fd_sc_hd__nand2_1 _20254_ (.A(net4103),
    .B(net4122),
    .Y(_03795_));
 sky130_fd_sc_hd__o211a_1 _20255_ (.A1(net4103),
    .A2(_03794_),
    .B1(net6001),
    .C1(_03765_),
    .X(_01244_));
 sky130_fd_sc_hd__a31o_1 _20256_ (.A1(net4024),
    .A2(net4103),
    .A3(net4122),
    .B1(_04459_),
    .X(_03796_));
 sky130_fd_sc_hd__a21oi_1 _20257_ (.A1(net4025),
    .A2(net6001),
    .B1(_03796_),
    .Y(_01245_));
 sky130_fd_sc_hd__inv_2 _20258_ (.A(net3970),
    .Y(_03797_));
 sky130_fd_sc_hd__a22o_1 _20259_ (.A1(net4111),
    .A2(_09733_),
    .B1(_03797_),
    .B2(_03794_),
    .X(_03798_));
 sky130_fd_sc_hd__a21o_1 _20260_ (.A1(net4024),
    .A2(net4103),
    .B1(net4111),
    .X(_03799_));
 sky130_fd_sc_hd__and3_1 _20261_ (.A(_09721_),
    .B(_03798_),
    .C(net4112),
    .X(_03800_));
 sky130_fd_sc_hd__clkbuf_1 _20262_ (.A(net4113),
    .X(_01246_));
 sky130_fd_sc_hd__a22o_1 _20263_ (.A1(_05673_),
    .A2(_09733_),
    .B1(net4096),
    .B2(_03794_),
    .X(_03801_));
 sky130_fd_sc_hd__o211a_1 _20264_ (.A1(_05673_),
    .A2(net3970),
    .B1(_03801_),
    .C1(_03765_),
    .X(_01247_));
 sky130_fd_sc_hd__xnor2_1 _20265_ (.A(net4128),
    .B(net4097),
    .Y(_03802_));
 sky130_fd_sc_hd__nor2_1 _20266_ (.A(_03352_),
    .B(net4129),
    .Y(_01248_));
 sky130_fd_sc_hd__and3_1 _20267_ (.A(net4178),
    .B(net4128),
    .C(net4097),
    .X(_03803_));
 sky130_fd_sc_hd__a21o_1 _20268_ (.A1(net4128),
    .A2(net4097),
    .B1(net4178),
    .X(_03804_));
 sky130_fd_sc_hd__and3b_1 _20269_ (.A_N(net4098),
    .B(net4179),
    .C(_09725_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _20270_ (.A(_03805_),
    .X(_01249_));
 sky130_fd_sc_hd__and2_1 _20271_ (.A(net4071),
    .B(net4098),
    .X(_03806_));
 sky130_fd_sc_hd__nor2_1 _20272_ (.A(_03689_),
    .B(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__o21a_1 _20273_ (.A1(net4071),
    .A2(net4098),
    .B1(_03807_),
    .X(_01250_));
 sky130_fd_sc_hd__and3_1 _20274_ (.A(net4092),
    .B(net4071),
    .C(net4098),
    .X(_03808_));
 sky130_fd_sc_hd__nor2_1 _20275_ (.A(_03689_),
    .B(net4099),
    .Y(_03809_));
 sky130_fd_sc_hd__o21a_1 _20276_ (.A1(net4092),
    .A2(_03806_),
    .B1(_03809_),
    .X(_01251_));
 sky130_fd_sc_hd__and2_1 _20277_ (.A(net5966),
    .B(net4099),
    .X(_03810_));
 sky130_fd_sc_hd__nor2_1 _20278_ (.A(_03689_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__o21a_1 _20279_ (.A1(net5966),
    .A2(net4099),
    .B1(_03811_),
    .X(_01252_));
 sky130_fd_sc_hd__o221a_1 _20280_ (.A1(_09733_),
    .A2(_03793_),
    .B1(_03810_),
    .B2(net3996),
    .C1(_09725_),
    .X(_03812_));
 sky130_fd_sc_hd__a21boi_1 _20281_ (.A1(net3996),
    .A2(_03810_),
    .B1_N(_03812_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor2_4 _20282_ (.A(_04102_),
    .B(net4816),
    .Y(_03813_));
 sky130_fd_sc_hd__buf_4 _20283_ (.A(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__mux2_1 _20284_ (.A0(net6275),
    .A1(net3897),
    .S(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _20285_ (.A(net1341),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _20286_ (.A0(net6552),
    .A1(net4028),
    .S(_03814_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _20287_ (.A(net1556),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _20288_ (.A0(net6374),
    .A1(net1492),
    .S(_03814_),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_1 _20289_ (.A(net6376),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _20290_ (.A0(net6409),
    .A1(net4074),
    .S(_03814_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _20291_ (.A(net1305),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _20292_ (.A0(net6510),
    .A1(net4038),
    .S(_03814_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_1 _20293_ (.A(net1460),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _20294_ (.A0(net6450),
    .A1(net2204),
    .S(_03814_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_1 _20295_ (.A(net6452),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _20296_ (.A0(net6283),
    .A1(net3863),
    .S(_03814_),
    .X(_03821_));
 sky130_fd_sc_hd__clkbuf_1 _20297_ (.A(net1264),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _20298_ (.A0(net6378),
    .A1(net3816),
    .S(_03814_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _20299_ (.A(net1442),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _20300_ (.A0(net6265),
    .A1(net3402),
    .S(_03814_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_1 _20301_ (.A(net1215),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _20302_ (.A0(net6309),
    .A1(net2953),
    .S(_03814_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _20303_ (.A(net6311),
    .X(_01263_));
 sky130_fd_sc_hd__buf_4 _20304_ (.A(_03813_),
    .X(_03825_));
 sky130_fd_sc_hd__mux2_1 _20305_ (.A0(net6446),
    .A1(net3838),
    .S(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__clkbuf_1 _20306_ (.A(net1475),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _20307_ (.A0(net6601),
    .A1(net3745),
    .S(_03825_),
    .X(_03827_));
 sky130_fd_sc_hd__clkbuf_1 _20308_ (.A(net1786),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _20309_ (.A0(net6257),
    .A1(net3596),
    .S(_03825_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_1 _20310_ (.A(net1201),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _20311_ (.A0(net6470),
    .A1(net3562),
    .S(_03825_),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_1 _20312_ (.A(net1503),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _20313_ (.A0(net6372),
    .A1(net3738),
    .S(_03825_),
    .X(_03830_));
 sky130_fd_sc_hd__clkbuf_1 _20314_ (.A(net1356),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _20315_ (.A0(net6570),
    .A1(net3592),
    .S(_03825_),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _20316_ (.A(net6572),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _20317_ (.A0(net6496),
    .A1(net3556),
    .S(_03825_),
    .X(_03832_));
 sky130_fd_sc_hd__clkbuf_1 _20318_ (.A(net6498),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _20319_ (.A0(net6677),
    .A1(net3674),
    .S(_03825_),
    .X(_03833_));
 sky130_fd_sc_hd__clkbuf_1 _20320_ (.A(net6679),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _20321_ (.A0(net6317),
    .A1(net3866),
    .S(_03825_),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _20322_ (.A(net6319),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _20323_ (.A0(net6683),
    .A1(net1447),
    .S(_03825_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_1 _20324_ (.A(net6685),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _20325_ (.A0(net6136),
    .A1(net3478),
    .S(_03813_),
    .X(_03836_));
 sky130_fd_sc_hd__clkbuf_1 _20326_ (.A(net6138),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _20327_ (.A0(net6080),
    .A1(net3481),
    .S(_03813_),
    .X(_03837_));
 sky130_fd_sc_hd__clkbuf_1 _20328_ (.A(net6082),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _20329_ (.A0(net6180),
    .A1(net3583),
    .S(_03813_),
    .X(_03838_));
 sky130_fd_sc_hd__clkbuf_1 _20330_ (.A(net6182),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _20331_ (.A0(net6176),
    .A1(net3631),
    .S(_03813_),
    .X(_03839_));
 sky130_fd_sc_hd__clkbuf_1 _20332_ (.A(net6178),
    .X(_01277_));
 sky130_fd_sc_hd__inv_2 _20333__91 (.A(clknet_1_0__leaf__03514_),
    .Y(net233));
 sky130_fd_sc_hd__inv_2 _20334__92 (.A(clknet_1_0__leaf__03514_),
    .Y(net234));
 sky130_fd_sc_hd__inv_2 _20335__93 (.A(clknet_1_0__leaf__03514_),
    .Y(net235));
 sky130_fd_sc_hd__inv_2 _20336__94 (.A(clknet_1_0__leaf__03514_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _20337__95 (.A(clknet_1_0__leaf__03514_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _20338__96 (.A(clknet_1_0__leaf__03514_),
    .Y(net238));
 sky130_fd_sc_hd__buf_1 _20339_ (.A(clknet_1_0__leaf__03513_),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _20340__97 (.A(clknet_1_0__leaf__03840_),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _20341__98 (.A(clknet_1_0__leaf__03840_),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _20342__99 (.A(clknet_1_0__leaf__03840_),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _20343__100 (.A(clknet_1_0__leaf__03840_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _20344__101 (.A(clknet_1_0__leaf__03840_),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _20345__102 (.A(clknet_1_0__leaf__03840_),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _20346__103 (.A(clknet_1_1__leaf__03840_),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _20347__104 (.A(clknet_1_1__leaf__03840_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _20348__105 (.A(clknet_1_1__leaf__03840_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _20349__106 (.A(clknet_1_1__leaf__03840_),
    .Y(net248));
 sky130_fd_sc_hd__buf_1 _20350_ (.A(clknet_1_0__leaf__03513_),
    .X(_03841_));
 sky130_fd_sc_hd__inv_2 _20351__107 (.A(clknet_1_0__leaf__03841_),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _20352__108 (.A(clknet_1_0__leaf__03841_),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _20353__109 (.A(clknet_1_0__leaf__03841_),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _20354__110 (.A(clknet_1_1__leaf__03841_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _20355__111 (.A(clknet_1_1__leaf__03841_),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _20356__112 (.A(clknet_1_1__leaf__03841_),
    .Y(net254));
 sky130_fd_sc_hd__inv_2 _20357__113 (.A(clknet_1_1__leaf__03841_),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _20358__114 (.A(clknet_1_1__leaf__03841_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _20359__115 (.A(clknet_1_0__leaf__03841_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _20360__116 (.A(clknet_1_0__leaf__03841_),
    .Y(net258));
 sky130_fd_sc_hd__buf_1 _20361_ (.A(clknet_1_1__leaf__03513_),
    .X(_03842_));
 sky130_fd_sc_hd__inv_2 _20362__117 (.A(clknet_1_0__leaf__03842_),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _20363__118 (.A(clknet_1_0__leaf__03842_),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _20364__119 (.A(clknet_1_0__leaf__03842_),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _20365__120 (.A(clknet_1_0__leaf__03842_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _20366__121 (.A(clknet_1_1__leaf__03842_),
    .Y(net263));
 sky130_fd_sc_hd__inv_2 _20367__122 (.A(clknet_1_1__leaf__03842_),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _20368__123 (.A(clknet_1_1__leaf__03842_),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _20369__124 (.A(clknet_1_1__leaf__03842_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _20370__125 (.A(clknet_1_1__leaf__03842_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _20371__126 (.A(clknet_1_0__leaf__03842_),
    .Y(net268));
 sky130_fd_sc_hd__buf_1 _20372_ (.A(clknet_1_1__leaf__03513_),
    .X(_03843_));
 sky130_fd_sc_hd__inv_2 _20373__127 (.A(clknet_1_0__leaf__03843_),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _20374__128 (.A(clknet_1_0__leaf__03843_),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _20375__129 (.A(clknet_1_0__leaf__03843_),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _20376__130 (.A(clknet_1_1__leaf__03843_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _20377__131 (.A(clknet_1_1__leaf__03843_),
    .Y(net273));
 sky130_fd_sc_hd__inv_2 _20378__132 (.A(clknet_1_1__leaf__03843_),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _20379__133 (.A(clknet_1_1__leaf__03843_),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _20380__134 (.A(clknet_1_1__leaf__03843_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _20381__135 (.A(clknet_1_0__leaf__03843_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _20382__136 (.A(clknet_1_0__leaf__03843_),
    .Y(net278));
 sky130_fd_sc_hd__buf_1 _20383_ (.A(clknet_1_1__leaf__03513_),
    .X(_03844_));
 sky130_fd_sc_hd__inv_2 _20384__137 (.A(clknet_1_1__leaf__03844_),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _20385__138 (.A(clknet_1_1__leaf__03844_),
    .Y(net280));
 sky130_fd_sc_hd__inv_2 _20386__139 (.A(clknet_1_1__leaf__03844_),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _20387__140 (.A(clknet_1_1__leaf__03844_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _20388__141 (.A(clknet_1_1__leaf__03844_),
    .Y(net283));
 sky130_fd_sc_hd__inv_2 _20389__142 (.A(clknet_1_1__leaf__03844_),
    .Y(net284));
 sky130_fd_sc_hd__inv_2 _20390__143 (.A(clknet_1_0__leaf__03844_),
    .Y(net285));
 sky130_fd_sc_hd__inv_2 _20391__144 (.A(clknet_1_0__leaf__03844_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _20392__145 (.A(clknet_1_0__leaf__03844_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _20393__146 (.A(clknet_1_0__leaf__03844_),
    .Y(net288));
 sky130_fd_sc_hd__buf_1 _20394_ (.A(clknet_1_1__leaf__03513_),
    .X(_03845_));
 sky130_fd_sc_hd__inv_2 _20395__147 (.A(clknet_1_1__leaf__03845_),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _20396__148 (.A(clknet_1_1__leaf__03845_),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _20397__149 (.A(clknet_1_1__leaf__03845_),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _20398__150 (.A(clknet_1_1__leaf__03845_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _20399__151 (.A(clknet_1_1__leaf__03845_),
    .Y(net293));
 sky130_fd_sc_hd__inv_2 _20400__152 (.A(clknet_1_1__leaf__03845_),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _20401__153 (.A(clknet_1_0__leaf__03845_),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _20402__154 (.A(clknet_1_0__leaf__03845_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _20403__155 (.A(clknet_1_0__leaf__03845_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _20404__156 (.A(clknet_1_0__leaf__03845_),
    .Y(net298));
 sky130_fd_sc_hd__buf_1 _20405_ (.A(clknet_1_0__leaf__03513_),
    .X(_03846_));
 sky130_fd_sc_hd__inv_2 _20406__157 (.A(clknet_1_0__leaf__03846_),
    .Y(net299));
 sky130_fd_sc_hd__inv_2 _20407__158 (.A(clknet_1_0__leaf__03846_),
    .Y(net300));
 sky130_fd_sc_hd__inv_2 _20408__159 (.A(clknet_1_1__leaf__03846_),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _20409__160 (.A(clknet_1_1__leaf__03846_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _20410__161 (.A(clknet_1_1__leaf__03846_),
    .Y(net303));
 sky130_fd_sc_hd__inv_2 _20411__162 (.A(clknet_1_1__leaf__03846_),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _20412__163 (.A(clknet_1_1__leaf__03846_),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _20413__164 (.A(clknet_1_1__leaf__03846_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _20414__165 (.A(clknet_1_0__leaf__03846_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _20415__166 (.A(clknet_1_0__leaf__03846_),
    .Y(net308));
 sky130_fd_sc_hd__buf_1 _20416_ (.A(clknet_1_1__leaf__03513_),
    .X(_03847_));
 sky130_fd_sc_hd__inv_2 _20417__167 (.A(clknet_1_1__leaf__03847_),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _20418__168 (.A(clknet_1_1__leaf__03847_),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 _20419__169 (.A(clknet_1_1__leaf__03847_),
    .Y(net311));
 sky130_fd_sc_hd__inv_2 _20420__170 (.A(clknet_1_1__leaf__03847_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _20421__171 (.A(clknet_1_1__leaf__03847_),
    .Y(net313));
 sky130_fd_sc_hd__inv_2 _20422__172 (.A(clknet_1_1__leaf__03847_),
    .Y(net314));
 sky130_fd_sc_hd__inv_2 _20423__173 (.A(clknet_1_0__leaf__03847_),
    .Y(net315));
 sky130_fd_sc_hd__inv_2 _20424__174 (.A(clknet_1_0__leaf__03847_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _20425__175 (.A(clknet_1_0__leaf__03847_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _20426__176 (.A(clknet_1_0__leaf__03847_),
    .Y(net318));
 sky130_fd_sc_hd__buf_1 _20427_ (.A(clknet_1_0__leaf__03513_),
    .X(_03848_));
 sky130_fd_sc_hd__inv_2 _20428__177 (.A(clknet_1_1__leaf__03848_),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 _20429__178 (.A(clknet_1_1__leaf__03848_),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _20430__179 (.A(clknet_1_1__leaf__03848_),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _20431__180 (.A(clknet_1_1__leaf__03848_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _20432__181 (.A(clknet_1_0__leaf__03848_),
    .Y(net323));
 sky130_fd_sc_hd__inv_2 _20433__182 (.A(clknet_1_0__leaf__03848_),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _20434__183 (.A(clknet_1_0__leaf__03848_),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _20435__184 (.A(clknet_1_0__leaf__03848_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _20436__185 (.A(clknet_1_0__leaf__03848_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _20437__186 (.A(clknet_1_0__leaf__03848_),
    .Y(net328));
 sky130_fd_sc_hd__buf_1 _20438_ (.A(clknet_1_0__leaf__05645_),
    .X(_03849_));
 sky130_fd_sc_hd__buf_1 _20439_ (.A(clknet_1_0__leaf__03849_),
    .X(_03850_));
 sky130_fd_sc_hd__inv_2 _20440__187 (.A(clknet_1_1__leaf__03850_),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _20441__188 (.A(clknet_1_1__leaf__03850_),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _20442__189 (.A(clknet_1_1__leaf__03850_),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _20443__190 (.A(clknet_1_1__leaf__03850_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _20444__191 (.A(clknet_1_1__leaf__03850_),
    .Y(net333));
 sky130_fd_sc_hd__inv_2 _20445__192 (.A(clknet_1_1__leaf__03850_),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _20446__193 (.A(clknet_1_0__leaf__03850_),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _20447__194 (.A(clknet_1_0__leaf__03850_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _20448__195 (.A(clknet_1_0__leaf__03850_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _20449__196 (.A(clknet_1_0__leaf__03850_),
    .Y(net338));
 sky130_fd_sc_hd__buf_1 _20450_ (.A(clknet_1_0__leaf__03849_),
    .X(_03851_));
 sky130_fd_sc_hd__inv_2 _20451__197 (.A(clknet_1_1__leaf__03851_),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _20452__198 (.A(clknet_1_1__leaf__03851_),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _20453__199 (.A(clknet_1_1__leaf__03851_),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _20454__200 (.A(clknet_1_1__leaf__03851_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _20455__201 (.A(clknet_1_0__leaf__03851_),
    .Y(net343));
 sky130_fd_sc_hd__inv_2 _20456__202 (.A(clknet_1_0__leaf__03851_),
    .Y(net344));
 sky130_fd_sc_hd__inv_2 _20457__203 (.A(clknet_1_0__leaf__03851_),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _20458__204 (.A(clknet_1_0__leaf__03851_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _20459__205 (.A(clknet_1_0__leaf__03851_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _20460__206 (.A(clknet_1_0__leaf__03851_),
    .Y(net348));
 sky130_fd_sc_hd__buf_1 _20461_ (.A(clknet_1_0__leaf__03849_),
    .X(_03852_));
 sky130_fd_sc_hd__inv_2 _20462__207 (.A(clknet_1_0__leaf__03852_),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _20463__208 (.A(clknet_1_0__leaf__03852_),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _20464__209 (.A(clknet_1_0__leaf__03852_),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _20465__210 (.A(clknet_1_0__leaf__03852_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _20466__211 (.A(clknet_1_0__leaf__03852_),
    .Y(net353));
 sky130_fd_sc_hd__inv_2 _20467__212 (.A(clknet_1_1__leaf__03852_),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _20468__213 (.A(clknet_1_1__leaf__03852_),
    .Y(net355));
 sky130_fd_sc_hd__inv_2 _20469__214 (.A(clknet_1_1__leaf__03852_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _20470__215 (.A(clknet_1_1__leaf__03852_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _20471__216 (.A(clknet_1_1__leaf__03852_),
    .Y(net358));
 sky130_fd_sc_hd__buf_1 _20472_ (.A(clknet_1_0__leaf__03849_),
    .X(_03853_));
 sky130_fd_sc_hd__inv_2 _20473__217 (.A(clknet_1_0__leaf__03853_),
    .Y(net359));
 sky130_fd_sc_hd__inv_2 _20474__218 (.A(clknet_1_0__leaf__03853_),
    .Y(net360));
 sky130_fd_sc_hd__inv_2 _20475__219 (.A(clknet_1_1__leaf__03853_),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 _20476__220 (.A(clknet_1_1__leaf__03853_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _20477__221 (.A(clknet_1_1__leaf__03853_),
    .Y(net363));
 sky130_fd_sc_hd__inv_2 _20478__222 (.A(clknet_1_1__leaf__03853_),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _20479__223 (.A(clknet_1_1__leaf__03853_),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _20480__224 (.A(clknet_1_0__leaf__03853_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _20481__225 (.A(clknet_1_0__leaf__03853_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _20482__226 (.A(clknet_1_1__leaf__03853_),
    .Y(net368));
 sky130_fd_sc_hd__buf_1 _20483_ (.A(clknet_1_1__leaf__03849_),
    .X(_03854_));
 sky130_fd_sc_hd__inv_2 _20484__227 (.A(clknet_1_1__leaf__03854_),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _20485__228 (.A(clknet_1_1__leaf__03854_),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _20486__229 (.A(clknet_1_1__leaf__03854_),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _20487__230 (.A(clknet_1_1__leaf__03854_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _20488__231 (.A(clknet_1_1__leaf__03854_),
    .Y(net373));
 sky130_fd_sc_hd__inv_2 _20489__232 (.A(clknet_1_1__leaf__03854_),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _20490__233 (.A(clknet_1_0__leaf__03854_),
    .Y(net375));
 sky130_fd_sc_hd__inv_2 _20491__234 (.A(clknet_1_0__leaf__03854_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _20492__235 (.A(clknet_1_0__leaf__03854_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _20493__236 (.A(clknet_1_0__leaf__03854_),
    .Y(net378));
 sky130_fd_sc_hd__buf_1 _20494_ (.A(clknet_1_1__leaf__03849_),
    .X(_03855_));
 sky130_fd_sc_hd__inv_2 _20495__237 (.A(clknet_1_1__leaf__03855_),
    .Y(net379));
 sky130_fd_sc_hd__inv_2 _20496__238 (.A(clknet_1_1__leaf__03855_),
    .Y(net380));
 sky130_fd_sc_hd__inv_2 _20497__239 (.A(clknet_1_0__leaf__03855_),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _20498__240 (.A(clknet_1_0__leaf__03855_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _20499__241 (.A(clknet_1_0__leaf__03855_),
    .Y(net383));
 sky130_fd_sc_hd__inv_2 _20500__242 (.A(clknet_1_0__leaf__03855_),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _20501__243 (.A(clknet_1_0__leaf__03855_),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _20502__244 (.A(clknet_1_1__leaf__03855_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _20503__245 (.A(clknet_1_1__leaf__03855_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _20504__246 (.A(clknet_1_1__leaf__03855_),
    .Y(net388));
 sky130_fd_sc_hd__buf_1 _20505_ (.A(clknet_1_1__leaf__03849_),
    .X(_03856_));
 sky130_fd_sc_hd__inv_2 _20506__247 (.A(clknet_1_1__leaf__03856_),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _20507__248 (.A(clknet_1_1__leaf__03856_),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _20508__249 (.A(clknet_1_1__leaf__03856_),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _20509__250 (.A(clknet_1_1__leaf__03856_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _20510__251 (.A(clknet_1_1__leaf__03856_),
    .Y(net393));
 sky130_fd_sc_hd__inv_2 _20511__252 (.A(clknet_1_0__leaf__03856_),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _20512__253 (.A(clknet_1_0__leaf__03856_),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _20513__254 (.A(clknet_1_0__leaf__03856_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _20514__255 (.A(clknet_1_0__leaf__03856_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _20515__256 (.A(clknet_1_0__leaf__03856_),
    .Y(net398));
 sky130_fd_sc_hd__buf_1 _20516_ (.A(clknet_1_1__leaf__03849_),
    .X(_03857_));
 sky130_fd_sc_hd__inv_2 _20517__257 (.A(clknet_1_1__leaf__03857_),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _20518__258 (.A(clknet_1_1__leaf__03857_),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _20519__259 (.A(clknet_1_0__leaf__03857_),
    .Y(net401));
 sky130_fd_sc_hd__inv_2 _20520__260 (.A(clknet_1_0__leaf__03857_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _20521__261 (.A(clknet_1_0__leaf__03857_),
    .Y(net403));
 sky130_fd_sc_hd__inv_2 _20522__262 (.A(clknet_1_0__leaf__03857_),
    .Y(net404));
 sky130_fd_sc_hd__inv_2 _20523__263 (.A(clknet_1_0__leaf__03857_),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _20524__264 (.A(clknet_1_0__leaf__03857_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _20525__265 (.A(clknet_1_1__leaf__03857_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _20526__266 (.A(clknet_1_1__leaf__03857_),
    .Y(net408));
 sky130_fd_sc_hd__buf_1 _20527_ (.A(clknet_1_1__leaf__03849_),
    .X(_03858_));
 sky130_fd_sc_hd__inv_2 _20528__267 (.A(clknet_1_0__leaf__03858_),
    .Y(net409));
 sky130_fd_sc_hd__inv_2 _20529__268 (.A(clknet_1_0__leaf__03858_),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _20530__269 (.A(clknet_1_1__leaf__03858_),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _20531__270 (.A(clknet_1_1__leaf__03858_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _20532__271 (.A(clknet_1_1__leaf__03858_),
    .Y(net413));
 sky130_fd_sc_hd__inv_2 _20533__272 (.A(clknet_1_1__leaf__03858_),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _20534__273 (.A(clknet_1_1__leaf__03858_),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _20535__274 (.A(clknet_1_0__leaf__03858_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _20536__275 (.A(clknet_1_0__leaf__03858_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _20537__276 (.A(clknet_1_0__leaf__03858_),
    .Y(net418));
 sky130_fd_sc_hd__buf_1 _20538_ (.A(clknet_1_0__leaf__03849_),
    .X(_03859_));
 sky130_fd_sc_hd__inv_2 _20539__277 (.A(clknet_1_1__leaf__03859_),
    .Y(net419));
 sky130_fd_sc_hd__inv_2 _20540__278 (.A(clknet_1_1__leaf__03859_),
    .Y(net420));
 sky130_fd_sc_hd__inv_2 _20541__279 (.A(clknet_1_1__leaf__03859_),
    .Y(net421));
 sky130_fd_sc_hd__inv_2 _20542__280 (.A(clknet_1_1__leaf__03859_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _20543__281 (.A(clknet_1_1__leaf__03859_),
    .Y(net423));
 sky130_fd_sc_hd__inv_2 _20544__282 (.A(clknet_1_1__leaf__03859_),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _20545__283 (.A(clknet_1_0__leaf__03859_),
    .Y(net425));
 sky130_fd_sc_hd__inv_2 _20546__284 (.A(clknet_1_0__leaf__03859_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _20547__285 (.A(clknet_1_0__leaf__03859_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _20548__286 (.A(clknet_1_0__leaf__03859_),
    .Y(net428));
 sky130_fd_sc_hd__buf_1 _20549_ (.A(clknet_1_0__leaf__05645_),
    .X(_03860_));
 sky130_fd_sc_hd__buf_1 _20550_ (.A(clknet_1_0__leaf__03860_),
    .X(_03861_));
 sky130_fd_sc_hd__inv_2 _20551__287 (.A(clknet_1_1__leaf__03861_),
    .Y(net429));
 sky130_fd_sc_hd__inv_2 _20552__288 (.A(clknet_1_0__leaf__03861_),
    .Y(net430));
 sky130_fd_sc_hd__inv_2 _20553__289 (.A(clknet_1_0__leaf__03861_),
    .Y(net431));
 sky130_fd_sc_hd__inv_2 _20554__290 (.A(clknet_1_0__leaf__03861_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _20555__291 (.A(clknet_1_0__leaf__03861_),
    .Y(net433));
 sky130_fd_sc_hd__inv_2 _20556__292 (.A(clknet_1_0__leaf__03861_),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _20557__293 (.A(clknet_1_0__leaf__03861_),
    .Y(net435));
 sky130_fd_sc_hd__inv_2 _20558__294 (.A(clknet_1_1__leaf__03861_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _20559__295 (.A(clknet_1_1__leaf__03861_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _20560__296 (.A(clknet_1_1__leaf__03861_),
    .Y(net438));
 sky130_fd_sc_hd__buf_1 _20561_ (.A(clknet_1_0__leaf__03860_),
    .X(_03862_));
 sky130_fd_sc_hd__inv_2 _20562__297 (.A(clknet_1_0__leaf__03862_),
    .Y(net439));
 sky130_fd_sc_hd__inv_2 _20563__298 (.A(clknet_1_0__leaf__03862_),
    .Y(net440));
 sky130_fd_sc_hd__inv_2 _20564__299 (.A(clknet_1_0__leaf__03862_),
    .Y(net441));
 sky130_fd_sc_hd__inv_2 _20565__300 (.A(clknet_1_0__leaf__03862_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _20566__301 (.A(clknet_1_0__leaf__03862_),
    .Y(net443));
 sky130_fd_sc_hd__inv_2 _20567__302 (.A(clknet_1_1__leaf__03862_),
    .Y(net444));
 sky130_fd_sc_hd__inv_2 _20568__303 (.A(clknet_1_1__leaf__03862_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _20569__304 (.A(clknet_1_1__leaf__03862_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _20570__305 (.A(clknet_1_1__leaf__03862_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _20571__306 (.A(clknet_1_1__leaf__03862_),
    .Y(net448));
 sky130_fd_sc_hd__buf_1 _20572_ (.A(clknet_1_1__leaf__03860_),
    .X(_03863_));
 sky130_fd_sc_hd__inv_2 _20573__307 (.A(clknet_1_0__leaf__03863_),
    .Y(net449));
 sky130_fd_sc_hd__inv_2 _20574__308 (.A(clknet_1_0__leaf__03863_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _20575__309 (.A(clknet_1_0__leaf__03863_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _20576__310 (.A(clknet_1_0__leaf__03863_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _20577__311 (.A(clknet_1_0__leaf__03863_),
    .Y(net453));
 sky130_fd_sc_hd__inv_2 _20578__312 (.A(clknet_1_1__leaf__03863_),
    .Y(net454));
 sky130_fd_sc_hd__inv_2 _20579__313 (.A(clknet_1_1__leaf__03863_),
    .Y(net455));
 sky130_fd_sc_hd__inv_2 _20580__314 (.A(clknet_1_1__leaf__03863_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _20581__315 (.A(clknet_1_1__leaf__03863_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _20582__316 (.A(clknet_1_1__leaf__03863_),
    .Y(net458));
 sky130_fd_sc_hd__buf_1 _20583_ (.A(clknet_1_1__leaf__03860_),
    .X(_03864_));
 sky130_fd_sc_hd__inv_2 _20584__317 (.A(clknet_1_0__leaf__03864_),
    .Y(net459));
 sky130_fd_sc_hd__inv_2 _20585__318 (.A(clknet_1_0__leaf__03864_),
    .Y(net460));
 sky130_fd_sc_hd__inv_2 _20586__319 (.A(clknet_1_0__leaf__03864_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _20587__320 (.A(clknet_1_0__leaf__03864_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _20588__321 (.A(clknet_1_1__leaf__03864_),
    .Y(net463));
 sky130_fd_sc_hd__inv_2 _20589__322 (.A(clknet_1_1__leaf__03864_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _20590__323 (.A(clknet_1_1__leaf__03864_),
    .Y(net465));
 sky130_fd_sc_hd__inv_2 _20591__324 (.A(clknet_1_1__leaf__03864_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _20592__325 (.A(clknet_1_0__leaf__03864_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _20593__326 (.A(clknet_1_0__leaf__03864_),
    .Y(net468));
 sky130_fd_sc_hd__buf_1 _20594_ (.A(clknet_1_1__leaf__03860_),
    .X(_03865_));
 sky130_fd_sc_hd__inv_2 _20595__327 (.A(clknet_1_0__leaf__03865_),
    .Y(net469));
 sky130_fd_sc_hd__inv_2 _20596__328 (.A(clknet_1_0__leaf__03865_),
    .Y(net470));
 sky130_fd_sc_hd__inv_2 _20597__329 (.A(clknet_1_0__leaf__03865_),
    .Y(net471));
 sky130_fd_sc_hd__inv_2 _20598__330 (.A(clknet_1_0__leaf__03865_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _20599__331 (.A(clknet_1_0__leaf__03865_),
    .Y(net473));
 sky130_fd_sc_hd__inv_2 _20600__332 (.A(clknet_1_1__leaf__03865_),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _20601__333 (.A(clknet_1_1__leaf__03865_),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _20602__334 (.A(clknet_1_1__leaf__03865_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _20603__335 (.A(clknet_1_1__leaf__03865_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _20604__336 (.A(clknet_1_1__leaf__03865_),
    .Y(net478));
 sky130_fd_sc_hd__buf_1 _20605_ (.A(clknet_1_1__leaf__03860_),
    .X(_03866_));
 sky130_fd_sc_hd__inv_2 _20606__337 (.A(clknet_1_0__leaf__03866_),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _20607__338 (.A(clknet_1_0__leaf__03866_),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _20608__339 (.A(clknet_1_0__leaf__03866_),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _20609__340 (.A(clknet_1_0__leaf__03866_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _20610__341 (.A(clknet_1_1__leaf__03866_),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _20611__342 (.A(clknet_1_1__leaf__03866_),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _20612__343 (.A(clknet_1_1__leaf__03866_),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _20613__344 (.A(clknet_1_1__leaf__03866_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _20614__345 (.A(clknet_1_1__leaf__03866_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _20615__346 (.A(clknet_1_1__leaf__03866_),
    .Y(net488));
 sky130_fd_sc_hd__buf_1 _20616_ (.A(clknet_1_0__leaf__03860_),
    .X(_03867_));
 sky130_fd_sc_hd__inv_2 _20617__347 (.A(clknet_1_1__leaf__03867_),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _20618__348 (.A(clknet_1_1__leaf__03867_),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _20619__349 (.A(clknet_1_0__leaf__03867_),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _20620__350 (.A(clknet_1_0__leaf__03867_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _20621__351 (.A(clknet_1_1__leaf__03867_),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _20622__352 (.A(clknet_1_1__leaf__03867_),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _20623__353 (.A(clknet_1_1__leaf__03867_),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _20624__354 (.A(clknet_1_0__leaf__03867_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _20625__355 (.A(clknet_1_0__leaf__03867_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _20626__356 (.A(clknet_1_0__leaf__03867_),
    .Y(net498));
 sky130_fd_sc_hd__buf_1 _20627_ (.A(clknet_1_0__leaf__03860_),
    .X(_03868_));
 sky130_fd_sc_hd__inv_2 _20628__357 (.A(clknet_1_0__leaf__03868_),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _20629__358 (.A(clknet_1_1__leaf__03868_),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _20630__359 (.A(clknet_1_1__leaf__03868_),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _20631__360 (.A(clknet_1_1__leaf__03868_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _20632__361 (.A(clknet_1_1__leaf__03868_),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _20633__362 (.A(clknet_1_0__leaf__03868_),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _20634__363 (.A(clknet_1_0__leaf__03868_),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _20635__364 (.A(clknet_1_0__leaf__03868_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _20636__365 (.A(clknet_1_0__leaf__03868_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _20637__366 (.A(clknet_1_0__leaf__03868_),
    .Y(net508));
 sky130_fd_sc_hd__buf_1 _20638_ (.A(clknet_1_0__leaf__03860_),
    .X(_03869_));
 sky130_fd_sc_hd__inv_2 _20639__367 (.A(clknet_1_0__leaf__03869_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _20640__368 (.A(clknet_1_0__leaf__03869_),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _20641__369 (.A(clknet_1_0__leaf__03869_),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _20642__370 (.A(clknet_1_0__leaf__03869_),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _20643__371 (.A(clknet_1_1__leaf__03869_),
    .Y(net513));
 sky130_fd_sc_hd__inv_2 _20644__372 (.A(clknet_1_1__leaf__03869_),
    .Y(net514));
 sky130_fd_sc_hd__inv_2 _20645__373 (.A(clknet_1_1__leaf__03869_),
    .Y(net515));
 sky130_fd_sc_hd__inv_2 _20646__374 (.A(clknet_1_1__leaf__03869_),
    .Y(net516));
 sky130_fd_sc_hd__inv_2 _20647__375 (.A(clknet_1_1__leaf__03869_),
    .Y(net517));
 sky130_fd_sc_hd__inv_2 _20648__376 (.A(clknet_1_1__leaf__03869_),
    .Y(net518));
 sky130_fd_sc_hd__buf_1 _20649_ (.A(clknet_1_0__leaf__03860_),
    .X(_03870_));
 sky130_fd_sc_hd__inv_2 _20650__377 (.A(clknet_1_0__leaf__03870_),
    .Y(net519));
 sky130_fd_sc_hd__inv_2 _20651__378 (.A(clknet_1_0__leaf__03870_),
    .Y(net520));
 sky130_fd_sc_hd__inv_2 _20652__379 (.A(clknet_1_0__leaf__03870_),
    .Y(net521));
 sky130_fd_sc_hd__inv_2 _20653__380 (.A(clknet_1_0__leaf__03870_),
    .Y(net522));
 sky130_fd_sc_hd__inv_2 _20654__381 (.A(clknet_1_0__leaf__03870_),
    .Y(net523));
 sky130_fd_sc_hd__inv_2 _20655__382 (.A(clknet_1_1__leaf__03870_),
    .Y(net524));
 sky130_fd_sc_hd__inv_2 _20656__383 (.A(clknet_1_1__leaf__03870_),
    .Y(net525));
 sky130_fd_sc_hd__inv_2 _20657__384 (.A(clknet_1_1__leaf__03870_),
    .Y(net526));
 sky130_fd_sc_hd__inv_2 _20658__385 (.A(clknet_1_1__leaf__03870_),
    .Y(net527));
 sky130_fd_sc_hd__inv_2 _20659__386 (.A(clknet_1_1__leaf__03870_),
    .Y(net528));
 sky130_fd_sc_hd__buf_1 _20660_ (.A(clknet_1_0__leaf__05645_),
    .X(_03871_));
 sky130_fd_sc_hd__inv_2 _20661__7 (.A(clknet_1_1__leaf__03871_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _20662__8 (.A(clknet_1_1__leaf__03871_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _20663__9 (.A(clknet_1_1__leaf__03871_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _20664__10 (.A(clknet_1_1__leaf__03871_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _20665__11 (.A(clknet_1_0__leaf__03871_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _20666__12 (.A(clknet_1_0__leaf__03871_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _20667__13 (.A(clknet_1_0__leaf__03871_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _20668__14 (.A(clknet_1_0__leaf__03871_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _20669__15 (.A(clknet_1_0__leaf__03871_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _20670__16 (.A(clknet_1_0__leaf__03871_),
    .Y(net158));
 sky130_fd_sc_hd__buf_1 _20671_ (.A(clknet_1_0__leaf__05645_),
    .X(_03872_));
 sky130_fd_sc_hd__inv_2 _20672__17 (.A(clknet_1_1__leaf__03872_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _20673__18 (.A(clknet_1_1__leaf__03872_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _20674__19 (.A(clknet_1_1__leaf__03872_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _20675__20 (.A(clknet_1_1__leaf__03872_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _20676__21 (.A(clknet_1_0__leaf__03872_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _20677__22 (.A(clknet_1_0__leaf__03872_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _20678__23 (.A(clknet_1_0__leaf__03872_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _20679__24 (.A(clknet_1_0__leaf__03872_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _20680__25 (.A(clknet_1_0__leaf__03872_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _20681__26 (.A(clknet_1_0__leaf__03872_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _20682__3 (.A(clknet_1_0__leaf__03506_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _20683__4 (.A(clknet_1_0__leaf__03506_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _20684__5 (.A(clknet_1_0__leaf__03506_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _20685__6 (.A(clknet_1_0__leaf__03506_),
    .Y(net148));
 sky130_fd_sc_hd__nor2_1 _20686_ (.A(net4922),
    .B(net63),
    .Y(_01598_));
 sky130_fd_sc_hd__xnor2_1 _20687_ (.A(net6058),
    .B(net4922),
    .Y(_03873_));
 sky130_fd_sc_hd__nor2_1 _20688_ (.A(_03352_),
    .B(net920),
    .Y(_01599_));
 sky130_fd_sc_hd__clkbuf_4 _20689_ (.A(_09727_),
    .X(_03874_));
 sky130_fd_sc_hd__or2_1 _20690_ (.A(net777),
    .B(net4968),
    .X(_03875_));
 sky130_fd_sc_hd__nand2_1 _20691_ (.A(net777),
    .B(net4968),
    .Y(_03876_));
 sky130_fd_sc_hd__clkbuf_4 _20692_ (.A(_03109_),
    .X(_03877_));
 sky130_fd_sc_hd__a32o_1 _20693_ (.A1(_03874_),
    .A2(_03875_),
    .A3(_03876_),
    .B1(_03877_),
    .B2(net4968),
    .X(_01600_));
 sky130_fd_sc_hd__clkbuf_4 _20694_ (.A(_09727_),
    .X(_03878_));
 sky130_fd_sc_hd__or2_1 _20695_ (.A(net756),
    .B(net4984),
    .X(_03879_));
 sky130_fd_sc_hd__nand2_1 _20696_ (.A(net756),
    .B(net4984),
    .Y(_03880_));
 sky130_fd_sc_hd__nand3b_1 _20697_ (.A_N(_03876_),
    .B(_03879_),
    .C(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__a21bo_1 _20698_ (.A1(_03879_),
    .A2(_03880_),
    .B1_N(_03876_),
    .X(_03882_));
 sky130_fd_sc_hd__clkbuf_4 _20699_ (.A(_03109_),
    .X(_03883_));
 sky130_fd_sc_hd__a32o_1 _20700_ (.A1(_03878_),
    .A2(_03881_),
    .A3(_03882_),
    .B1(_03883_),
    .B2(net4984),
    .X(_01601_));
 sky130_fd_sc_hd__and2_1 _20701_ (.A(_03880_),
    .B(_03881_),
    .X(_03884_));
 sky130_fd_sc_hd__nor2_1 _20702_ (.A(net967),
    .B(net5384),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _20703_ (.A(net967),
    .B(net5384),
    .Y(_03886_));
 sky130_fd_sc_hd__and2b_1 _20704_ (.A_N(_03885_),
    .B(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__xnor2_1 _20705_ (.A(_03884_),
    .B(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__a22o_1 _20706_ (.A1(net5384),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03888_),
    .X(_01602_));
 sky130_fd_sc_hd__o21a_1 _20707_ (.A1(_03884_),
    .A2(_03885_),
    .B1(_03886_),
    .X(_03889_));
 sky130_fd_sc_hd__nor2_1 _20708_ (.A(net754),
    .B(net5400),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _20709_ (.A(net754),
    .B(net5400),
    .Y(_03891_));
 sky130_fd_sc_hd__and2b_1 _20710_ (.A_N(_03890_),
    .B(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__xnor2_1 _20711_ (.A(_03889_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__a22o_1 _20712_ (.A1(net5400),
    .A2(_03877_),
    .B1(_03874_),
    .B2(net8232),
    .X(_01603_));
 sky130_fd_sc_hd__o21a_1 _20713_ (.A1(_03889_),
    .A2(_03890_),
    .B1(_03891_),
    .X(_03894_));
 sky130_fd_sc_hd__nor2_1 _20714_ (.A(net960),
    .B(net5380),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_1 _20715_ (.A(net960),
    .B(net5380),
    .Y(_03896_));
 sky130_fd_sc_hd__and2b_1 _20716_ (.A_N(_03895_),
    .B(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__xnor2_1 _20717_ (.A(_03894_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__a22o_1 _20718_ (.A1(net5380),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03898_),
    .X(_01604_));
 sky130_fd_sc_hd__o21a_1 _20719_ (.A1(_03894_),
    .A2(_03895_),
    .B1(_03896_),
    .X(_03899_));
 sky130_fd_sc_hd__nor2_1 _20720_ (.A(net1048),
    .B(net5404),
    .Y(_03900_));
 sky130_fd_sc_hd__nand2_1 _20721_ (.A(net1048),
    .B(net5404),
    .Y(_03901_));
 sky130_fd_sc_hd__and2b_1 _20722_ (.A_N(_03900_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__xnor2_1 _20723_ (.A(_03899_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__a22o_1 _20724_ (.A1(net5404),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03903_),
    .X(_01605_));
 sky130_fd_sc_hd__o21a_1 _20725_ (.A1(_03899_),
    .A2(_03900_),
    .B1(_03901_),
    .X(_03904_));
 sky130_fd_sc_hd__nor2_1 _20726_ (.A(net1120),
    .B(net5252),
    .Y(_03905_));
 sky130_fd_sc_hd__nand2_1 _20727_ (.A(net1120),
    .B(net5252),
    .Y(_03906_));
 sky130_fd_sc_hd__and2b_1 _20728_ (.A_N(_03905_),
    .B(_03906_),
    .X(_03907_));
 sky130_fd_sc_hd__xnor2_1 _20729_ (.A(_03904_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__a22o_1 _20730_ (.A1(net5252),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03908_),
    .X(_01606_));
 sky130_fd_sc_hd__o21a_1 _20731_ (.A1(_03904_),
    .A2(_03905_),
    .B1(_03906_),
    .X(_03909_));
 sky130_fd_sc_hd__nor2_1 _20732_ (.A(net1106),
    .B(net5340),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _20733_ (.A(net1106),
    .B(net5340),
    .Y(_03911_));
 sky130_fd_sc_hd__and2b_1 _20734_ (.A_N(_03910_),
    .B(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__xnor2_1 _20735_ (.A(_03909_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__a22o_1 _20736_ (.A1(net5340),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03913_),
    .X(_01607_));
 sky130_fd_sc_hd__o21a_1 _20737_ (.A1(_03909_),
    .A2(_03910_),
    .B1(_03911_),
    .X(_03914_));
 sky130_fd_sc_hd__nor2_1 _20738_ (.A(net896),
    .B(net5376),
    .Y(_03915_));
 sky130_fd_sc_hd__nand2_1 _20739_ (.A(net896),
    .B(net5376),
    .Y(_03916_));
 sky130_fd_sc_hd__and2b_1 _20740_ (.A_N(_03915_),
    .B(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__xnor2_1 _20741_ (.A(_03914_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__a22o_1 _20742_ (.A1(net5376),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03918_),
    .X(_01608_));
 sky130_fd_sc_hd__o21ai_2 _20743_ (.A1(_03914_),
    .A2(_03915_),
    .B1(_03916_),
    .Y(_03919_));
 sky130_fd_sc_hd__or2_1 _20744_ (.A(net834),
    .B(net4972),
    .X(_03920_));
 sky130_fd_sc_hd__nand2_1 _20745_ (.A(net834),
    .B(net4972),
    .Y(_03921_));
 sky130_fd_sc_hd__nand3_1 _20746_ (.A(_03919_),
    .B(_03920_),
    .C(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__a21o_1 _20747_ (.A1(_03920_),
    .A2(_03921_),
    .B1(_03919_),
    .X(_03923_));
 sky130_fd_sc_hd__a32o_1 _20748_ (.A1(_03878_),
    .A2(_03922_),
    .A3(_03923_),
    .B1(_03883_),
    .B2(net4972),
    .X(_01609_));
 sky130_fd_sc_hd__or2_1 _20749_ (.A(net822),
    .B(net4980),
    .X(_03924_));
 sky130_fd_sc_hd__nand2_1 _20750_ (.A(net822),
    .B(net4980),
    .Y(_03925_));
 sky130_fd_sc_hd__a21bo_1 _20751_ (.A1(_03919_),
    .A2(_03920_),
    .B1_N(_03921_),
    .X(_03926_));
 sky130_fd_sc_hd__and3_1 _20752_ (.A(_03924_),
    .B(_03925_),
    .C(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__inv_2 _20753_ (.A(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__a21o_1 _20754_ (.A1(_03924_),
    .A2(_03925_),
    .B1(_03926_),
    .X(_03929_));
 sky130_fd_sc_hd__a32o_1 _20755_ (.A1(_03878_),
    .A2(_03928_),
    .A3(net8197),
    .B1(_03883_),
    .B2(net4980),
    .X(_01610_));
 sky130_fd_sc_hd__or2_1 _20756_ (.A(net984),
    .B(net5448),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_1 _20757_ (.A(net984),
    .B(net5448),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _20758_ (.A(_03925_),
    .B(_03928_),
    .Y(_03932_));
 sky130_fd_sc_hd__a21o_1 _20759_ (.A1(_03930_),
    .A2(_03931_),
    .B1(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__and3_1 _20760_ (.A(_03930_),
    .B(_03931_),
    .C(_03932_),
    .X(_03934_));
 sky130_fd_sc_hd__inv_2 _20761_ (.A(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__a32o_1 _20762_ (.A1(_03878_),
    .A2(net8181),
    .A3(_03935_),
    .B1(_03883_),
    .B2(net5448),
    .X(_01611_));
 sky130_fd_sc_hd__or2_1 _20763_ (.A(net948),
    .B(net5492),
    .X(_03936_));
 sky130_fd_sc_hd__nand2_1 _20764_ (.A(net948),
    .B(net5492),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _20765_ (.A(_03931_),
    .B(_03935_),
    .Y(_03938_));
 sky130_fd_sc_hd__and3_1 _20766_ (.A(_03936_),
    .B(_03937_),
    .C(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__inv_2 _20767_ (.A(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__a21o_1 _20768_ (.A1(_03936_),
    .A2(_03937_),
    .B1(_03938_),
    .X(_03941_));
 sky130_fd_sc_hd__a32o_1 _20769_ (.A1(_03878_),
    .A2(_03940_),
    .A3(_03941_),
    .B1(_03883_),
    .B2(net5492),
    .X(_01612_));
 sky130_fd_sc_hd__or2_1 _20770_ (.A(net864),
    .B(net5488),
    .X(_03942_));
 sky130_fd_sc_hd__nand2_1 _20771_ (.A(net864),
    .B(net5488),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _20772_ (.A(_03937_),
    .B(_03940_),
    .Y(_03944_));
 sky130_fd_sc_hd__a21o_1 _20773_ (.A1(_03942_),
    .A2(_03943_),
    .B1(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__and3_1 _20774_ (.A(_03942_),
    .B(_03943_),
    .C(_03944_),
    .X(_03946_));
 sky130_fd_sc_hd__inv_2 _20775_ (.A(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__a32o_1 _20776_ (.A1(_03878_),
    .A2(_03945_),
    .A3(_03947_),
    .B1(_03883_),
    .B2(net5488),
    .X(_01613_));
 sky130_fd_sc_hd__or2_1 _20777_ (.A(net1009),
    .B(net5622),
    .X(_03948_));
 sky130_fd_sc_hd__nand2_1 _20778_ (.A(net1009),
    .B(net5622),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_1 _20779_ (.A(_03943_),
    .B(_03947_),
    .Y(_03950_));
 sky130_fd_sc_hd__and3_1 _20780_ (.A(_03948_),
    .B(_03949_),
    .C(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__inv_2 _20781_ (.A(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__a21o_1 _20782_ (.A1(_03948_),
    .A2(_03949_),
    .B1(_03950_),
    .X(_03953_));
 sky130_fd_sc_hd__a32o_1 _20783_ (.A1(_03878_),
    .A2(_03952_),
    .A3(_03953_),
    .B1(_03883_),
    .B2(net5622),
    .X(_01614_));
 sky130_fd_sc_hd__or2_1 _20784_ (.A(net1038),
    .B(net5581),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_1 _20785_ (.A(net1038),
    .B(net5581),
    .Y(_03955_));
 sky130_fd_sc_hd__nand2_1 _20786_ (.A(_03949_),
    .B(_03952_),
    .Y(_03956_));
 sky130_fd_sc_hd__a21o_1 _20787_ (.A1(_03954_),
    .A2(_03955_),
    .B1(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__nand3_1 _20788_ (.A(_03954_),
    .B(_03955_),
    .C(_03956_),
    .Y(_03958_));
 sky130_fd_sc_hd__a32o_1 _20789_ (.A1(_03878_),
    .A2(_03957_),
    .A3(net8209),
    .B1(_03883_),
    .B2(net5581),
    .X(_01615_));
 sky130_fd_sc_hd__a21boi_1 _20790_ (.A1(_03954_),
    .A2(_03956_),
    .B1_N(_03955_),
    .Y(_03959_));
 sky130_fd_sc_hd__nor2_1 _20791_ (.A(net969),
    .B(net5692),
    .Y(_03960_));
 sky130_fd_sc_hd__and2_1 _20792_ (.A(net969),
    .B(net5692),
    .X(_03961_));
 sky130_fd_sc_hd__or3_1 _20793_ (.A(_03959_),
    .B(_03960_),
    .C(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__o21ai_1 _20794_ (.A1(_03960_),
    .A2(_03961_),
    .B1(_03959_),
    .Y(_03963_));
 sky130_fd_sc_hd__a32o_1 _20795_ (.A1(_03878_),
    .A2(_03962_),
    .A3(_03963_),
    .B1(_03883_),
    .B2(net5692),
    .X(_01616_));
 sky130_fd_sc_hd__o21ba_1 _20796_ (.A1(_03959_),
    .A2(_03960_),
    .B1_N(_03961_),
    .X(_03964_));
 sky130_fd_sc_hd__nor2_1 _20797_ (.A(net1015),
    .B(net5522),
    .Y(_03965_));
 sky130_fd_sc_hd__and2_1 _20798_ (.A(net1015),
    .B(net5522),
    .X(_03966_));
 sky130_fd_sc_hd__or3_1 _20799_ (.A(_03964_),
    .B(_03965_),
    .C(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__o21ai_1 _20800_ (.A1(_03965_),
    .A2(_03966_),
    .B1(_03964_),
    .Y(_03968_));
 sky130_fd_sc_hd__a32o_1 _20801_ (.A1(_03878_),
    .A2(_03967_),
    .A3(net8229),
    .B1(_03883_),
    .B2(net5522),
    .X(_01617_));
 sky130_fd_sc_hd__o21ba_1 _20802_ (.A1(_03964_),
    .A2(_03965_),
    .B1_N(_03966_),
    .X(_03969_));
 sky130_fd_sc_hd__nor2_1 _20803_ (.A(net971),
    .B(net5726),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _20804_ (.A(net971),
    .B(net5726),
    .Y(_03971_));
 sky130_fd_sc_hd__and2b_1 _20805_ (.A_N(_03970_),
    .B(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__xnor2_1 _20806_ (.A(_03969_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__a22o_1 _20807_ (.A1(net5726),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03973_),
    .X(_01618_));
 sky130_fd_sc_hd__o21a_1 _20808_ (.A1(_03969_),
    .A2(_03970_),
    .B1(_03971_),
    .X(_03974_));
 sky130_fd_sc_hd__nor2_1 _20809_ (.A(net991),
    .B(net5739),
    .Y(_03975_));
 sky130_fd_sc_hd__and2_1 _20810_ (.A(net991),
    .B(net5739),
    .X(_03976_));
 sky130_fd_sc_hd__nor2_1 _20811_ (.A(_03975_),
    .B(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__xnor2_1 _20812_ (.A(net8222),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__a22o_1 _20813_ (.A1(net5739),
    .A2(_03877_),
    .B1(_03874_),
    .B2(_03978_),
    .X(_01619_));
 sky130_fd_sc_hd__nor2_1 _20814_ (.A(_03974_),
    .B(_03975_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_2 _20815_ (.A(net1028),
    .B(net5480),
    .Y(_03980_));
 sky130_fd_sc_hd__or2_1 _20816_ (.A(net1028),
    .B(net5480),
    .X(_03981_));
 sky130_fd_sc_hd__o211ai_2 _20817_ (.A1(_03976_),
    .A2(_03979_),
    .B1(_03980_),
    .C1(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__a211o_1 _20818_ (.A1(_03981_),
    .A2(_03980_),
    .B1(_03979_),
    .C1(_03976_),
    .X(_03983_));
 sky130_fd_sc_hd__a32o_1 _20819_ (.A1(_09727_),
    .A2(net8200),
    .A3(_03983_),
    .B1(_03689_),
    .B2(net5480),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_1 _20820_ (.A(net850),
    .B(net5609),
    .Y(_03984_));
 sky130_fd_sc_hd__a21oi_1 _20821_ (.A1(_03980_),
    .A2(_03982_),
    .B1(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__a31o_1 _20822_ (.A1(_03980_),
    .A2(_03982_),
    .A3(_03984_),
    .B1(_09720_),
    .X(_03986_));
 sky130_fd_sc_hd__a2bb2o_1 _20823_ (.A1_N(_03985_),
    .A2_N(_03986_),
    .B1(net5609),
    .B2(net63),
    .X(_01621_));
 sky130_fd_sc_hd__o21ai_1 _20824_ (.A1(net4083),
    .A2(net3452),
    .B1(_04485_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_1 _20825_ (.A(_04485_),
    .B(net4122),
    .Y(_03988_));
 sky130_fd_sc_hd__a41o_1 _20826_ (.A1(net3871),
    .A2(net3976),
    .A3(net4083),
    .A4(_03988_),
    .B1(_06237_),
    .X(_03989_));
 sky130_fd_sc_hd__mux2_1 _20827_ (.A0(net4084),
    .A1(_04485_),
    .S(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__and2_1 _20828_ (.A(_08038_),
    .B(net4085),
    .X(_03991_));
 sky130_fd_sc_hd__clkbuf_1 _20829_ (.A(net4086),
    .X(_01622_));
 sky130_fd_sc_hd__o211a_1 _20830_ (.A1(net3628),
    .A2(net5923),
    .B1(_01633_),
    .C1(_04476_),
    .X(_01623_));
 sky130_fd_sc_hd__nor2_1 _20831_ (.A(net3628),
    .B(net5923),
    .Y(_03992_));
 sky130_fd_sc_hd__a21oi_1 _20832_ (.A1(net3976),
    .A2(_03992_),
    .B1(_04490_),
    .Y(_03993_));
 sky130_fd_sc_hd__o21a_1 _20833_ (.A1(net3976),
    .A2(_03992_),
    .B1(_03993_),
    .X(_01624_));
 sky130_fd_sc_hd__a21boi_1 _20834_ (.A1(_04474_),
    .A2(net4083),
    .B1_N(net3871),
    .Y(_03994_));
 sky130_fd_sc_hd__o31a_1 _20835_ (.A1(_09413_),
    .A2(net5923),
    .A3(net3872),
    .B1(_01633_),
    .X(_01625_));
 sky130_fd_sc_hd__and2_2 _20836_ (.A(_03320_),
    .B(clknet_1_0__leaf__05688_),
    .X(_03995_));
 sky130_fd_sc_hd__buf_1 _20837_ (.A(_03995_),
    .X(_01626_));
 sky130_fd_sc_hd__and2_2 _20838_ (.A(_03320_),
    .B(clknet_1_1__leaf__05742_),
    .X(_03996_));
 sky130_fd_sc_hd__buf_1 _20839_ (.A(_03996_),
    .X(_01627_));
 sky130_fd_sc_hd__and2_2 _20840_ (.A(_03320_),
    .B(clknet_1_0__leaf__05794_),
    .X(_03997_));
 sky130_fd_sc_hd__buf_1 _20841_ (.A(_03997_),
    .X(_01628_));
 sky130_fd_sc_hd__and2_2 _20842_ (.A(_09721_),
    .B(clknet_1_0__leaf__05847_),
    .X(_03998_));
 sky130_fd_sc_hd__buf_1 _20843_ (.A(_03998_),
    .X(_01629_));
 sky130_fd_sc_hd__and2_2 _20844_ (.A(_09721_),
    .B(clknet_1_0__leaf__05898_),
    .X(_03999_));
 sky130_fd_sc_hd__buf_1 _20845_ (.A(_03999_),
    .X(_01630_));
 sky130_fd_sc_hd__and2_2 _20846_ (.A(_09721_),
    .B(clknet_1_0__leaf__05946_),
    .X(_04000_));
 sky130_fd_sc_hd__buf_1 _20847_ (.A(_04000_),
    .X(_01631_));
 sky130_fd_sc_hd__nor2_1 _20848_ (.A(net5657),
    .B(net63),
    .Y(_01632_));
 sky130_fd_sc_hd__a22o_1 _20849_ (.A1(net4192),
    .A2(_09745_),
    .B1(_09746_),
    .B2(_09091_),
    .X(_01634_));
 sky130_fd_sc_hd__clkbuf_4 _20850_ (.A(_09736_),
    .X(_04001_));
 sky130_fd_sc_hd__clkbuf_4 _20851_ (.A(_09738_),
    .X(_04002_));
 sky130_fd_sc_hd__a22o_1 _20852_ (.A1(net4206),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_09089_),
    .X(_01635_));
 sky130_fd_sc_hd__a22o_1 _20853_ (.A1(net4202),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_09084_),
    .X(_01636_));
 sky130_fd_sc_hd__a22o_1 _20854_ (.A1(net4211),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_09209_),
    .X(_01637_));
 sky130_fd_sc_hd__a22o_1 _20855_ (.A1(net4213),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_09326_),
    .X(_01638_));
 sky130_fd_sc_hd__a22o_1 _20856_ (.A1(net4215),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_09450_),
    .X(_01639_));
 sky130_fd_sc_hd__a22o_1 _20857_ (.A1(net4219),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_09577_),
    .X(_01640_));
 sky130_fd_sc_hd__a22o_1 _20858_ (.A1(net4224),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_09711_),
    .X(_01641_));
 sky130_fd_sc_hd__a22o_1 _20859_ (.A1(net4229),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_10009_),
    .X(_01642_));
 sky130_fd_sc_hd__a22o_1 _20860_ (.A1(net4217),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_10132_),
    .X(_01643_));
 sky130_fd_sc_hd__a22o_1 _20861_ (.A1(net4204),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_10257_),
    .X(_01644_));
 sky130_fd_sc_hd__nor2_1 _20862_ (.A(net4932),
    .B(net63),
    .Y(_01645_));
 sky130_fd_sc_hd__xnor2_1 _20863_ (.A(net4932),
    .B(net6122),
    .Y(_04003_));
 sky130_fd_sc_hd__nor2_1 _20864_ (.A(_03312_),
    .B(net1093),
    .Y(_01646_));
 sky130_fd_sc_hd__or2_1 _20865_ (.A(net3565),
    .B(net5033),
    .X(_04004_));
 sky130_fd_sc_hd__a32o_1 _20866_ (.A1(_09739_),
    .A2(_02512_),
    .A3(_04004_),
    .B1(_02508_),
    .B2(net5033),
    .X(_01647_));
 sky130_fd_sc_hd__a21bo_1 _20867_ (.A1(_02511_),
    .A2(net4714),
    .B1_N(_02512_),
    .X(_04005_));
 sky130_fd_sc_hd__a32o_1 _20868_ (.A1(_09739_),
    .A2(_02514_),
    .A3(net4715),
    .B1(_02508_),
    .B2(net8105),
    .X(_01648_));
 sky130_fd_sc_hd__or2b_1 _20869_ (.A(_02510_),
    .B_N(_02516_),
    .X(_04006_));
 sky130_fd_sc_hd__xor2_1 _20870_ (.A(_02515_),
    .B(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__a22o_1 _20871_ (.A1(net4887),
    .A2(_02508_),
    .B1(_02559_),
    .B2(_04007_),
    .X(_01649_));
 sky130_fd_sc_hd__and2b_1 _20872_ (.A_N(_02509_),
    .B(_02518_),
    .X(_04008_));
 sky130_fd_sc_hd__xnor2_1 _20873_ (.A(_02517_),
    .B(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__a22o_1 _20874_ (.A1(net4852),
    .A2(_02508_),
    .B1(_02559_),
    .B2(_04009_),
    .X(_01650_));
 sky130_fd_sc_hd__or2_1 _20875_ (.A(net4423),
    .B(net652),
    .X(_04010_));
 sky130_fd_sc_hd__a32o_1 _20876_ (.A1(_09739_),
    .A2(net4424),
    .A3(_04010_),
    .B1(_02508_),
    .B2(net8097),
    .X(_01651_));
 sky130_fd_sc_hd__a21bo_1 _20877_ (.A1(_02753_),
    .A2(net4599),
    .B1_N(net4424),
    .X(_04011_));
 sky130_fd_sc_hd__a32o_1 _20878_ (.A1(_09739_),
    .A2(_02756_),
    .A3(net4600),
    .B1(_02508_),
    .B2(net8100),
    .X(_01652_));
 sky130_fd_sc_hd__or2b_1 _20879_ (.A(_02752_),
    .B_N(_02758_),
    .X(_04012_));
 sky130_fd_sc_hd__xor2_1 _20880_ (.A(_02757_),
    .B(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__a22o_1 _20881_ (.A1(net4879),
    .A2(_02508_),
    .B1(_02559_),
    .B2(net8249),
    .X(_01653_));
 sky130_fd_sc_hd__and2b_1 _20882_ (.A_N(_02751_),
    .B(net4529),
    .X(_04014_));
 sky130_fd_sc_hd__xnor2_1 _20883_ (.A(_02759_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__a22o_1 _20884_ (.A1(net4848),
    .A2(_02508_),
    .B1(_02559_),
    .B2(_04015_),
    .X(_01654_));
 sky130_fd_sc_hd__nor2_1 _20885_ (.A(net4940),
    .B(net63),
    .Y(_01655_));
 sky130_fd_sc_hd__xnor2_1 _20886_ (.A(net4940),
    .B(net6100),
    .Y(_04016_));
 sky130_fd_sc_hd__nor2_1 _20887_ (.A(_03312_),
    .B(net1096),
    .Y(_01656_));
 sky130_fd_sc_hd__nor2_1 _20888_ (.A(net4948),
    .B(net63),
    .Y(_01657_));
 sky130_fd_sc_hd__xnor2_1 _20889_ (.A(net6041),
    .B(net4948),
    .Y(_04017_));
 sky130_fd_sc_hd__nor2_1 _20890_ (.A(_03312_),
    .B(net679),
    .Y(_01658_));
 sky130_fd_sc_hd__nor2_1 _20891_ (.A(net4928),
    .B(net63),
    .Y(_01659_));
 sky130_fd_sc_hd__xnor2_1 _20892_ (.A(net4928),
    .B(net6627),
    .Y(_04018_));
 sky130_fd_sc_hd__nor2_1 _20893_ (.A(_03312_),
    .B(net2614),
    .Y(_01660_));
 sky130_fd_sc_hd__nor2_1 _20894_ (.A(net4936),
    .B(net63),
    .Y(_01661_));
 sky130_fd_sc_hd__xnor2_1 _20895_ (.A(net4936),
    .B(net6111),
    .Y(_04019_));
 sky130_fd_sc_hd__nor2_1 _20896_ (.A(_03312_),
    .B(net1099),
    .Y(_01662_));
 sky130_fd_sc_hd__dfxtp_2 _20897_ (.CLK(clknet_leaf_84_i_clk),
    .D(net5781),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20898_ (.CLK(clknet_4_7__leaf_i_clk),
    .D(net4813),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20899_ (.CLK(clknet_leaf_32_i_clk),
    .D(net5607),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20900_ (.CLK(clknet_leaf_32_i_clk),
    .D(net5533),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20901_ (.CLK(clknet_leaf_37_i_clk),
    .D(net5430),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20902_ (.CLK(clknet_leaf_37_i_clk),
    .D(net5620),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20903_ (.CLK(clknet_leaf_37_i_clk),
    .D(net5410),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20904_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00391_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20905_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00392_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20906_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00393_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20907_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00394_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20908_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00395_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20909_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00396_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20910_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00397_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20911_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00398_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20912_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00399_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20913_ (.CLK(clknet_4_12__leaf_i_clk),
    .D(_00400_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20914_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00401_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20915_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00402_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20916_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00403_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20917_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00404_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20918_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00405_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20919_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20920_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20921_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20922_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20923_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20924_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20925_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20926_ (.CLK(clknet_leaf_60_i_clk),
    .D(net4545),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_2 _20927_ (.CLK(clknet_leaf_75_i_clk),
    .D(net4681),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _20928_ (.CLK(clknet_leaf_60_i_clk),
    .D(net4673),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _20929_ (.CLK(clknet_leaf_60_i_clk),
    .D(net4746),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(clknet_leaf_60_i_clk),
    .D(net4573),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20931_ (.CLK(clknet_leaf_60_i_clk),
    .D(net4549),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20932_ (.CLK(clknet_leaf_80_i_clk),
    .D(net4510),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20933_ (.CLK(clknet_leaf_78_i_clk),
    .D(net4685),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(clknet_leaf_78_i_clk),
    .D(net4732),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20935_ (.CLK(clknet_leaf_78_i_clk),
    .D(net4553),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20936_ (.CLK(clknet_leaf_76_i_clk),
    .D(net4579),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20937_ (.CLK(clknet_leaf_77_i_clk),
    .D(net4587),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20938_ (.CLK(clknet_leaf_77_i_clk),
    .D(net4697),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20939_ (.CLK(clknet_leaf_76_i_clk),
    .D(net4693),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20940_ (.CLK(clknet_leaf_77_i_clk),
    .D(net4740),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20941_ (.CLK(clknet_leaf_77_i_clk),
    .D(net4760),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20942_ (.CLK(clknet_leaf_70_i_clk),
    .D(net4754),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20943_ (.CLK(clknet_leaf_70_i_clk),
    .D(net4721),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20944_ (.CLK(clknet_leaf_70_i_clk),
    .D(net4708),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20945_ (.CLK(clknet_leaf_69_i_clk),
    .D(net4677),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20946_ (.CLK(clknet_leaf_69_i_clk),
    .D(net4663),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20947_ (.CLK(clknet_leaf_77_i_clk),
    .D(net4334),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20948_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20949_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20950_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20951_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20952_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20953_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20954_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20955_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20956_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20957_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20958_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20959_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20960_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20961_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20962_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20963_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20964_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20965_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20966_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20967_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20970_ (.CLK(clknet_leaf_111_i_clk),
    .D(net4158),
    .Q(\reg_rgb[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(clknet_leaf_108_i_clk),
    .D(net4069),
    .Q(\reg_rgb[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(clknet_leaf_111_i_clk),
    .D(net4151),
    .Q(\reg_rgb[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20973_ (.CLK(clknet_leaf_111_i_clk),
    .D(net4143),
    .Q(\reg_rgb[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(clknet_leaf_110_i_clk),
    .D(net4166),
    .Q(\reg_rgb[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_110_i_clk),
    .D(net4175),
    .Q(\reg_rgb[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20976_ (.CLK(clknet_leaf_42_i_clk),
    .D(net3989),
    .Q(\rbzero.wall_hot[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20977_ (.CLK(clknet_leaf_42_i_clk),
    .D(net4014),
    .Q(\rbzero.wall_hot[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(clknet_leaf_81_i_clk),
    .D(net4184),
    .Q(\rbzero.side_hot ));
 sky130_fd_sc_hd__dfxtp_2 _20979_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00466_),
    .Q(\rbzero.texu_hot[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20980_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00467_),
    .Q(\rbzero.texu_hot[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20981_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00468_),
    .Q(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20982_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00469_),
    .Q(\rbzero.texu_hot[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20983_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00470_),
    .Q(\rbzero.texu_hot[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20984_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00471_),
    .Q(\rbzero.texu_hot[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20985_ (.CLK(clknet_leaf_29_i_clk),
    .D(net4125),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3860),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(clknet_leaf_113_i_clk),
    .D(net3958),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_112_i_clk),
    .D(net3920),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_112_i_clk),
    .D(net4060),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_110_i_clk),
    .D(net4109),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_110_i_clk),
    .D(net3518),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20992_ (.CLK(clknet_leaf_111_i_clk),
    .D(net4119),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20993_ (.CLK(clknet_leaf_112_i_clk),
    .D(net4136),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20994_ (.CLK(clknet_leaf_112_i_clk),
    .D(net5951),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20995_ (.CLK(clknet_leaf_52_i_clk),
    .D(net4081),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _20996_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00483_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20997_ (.CLK(clknet_4_15__leaf_i_clk),
    .D(_00484_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20998_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00485_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20999_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00486_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21000_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00487_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21001_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00488_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21002_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00489_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21003_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00490_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21004_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00491_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21005_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00492_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21006_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00493_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21007_ (.CLK(clknet_leaf_37_i_clk),
    .D(net4323),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21008_ (.CLK(clknet_leaf_38_i_clk),
    .D(net4261),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21009_ (.CLK(clknet_leaf_37_i_clk),
    .D(net4337),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21010_ (.CLK(clknet_leaf_38_i_clk),
    .D(net4273),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21011_ (.CLK(clknet_leaf_38_i_clk),
    .D(net1823),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21012_ (.CLK(clknet_leaf_62_i_clk),
    .D(net4289),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21013_ (.CLK(clknet_leaf_62_i_clk),
    .D(net4244),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21014_ (.CLK(clknet_leaf_62_i_clk),
    .D(net4298),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21015_ (.CLK(clknet_leaf_62_i_clk),
    .D(net4320),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21016_ (.CLK(clknet_leaf_59_i_clk),
    .D(net4279),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21017_ (.CLK(clknet_leaf_57_i_clk),
    .D(net4270),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21018_ (.CLK(clknet_leaf_59_i_clk),
    .D(net4238),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(clknet_leaf_57_i_clk),
    .D(net4282),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21020_ (.CLK(clknet_leaf_55_i_clk),
    .D(net4295),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21021_ (.CLK(clknet_leaf_54_i_clk),
    .D(net4241),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21022_ (.CLK(clknet_leaf_63_i_clk),
    .D(net4258),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21023_ (.CLK(clknet_leaf_63_i_clk),
    .D(net4276),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21024_ (.CLK(clknet_leaf_63_i_clk),
    .D(net4301),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21025_ (.CLK(clknet_leaf_53_i_clk),
    .D(net4222),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21026_ (.CLK(clknet_leaf_53_i_clk),
    .D(net4255),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21027_ (.CLK(clknet_leaf_53_i_clk),
    .D(net4264),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21028_ (.CLK(clknet_leaf_53_i_clk),
    .D(net4249),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21029_ (.CLK(clknet_leaf_53_i_clk),
    .D(net4235),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(clknet_leaf_53_i_clk),
    .D(net4227),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21031_ (.CLK(clknet_leaf_55_i_clk),
    .D(net4292),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21032_ (.CLK(clknet_leaf_55_i_clk),
    .D(net4267),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21033_ (.CLK(clknet_leaf_55_i_clk),
    .D(net4252),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21034_ (.CLK(clknet_leaf_34_i_clk),
    .D(net3783),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(clknet_leaf_34_i_clk),
    .D(net3650),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(clknet_leaf_31_i_clk),
    .D(net5556),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21037_ (.CLK(clknet_leaf_56_i_clk),
    .D(net5668),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21038_ (.CLK(clknet_leaf_31_i_clk),
    .D(net5474),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21039_ (.CLK(clknet_leaf_56_i_clk),
    .D(net5724),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21040_ (.CLK(clknet_leaf_56_i_clk),
    .D(net5330),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21041_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00528_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21042_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00529_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21043_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00530_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21044_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00531_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21045_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00532_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21046_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00533_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21047_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00534_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21048_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00535_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21049_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00536_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21050_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00537_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21051_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00538_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21052_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00539_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21053_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00540_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21054_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21055_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21056_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21057_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21058_ (.CLK(clknet_4_13__leaf_i_clk),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21059_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21060_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21061_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21062_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21068_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21071_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21073_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21074_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21080_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21081_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(clknet_leaf_46_i_clk),
    .D(net1288),
    .Q(\rbzero.spi_registers.new_texadd[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(clknet_leaf_46_i_clk),
    .D(net1398),
    .Q(\rbzero.spi_registers.new_texadd[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1424),
    .Q(\rbzero.spi_registers.new_texadd[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21088_ (.CLK(clknet_leaf_13_i_clk),
    .D(net1283),
    .Q(\rbzero.spi_registers.new_texadd[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(clknet_leaf_46_i_clk),
    .D(net1243),
    .Q(\rbzero.spi_registers.new_texadd[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(clknet_leaf_46_i_clk),
    .D(net1421),
    .Q(\rbzero.spi_registers.new_texadd[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21091_ (.CLK(clknet_leaf_47_i_clk),
    .D(net1540),
    .Q(\rbzero.spi_registers.new_texadd[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21092_ (.CLK(clknet_leaf_47_i_clk),
    .D(net1633),
    .Q(\rbzero.spi_registers.new_texadd[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21093_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1510),
    .Q(\rbzero.spi_registers.new_texadd[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1516),
    .Q(\rbzero.spi_registers.new_texadd[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(clknet_leaf_11_i_clk),
    .D(net1437),
    .Q(\rbzero.spi_registers.new_texadd[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(clknet_leaf_11_i_clk),
    .D(net1861),
    .Q(\rbzero.spi_registers.new_texadd[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21097_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1458),
    .Q(\rbzero.spi_registers.new_texadd[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21098_ (.CLK(clknet_leaf_5_i_clk),
    .D(net1679),
    .Q(\rbzero.spi_registers.new_texadd[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21099_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1382),
    .Q(\rbzero.spi_registers.new_texadd[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21100_ (.CLK(clknet_leaf_7_i_clk),
    .D(net1446),
    .Q(\rbzero.spi_registers.new_texadd[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21101_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1373),
    .Q(\rbzero.spi_registers.new_texadd[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21102_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1720),
    .Q(\rbzero.spi_registers.new_texadd[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21103_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1604),
    .Q(\rbzero.spi_registers.new_texadd[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21104_ (.CLK(clknet_leaf_1_i_clk),
    .D(net1449),
    .Q(\rbzero.spi_registers.new_texadd[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21105_ (.CLK(clknet_leaf_4_i_clk),
    .D(net1345),
    .Q(\rbzero.spi_registers.new_texadd[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21106_ (.CLK(clknet_leaf_20_i_clk),
    .D(net1507),
    .Q(\rbzero.spi_registers.new_texadd[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21107_ (.CLK(clknet_leaf_20_i_clk),
    .D(net1601),
    .Q(\rbzero.spi_registers.new_texadd[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21108_ (.CLK(clknet_leaf_17_i_clk),
    .D(net1391),
    .Q(\rbzero.spi_registers.new_texadd[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21109_ (.CLK(clknet_leaf_94_i_clk),
    .D(net4885),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21110_ (.CLK(clknet_leaf_93_i_clk),
    .D(net3143),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21111_ (.CLK(clknet_leaf_94_i_clk),
    .D(net3636),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21112_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3717),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21113_ (.CLK(clknet_leaf_105_i_clk),
    .D(net4787),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21114_ (.CLK(clknet_leaf_105_i_clk),
    .D(net3829),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21115_ (.CLK(clknet_leaf_93_i_clk),
    .D(net4728),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21116_ (.CLK(clknet_leaf_93_i_clk),
    .D(net3606),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21117_ (.CLK(clknet_leaf_92_i_clk),
    .D(net4795),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21118_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3814),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21119_ (.CLK(clknet_leaf_92_i_clk),
    .D(net4823),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21120_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3892),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(clknet_leaf_107_i_clk),
    .D(net4871),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21122_ (.CLK(clknet_leaf_106_i_clk),
    .D(net3736),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(clknet_leaf_92_i_clk),
    .D(net4830),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(clknet_leaf_107_i_clk),
    .D(net3780),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21125_ (.CLK(clknet_leaf_33_i_clk),
    .D(net3895),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(clknet_leaf_33_i_clk),
    .D(net4056),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_1 _21127_ (.CLK(clknet_leaf_33_i_clk),
    .D(net3850),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_1 _21128_ (.CLK(clknet_leaf_33_i_clk),
    .D(net4046),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_1 _21129_ (.CLK(clknet_leaf_32_i_clk),
    .D(net3809),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21130_ (.CLK(clknet_leaf_32_i_clk),
    .D(net3449),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21131_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3963),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(clknet_leaf_29_i_clk),
    .D(net4036),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_1 _21133_ (.CLK(clknet_leaf_29_i_clk),
    .D(net5920),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_1 _21134_ (.CLK(clknet_leaf_31_i_clk),
    .D(net4001),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_1 _21135_ (.CLK(clknet_leaf_29_i_clk),
    .D(net4051),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21136_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3886),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(clknet_leaf_95_i_clk),
    .D(net4533),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21138_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3310),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_4 _21139_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3528),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _21140_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3525),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _21141_ (.CLK(clknet_leaf_99_i_clk),
    .D(net4774),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_4 _21142_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3500),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21143_ (.CLK(clknet_leaf_100_i_clk),
    .D(net4767),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21144_ (.CLK(clknet_leaf_102_i_clk),
    .D(net3754),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21145_ (.CLK(clknet_leaf_104_i_clk),
    .D(net4801),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21146_ (.CLK(clknet_leaf_103_i_clk),
    .D(net3465),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21147_ (.CLK(clknet_leaf_104_i_clk),
    .D(net4810),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21148_ (.CLK(clknet_leaf_103_i_clk),
    .D(net3743),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21149_ (.CLK(clknet_leaf_104_i_clk),
    .D(net4860),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21150_ (.CLK(clknet_leaf_104_i_clk),
    .D(net3603),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21151_ (.CLK(clknet_leaf_106_i_clk),
    .D(net4840),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21152_ (.CLK(clknet_leaf_106_i_clk),
    .D(net3613),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21153_ (.CLK(clknet_leaf_122_i_clk),
    .D(net5847),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21154_ (.CLK(clknet_leaf_23_i_clk),
    .D(net3912),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21155_ (.CLK(clknet_leaf_122_i_clk),
    .D(net5881),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21156_ (.CLK(clknet_leaf_122_i_clk),
    .D(net3938),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21157_ (.CLK(clknet_leaf_2_i_clk),
    .D(net5866),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21158_ (.CLK(clknet_leaf_2_i_clk),
    .D(net5802),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21159_ (.CLK(clknet_4_1__leaf_i_clk),
    .D(net3698),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(clknet_leaf_130_i_clk),
    .D(net3331),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(clknet_leaf_130_i_clk),
    .D(net3353),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21162_ (.CLK(clknet_leaf_130_i_clk),
    .D(net2766),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21163_ (.CLK(clknet_leaf_134_i_clk),
    .D(net1864),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21164_ (.CLK(clknet_leaf_131_i_clk),
    .D(net1575),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(clknet_leaf_132_i_clk),
    .D(net1972),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21166_ (.CLK(clknet_leaf_131_i_clk),
    .D(net1684),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(clknet_leaf_132_i_clk),
    .D(net2470),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3021),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(clknet_leaf_132_i_clk),
    .D(net2958),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(clknet_leaf_132_i_clk),
    .D(net3113),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21171_ (.CLK(clknet_leaf_132_i_clk),
    .D(net2945),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(clknet_leaf_97_i_clk),
    .D(net1196),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21173_ (.CLK(clknet_leaf_97_i_clk),
    .D(net1170),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(clknet_leaf_97_i_clk),
    .D(net2081),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21175_ (.CLK(clknet_leaf_97_i_clk),
    .D(net2163),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21176_ (.CLK(clknet_leaf_97_i_clk),
    .D(net2127),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21177_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1754),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1877),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(clknet_leaf_99_i_clk),
    .D(net2366),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(clknet_leaf_101_i_clk),
    .D(net1948),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(clknet_leaf_128_i_clk),
    .D(net3058),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21182_ (.CLK(clknet_leaf_128_i_clk),
    .D(net3184),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(clknet_leaf_127_i_clk),
    .D(net1224),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21184_ (.CLK(clknet_leaf_101_i_clk),
    .D(net3291),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(clknet_leaf_102_i_clk),
    .D(net2487),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(clknet_leaf_102_i_clk),
    .D(net1917),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3197),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3181),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21189_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3294),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3209),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3278),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3082),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(clknet_leaf_124_i_clk),
    .D(net1246),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(clknet_leaf_126_i_clk),
    .D(net3275),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21195_ (.CLK(clknet_leaf_126_i_clk),
    .D(net1648),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21196_ (.CLK(clknet_leaf_125_i_clk),
    .D(net3364),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(clknet_leaf_126_i_clk),
    .D(net1620),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21198_ (.CLK(clknet_leaf_127_i_clk),
    .D(net1104),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(clknet_leaf_127_i_clk),
    .D(net1934),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(clknet_leaf_127_i_clk),
    .D(net2586),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(clknet_leaf_116_i_clk),
    .D(net3133),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(clknet_leaf_109_i_clk),
    .D(net2332),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(clknet_leaf_109_i_clk),
    .D(net2090),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(clknet_leaf_116_i_clk),
    .D(net2760),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21205_ (.CLK(clknet_leaf_117_i_clk),
    .D(net2840),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21206_ (.CLK(clknet_leaf_117_i_clk),
    .D(net3254),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(clknet_leaf_116_i_clk),
    .D(net1908),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(clknet_leaf_127_i_clk),
    .D(net1147),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21209_ (.CLK(clknet_leaf_117_i_clk),
    .D(net1790),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21210_ (.CLK(clknet_leaf_117_i_clk),
    .D(net2195),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(clknet_leaf_117_i_clk),
    .D(net3325),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21212_ (.CLK(clknet_leaf_118_i_clk),
    .D(net2876),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(clknet_leaf_118_i_clk),
    .D(net2428),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21214_ (.CLK(clknet_leaf_120_i_clk),
    .D(net1560),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21215_ (.CLK(clknet_leaf_120_i_clk),
    .D(net2831),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21216_ (.CLK(clknet_leaf_121_i_clk),
    .D(net3225),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(clknet_leaf_120_i_clk),
    .D(net3040),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_120_i_clk),
    .D(net2942),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_120_i_clk),
    .D(net3100),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21220_ (.CLK(clknet_leaf_119_i_clk),
    .D(net1537),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3413),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3271),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(clknet_leaf_24_i_clk),
    .D(net1473),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_23_i_clk),
    .D(net2865),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21225_ (.CLK(clknet_leaf_23_i_clk),
    .D(net3268),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21226_ (.CLK(clknet_leaf_121_i_clk),
    .D(net1711),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21227_ (.CLK(clknet_leaf_121_i_clk),
    .D(net1705),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_121_i_clk),
    .D(net3281),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(clknet_leaf_123_i_clk),
    .D(net3193),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(clknet_leaf_126_i_clk),
    .D(net1981),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(clknet_leaf_125_i_clk),
    .D(net3017),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(clknet_leaf_123_i_clk),
    .D(net3347),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(clknet_leaf_123_i_clk),
    .D(net1615),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(clknet_leaf_15_i_clk),
    .D(net3901),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00722_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_13_i_clk),
    .D(net4032),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_13_i_clk),
    .D(net4078),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_45_i_clk),
    .D(net4018),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(clknet_leaf_45_i_clk),
    .D(net4042),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(clknet_leaf_44_i_clk),
    .D(net3865),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(clknet_leaf_44_i_clk),
    .D(net3879),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_43_i_clk),
    .D(net3818),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(clknet_leaf_16_i_clk),
    .D(net3404),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(clknet_leaf_11_i_clk),
    .D(net3840),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21245_ (.CLK(clknet_leaf_11_i_clk),
    .D(net3747),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(clknet_leaf_8_i_clk),
    .D(net3400),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21247_ (.CLK(clknet_leaf_21_i_clk),
    .D(net3598),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21248_ (.CLK(clknet_leaf_2_i_clk),
    .D(net3564),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(clknet_leaf_2_i_clk),
    .D(net3740),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3594),
    .Q(\rbzero.spi_registers.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3558),
    .Q(\rbzero.spi_registers.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3676),
    .Q(\rbzero.spi_registers.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(clknet_leaf_1_i_clk),
    .D(net3868),
    .Q(\rbzero.spi_registers.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(clknet_leaf_2_i_clk),
    .D(net3480),
    .Q(\rbzero.spi_registers.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(clknet_leaf_3_i_clk),
    .D(net3483),
    .Q(\rbzero.spi_registers.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(clknet_leaf_2_i_clk),
    .D(net3585),
    .Q(\rbzero.spi_registers.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(clknet_leaf_22_i_clk),
    .D(net3633),
    .Q(\rbzero.spi_registers.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21258_ (.CLK(clknet_leaf_22_i_clk),
    .D(net3795),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21259_ (.CLK(clknet_leaf_22_i_clk),
    .D(net3772),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21260_ (.CLK(clknet_leaf_22_i_clk),
    .D(net3942),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21261_ (.CLK(clknet_leaf_23_i_clk),
    .D(net3853),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21262_ (.CLK(clknet_leaf_122_i_clk),
    .D(net1729),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(clknet_leaf_122_i_clk),
    .D(net2048),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21264_ (.CLK(clknet_leaf_123_i_clk),
    .D(net2437),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(clknet_leaf_122_i_clk),
    .D(net3034),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(clknet_leaf_123_i_clk),
    .D(net2057),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21267_ (.CLK(clknet_leaf_123_i_clk),
    .D(net2184),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(clknet_leaf_122_i_clk),
    .D(net3043),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21269_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5757),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(clknet_leaf_27_i_clk),
    .D(net4311),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(clknet_leaf_27_i_clk),
    .D(net4317),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(clknet_leaf_24_i_clk),
    .D(net4349),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5573),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5529),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21275_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5543),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21276_ (.CLK(clknet_leaf_25_i_clk),
    .D(net4326),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21277_ (.CLK(clknet_leaf_25_i_clk),
    .D(net4308),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21278_ (.CLK(clknet_leaf_27_i_clk),
    .D(net5538),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_25_i_clk),
    .D(net4453),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21280_ (.CLK(clknet_leaf_25_i_clk),
    .D(net4356),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(clknet_leaf_24_i_clk),
    .D(net4371),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(clknet_leaf_24_i_clk),
    .D(net4422),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_24_i_clk),
    .D(net4433),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(clknet_leaf_23_i_clk),
    .D(net5507),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(clknet_leaf_24_i_clk),
    .D(net5434),
    .Q(\rbzero.map_overlay.i_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(clknet_leaf_27_i_clk),
    .D(net5616),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(clknet_leaf_27_i_clk),
    .D(net4368),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_27_i_clk),
    .D(net4395),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_27_i_clk),
    .D(net4386),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(clknet_leaf_26_i_clk),
    .D(net4359),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(clknet_leaf_26_i_clk),
    .D(net5470),
    .Q(\rbzero.map_overlay.i_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(clknet_leaf_34_i_clk),
    .D(net5159),
    .Q(\rbzero.mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21293_ (.CLK(clknet_leaf_34_i_clk),
    .D(net5418),
    .Q(\rbzero.mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21294_ (.CLK(clknet_leaf_34_i_clk),
    .D(net5422),
    .Q(\rbzero.mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5394),
    .Q(\rbzero.mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5095),
    .Q(\rbzero.spi_registers.texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21297_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5055),
    .Q(\rbzero.spi_registers.texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(clknet_leaf_43_i_clk),
    .D(net5238),
    .Q(\rbzero.spi_registers.texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(clknet_leaf_43_i_clk),
    .D(net5007),
    .Q(\rbzero.spi_registers.texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(clknet_leaf_44_i_clk),
    .D(net5083),
    .Q(\rbzero.spi_registers.texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21301_ (.CLK(clknet_leaf_43_i_clk),
    .D(net5187),
    .Q(\rbzero.spi_registers.texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(clknet_leaf_48_i_clk),
    .D(net5366),
    .Q(\rbzero.spi_registers.texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(clknet_leaf_48_i_clk),
    .D(net5258),
    .Q(\rbzero.spi_registers.texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(clknet_leaf_47_i_clk),
    .D(net5242),
    .Q(\rbzero.spi_registers.texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(clknet_leaf_12_i_clk),
    .D(net5326),
    .Q(\rbzero.spi_registers.texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(clknet_leaf_10_i_clk),
    .D(net5214),
    .Q(\rbzero.spi_registers.texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(clknet_leaf_10_i_clk),
    .D(net5294),
    .Q(\rbzero.spi_registers.texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(clknet_leaf_8_i_clk),
    .D(net5246),
    .Q(\rbzero.spi_registers.texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21309_ (.CLK(clknet_leaf_5_i_clk),
    .D(net5374),
    .Q(\rbzero.spi_registers.texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21310_ (.CLK(clknet_leaf_9_i_clk),
    .D(net5123),
    .Q(\rbzero.spi_registers.texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(clknet_leaf_7_i_clk),
    .D(net5234),
    .Q(\rbzero.spi_registers.texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(clknet_leaf_7_i_clk),
    .D(net5067),
    .Q(\rbzero.spi_registers.texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5151),
    .Q(\rbzero.spi_registers.texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(clknet_leaf_3_i_clk),
    .D(net5167),
    .Q(\rbzero.spi_registers.texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(clknet_leaf_3_i_clk),
    .D(net5222),
    .Q(\rbzero.spi_registers.texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5338),
    .Q(\rbzero.spi_registers.texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5350),
    .Q(\rbzero.spi_registers.texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(clknet_leaf_21_i_clk),
    .D(net5438),
    .Q(\rbzero.spi_registers.texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(clknet_leaf_14_i_clk),
    .D(net5446),
    .Q(\rbzero.spi_registers.texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(clknet_leaf_13_i_clk),
    .D(net5266),
    .Q(\rbzero.spi_registers.texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(clknet_leaf_14_i_clk),
    .D(net5334),
    .Q(\rbzero.spi_registers.texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(clknet_leaf_12_i_clk),
    .D(net5127),
    .Q(\rbzero.spi_registers.texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(clknet_leaf_12_i_clk),
    .D(net5354),
    .Q(\rbzero.spi_registers.texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(clknet_leaf_45_i_clk),
    .D(net5099),
    .Q(\rbzero.spi_registers.texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(clknet_leaf_45_i_clk),
    .D(net5143),
    .Q(\rbzero.spi_registers.texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(clknet_leaf_45_i_clk),
    .D(net5230),
    .Q(\rbzero.spi_registers.texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(clknet_leaf_45_i_clk),
    .D(net5031),
    .Q(\rbzero.spi_registers.texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(clknet_leaf_47_i_clk),
    .D(net5079),
    .Q(\rbzero.spi_registers.texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(clknet_leaf_12_i_clk),
    .D(net5063),
    .Q(\rbzero.spi_registers.texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(clknet_leaf_8_i_clk),
    .D(net5390),
    .Q(\rbzero.spi_registers.texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(clknet_leaf_8_i_clk),
    .D(net5426),
    .Q(\rbzero.spi_registers.texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(clknet_leaf_8_i_clk),
    .D(net5147),
    .Q(\rbzero.spi_registers.texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5171),
    .Q(\rbzero.spi_registers.texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(clknet_leaf_9_i_clk),
    .D(net4209),
    .Q(\rbzero.spi_registers.texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5322),
    .Q(\rbzero.spi_registers.texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5286),
    .Q(\rbzero.spi_registers.texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5111),
    .Q(\rbzero.spi_registers.texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5310),
    .Q(\rbzero.spi_registers.texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5414),
    .Q(\rbzero.spi_registers.texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5059),
    .Q(\rbzero.spi_registers.texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5039),
    .Q(\rbzero.spi_registers.texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5370),
    .Q(\rbzero.spi_registers.texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(clknet_leaf_19_i_clk),
    .D(net5091),
    .Q(\rbzero.spi_registers.texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(clknet_leaf_46_i_clk),
    .D(net5131),
    .Q(\rbzero.spi_registers.texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(clknet_leaf_13_i_clk),
    .D(net4200),
    .Q(\rbzero.spi_registers.texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(clknet_leaf_13_i_clk),
    .D(net5163),
    .Q(\rbzero.spi_registers.texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(clknet_leaf_13_i_clk),
    .D(net5270),
    .Q(\rbzero.spi_registers.texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(clknet_leaf_45_i_clk),
    .D(net5203),
    .Q(\rbzero.spi_registers.texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(clknet_leaf_45_i_clk),
    .D(net5218),
    .Q(\rbzero.spi_registers.texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(clknet_leaf_47_i_clk),
    .D(net5119),
    .Q(\rbzero.spi_registers.texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(clknet_leaf_47_i_clk),
    .D(net5298),
    .Q(\rbzero.spi_registers.texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(clknet_leaf_47_i_clk),
    .D(net5075),
    .Q(\rbzero.spi_registers.texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(clknet_leaf_12_i_clk),
    .D(net5139),
    .Q(\rbzero.spi_registers.texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(clknet_leaf_10_i_clk),
    .D(net5262),
    .Q(\rbzero.spi_registers.texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(clknet_leaf_10_i_clk),
    .D(net5087),
    .Q(\rbzero.spi_registers.texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(clknet_leaf_8_i_clk),
    .D(net5302),
    .Q(\rbzero.spi_registers.texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(clknet_leaf_5_i_clk),
    .D(net5318),
    .Q(\rbzero.spi_registers.texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(clknet_leaf_14_i_clk),
    .D(net5458),
    .Q(\rbzero.spi_registers.texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(clknet_leaf_7_i_clk),
    .D(net5179),
    .Q(\rbzero.spi_registers.texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5183),
    .Q(\rbzero.spi_registers.texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5278),
    .Q(\rbzero.spi_registers.texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(clknet_leaf_3_i_clk),
    .D(net5135),
    .Q(\rbzero.spi_registers.texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4197),
    .Q(\rbzero.spi_registers.texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5015),
    .Q(\rbzero.spi_registers.texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5071),
    .Q(\rbzero.spi_registers.texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5306),
    .Q(\rbzero.spi_registers.texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(clknet_leaf_18_i_clk),
    .D(net5346),
    .Q(\rbzero.spi_registers.texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(clknet_leaf_14_i_clk),
    .D(net5019),
    .Q(\rbzero.spi_registers.texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(clknet_leaf_14_i_clk),
    .D(net5043),
    .Q(\rbzero.spi_registers.texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(clknet_leaf_10_i_clk),
    .D(net5195),
    .Q(\rbzero.spi_registers.texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(clknet_leaf_10_i_clk),
    .D(net4994),
    .Q(\rbzero.spi_registers.texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(clknet_leaf_44_i_clk),
    .D(net5115),
    .Q(\rbzero.spi_registers.texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(clknet_leaf_44_i_clk),
    .D(net5362),
    .Q(\rbzero.spi_registers.texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(clknet_leaf_48_i_clk),
    .D(net5398),
    .Q(\rbzero.spi_registers.texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(clknet_leaf_45_i_clk),
    .D(net5314),
    .Q(\rbzero.spi_registers.texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(clknet_leaf_46_i_clk),
    .D(net5107),
    .Q(\rbzero.spi_registers.texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(clknet_leaf_12_i_clk),
    .D(net5290),
    .Q(\rbzero.spi_registers.texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(clknet_leaf_9_i_clk),
    .D(net5023),
    .Q(\rbzero.spi_registers.texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(clknet_leaf_9_i_clk),
    .D(net5011),
    .Q(\rbzero.spi_registers.texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(clknet_leaf_9_i_clk),
    .D(net5027),
    .Q(\rbzero.spi_registers.texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(clknet_leaf_3_i_clk),
    .D(net5003),
    .Q(\rbzero.spi_registers.texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(clknet_leaf_9_i_clk),
    .D(net5103),
    .Q(\rbzero.spi_registers.texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5226),
    .Q(\rbzero.spi_registers.texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5155),
    .Q(\rbzero.spi_registers.texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(clknet_leaf_6_i_clk),
    .D(net5175),
    .Q(\rbzero.spi_registers.texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(clknet_leaf_3_i_clk),
    .D(net5191),
    .Q(\rbzero.spi_registers.texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(clknet_leaf_3_i_clk),
    .D(net5199),
    .Q(\rbzero.spi_registers.texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(clknet_leaf_20_i_clk),
    .D(net4990),
    .Q(\rbzero.spi_registers.texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5250),
    .Q(\rbzero.spi_registers.texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(clknet_leaf_21_i_clk),
    .D(net5274),
    .Q(\rbzero.spi_registers.texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(clknet_leaf_19_i_clk),
    .D(net4978),
    .Q(\rbzero.spi_registers.texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(clknet_leaf_39_i_clk),
    .D(net5442),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(clknet_leaf_39_i_clk),
    .D(net5462),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(clknet_leaf_39_i_clk),
    .D(net5486),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(clknet_leaf_39_i_clk),
    .D(net5503),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(clknet_leaf_39_i_clk),
    .D(net5520),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(clknet_leaf_39_i_clk),
    .D(net5511),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(clknet_leaf_41_i_clk),
    .D(net5358),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(clknet_leaf_41_i_clk),
    .D(net3572),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(clknet_leaf_41_i_clk),
    .D(net4966),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(clknet_leaf_41_i_clk),
    .D(net3673),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(clknet_leaf_41_i_clk),
    .D(net5051),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(clknet_leaf_41_i_clk),
    .D(net3654),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(clknet_leaf_36_i_clk),
    .D(net3659),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(clknet_leaf_35_i_clk),
    .D(net4962),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(clknet_leaf_36_i_clk),
    .D(net3550),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(clknet_leaf_35_i_clk),
    .D(net4954),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(clknet_leaf_36_i_clk),
    .D(net3647),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21409_ (.CLK(clknet_leaf_36_i_clk),
    .D(net4958),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21410_ (.CLK(clknet_leaf_38_i_clk),
    .D(net4314),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21411_ (.CLK(clknet_leaf_38_i_clk),
    .D(net5516),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21412_ (.CLK(clknet_leaf_38_i_clk),
    .D(net5565),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21413_ (.CLK(clknet_leaf_38_i_clk),
    .D(net4232),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(clknet_leaf_52_i_clk),
    .D(net5466),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(clknet_leaf_38_i_clk),
    .D(net5454),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21416_ (.CLK(clknet_leaf_2_i_clk),
    .D(net3908),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(clknet_leaf_41_i_clk),
    .D(net1735),
    .Q(\rbzero.spi_registers.new_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(clknet_leaf_42_i_clk),
    .D(net1534),
    .Q(\rbzero.spi_registers.new_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21419_ (.CLK(clknet_leaf_40_i_clk),
    .D(net2323),
    .Q(\rbzero.spi_registers.new_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(clknet_leaf_41_i_clk),
    .D(net1726),
    .Q(\rbzero.spi_registers.new_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(clknet_leaf_41_i_clk),
    .D(net2443),
    .Q(\rbzero.spi_registers.new_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(clknet_leaf_41_i_clk),
    .D(net2062),
    .Q(\rbzero.spi_registers.new_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(clknet_leaf_18_i_clk),
    .D(net3904),
    .Q(\rbzero.spi_registers.got_new_sky ));
 sky130_fd_sc_hd__dfxtp_1 _21424_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1482),
    .Q(\rbzero.spi_registers.new_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21425_ (.CLK(clknet_leaf_35_i_clk),
    .D(net1595),
    .Q(\rbzero.spi_registers.new_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(clknet_leaf_40_i_clk),
    .D(net1566),
    .Q(\rbzero.spi_registers.new_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(clknet_leaf_35_i_clk),
    .D(net1627),
    .Q(\rbzero.spi_registers.new_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(clknet_leaf_36_i_clk),
    .D(net2234),
    .Q(\rbzero.spi_registers.new_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1563),
    .Q(\rbzero.spi_registers.new_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(clknet_leaf_26_i_clk),
    .D(net3522),
    .Q(\rbzero.spi_registers.got_new_floor ));
 sky130_fd_sc_hd__dfxtp_1 _21431_ (.CLK(clknet_leaf_40_i_clk),
    .D(net2449),
    .Q(\rbzero.spi_registers.new_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21432_ (.CLK(clknet_leaf_40_i_clk),
    .D(net1645),
    .Q(\rbzero.spi_registers.new_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21433_ (.CLK(clknet_leaf_40_i_clk),
    .D(net2258),
    .Q(\rbzero.spi_registers.new_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21434_ (.CLK(clknet_leaf_40_i_clk),
    .D(net1636),
    .Q(\rbzero.spi_registers.new_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(clknet_leaf_40_i_clk),
    .D(net1673),
    .Q(\rbzero.spi_registers.new_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21436_ (.CLK(clknet_leaf_40_i_clk),
    .D(net2148),
    .Q(\rbzero.spi_registers.new_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21437_ (.CLK(clknet_leaf_18_i_clk),
    .D(net3219),
    .Q(\rbzero.spi_registers.got_new_leak ));
 sky130_fd_sc_hd__dfxtp_1 _21438_ (.CLK(clknet_leaf_25_i_clk),
    .D(net1642),
    .Q(\rbzero.spi_registers.new_other[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(clknet_leaf_25_i_clk),
    .D(net1738),
    .Q(\rbzero.spi_registers.new_other[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21440_ (.CLK(clknet_leaf_26_i_clk),
    .D(net1495),
    .Q(\rbzero.spi_registers.new_other[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21441_ (.CLK(clknet_leaf_26_i_clk),
    .D(net1428),
    .Q(\rbzero.spi_registers.new_other[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(clknet_leaf_26_i_clk),
    .D(net1702),
    .Q(\rbzero.spi_registers.new_other[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(clknet_leaf_17_i_clk),
    .D(net3369),
    .Q(\rbzero.spi_registers.new_other[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(clknet_leaf_18_i_clk),
    .D(net3335),
    .Q(\rbzero.spi_registers.new_other[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(clknet_leaf_17_i_clk),
    .D(net3088),
    .Q(\rbzero.spi_registers.new_other[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(clknet_leaf_19_i_clk),
    .D(net2955),
    .Q(\rbzero.spi_registers.new_other[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21447_ (.CLK(clknet_leaf_25_i_clk),
    .D(net1766),
    .Q(\rbzero.spi_registers.new_other[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(clknet_leaf_19_i_clk),
    .D(net3625),
    .Q(\rbzero.spi_registers.got_new_other ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(clknet_leaf_39_i_clk),
    .D(net1624),
    .Q(\rbzero.spi_registers.new_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21450_ (.CLK(clknet_leaf_38_i_clk),
    .D(net1584),
    .Q(\rbzero.spi_registers.new_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1404),
    .Q(\rbzero.spi_registers.new_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(clknet_leaf_39_i_clk),
    .D(net2100),
    .Q(\rbzero.spi_registers.new_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1744),
    .Q(\rbzero.spi_registers.new_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(clknet_leaf_39_i_clk),
    .D(net2225),
    .Q(\rbzero.spi_registers.new_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(clknet_leaf_26_i_clk),
    .D(net3981),
    .Q(\rbzero.spi_registers.got_new_vshift ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(clknet_leaf_19_i_clk),
    .D(net1884),
    .Q(\rbzero.spi_registers.new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(clknet_leaf_25_i_clk),
    .D(net3377),
    .Q(\rbzero.spi_registers.got_new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(clknet_leaf_42_i_clk),
    .D(net1431),
    .Q(\rbzero.spi_registers.new_mapd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(clknet_leaf_42_i_clk),
    .D(net1999),
    .Q(\rbzero.spi_registers.new_mapd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21460_ (.CLK(clknet_leaf_41_i_clk),
    .D(net1321),
    .Q(\rbzero.spi_registers.new_mapd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21461_ (.CLK(clknet_leaf_42_i_clk),
    .D(net3004),
    .Q(\rbzero.spi_registers.new_mapd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21462_ (.CLK(clknet_leaf_18_i_clk),
    .D(net2106),
    .Q(\rbzero.spi_registers.new_mapd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21463_ (.CLK(clknet_leaf_42_i_clk),
    .D(net2207),
    .Q(\rbzero.spi_registers.new_mapd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(clknet_leaf_17_i_clk),
    .D(net2646),
    .Q(\rbzero.spi_registers.new_mapd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21465_ (.CLK(clknet_leaf_17_i_clk),
    .D(net2600),
    .Q(\rbzero.spi_registers.new_mapd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(clknet_leaf_42_i_clk),
    .D(net2005),
    .Q(\rbzero.spi_registers.new_mapd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(clknet_leaf_18_i_clk),
    .D(net1294),
    .Q(\rbzero.spi_registers.new_mapd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21468_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1479),
    .Q(\rbzero.spi_registers.new_mapd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21469_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1394),
    .Q(\rbzero.spi_registers.new_mapd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21470_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1543),
    .Q(\rbzero.spi_registers.new_mapd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1657),
    .Q(\rbzero.spi_registers.new_mapd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21472_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1781),
    .Q(\rbzero.spi_registers.new_mapd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21473_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1639),
    .Q(\rbzero.spi_registers.new_mapd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21474_ (.CLK(clknet_leaf_18_i_clk),
    .D(net888),
    .Q(\rbzero.spi_registers.got_new_mapd ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(clknet_leaf_21_i_clk),
    .D(net3845),
    .Q(\rbzero.spi_registers.got_new_texadd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21476_ (.CLK(clknet_leaf_18_i_clk),
    .D(net4837),
    .Q(\rbzero.spi_registers.got_new_texadd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(clknet_leaf_18_i_clk),
    .D(net4846),
    .Q(\rbzero.spi_registers.got_new_texadd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(clknet_leaf_19_i_clk),
    .D(net4818),
    .Q(\rbzero.spi_registers.got_new_texadd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(clknet_leaf_15_i_clk),
    .D(net1303),
    .Q(\rbzero.spi_registers.new_texadd[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(clknet_leaf_16_i_clk),
    .D(net1379),
    .Q(\rbzero.spi_registers.new_texadd[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(clknet_leaf_43_i_clk),
    .D(net1213),
    .Q(\rbzero.spi_registers.new_texadd[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(clknet_leaf_43_i_clk),
    .D(net1249),
    .Q(\rbzero.spi_registers.new_texadd[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21483_ (.CLK(clknet_leaf_44_i_clk),
    .D(net1546),
    .Q(\rbzero.spi_registers.new_texadd[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(clknet_leaf_44_i_clk),
    .D(net1376),
    .Q(\rbzero.spi_registers.new_texadd[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(clknet_leaf_48_i_clk),
    .D(net1297),
    .Q(\rbzero.spi_registers.new_texadd[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21486_ (.CLK(clknet_leaf_48_i_clk),
    .D(net1670),
    .Q(\rbzero.spi_registers.new_texadd[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(clknet_leaf_47_i_clk),
    .D(net1280),
    .Q(\rbzero.spi_registers.new_texadd[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21488_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1630),
    .Q(\rbzero.spi_registers.new_texadd[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21489_ (.CLK(clknet_leaf_11_i_clk),
    .D(net1470),
    .Q(\rbzero.spi_registers.new_texadd[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21490_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1925),
    .Q(\rbzero.spi_registers.new_texadd[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21491_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1485),
    .Q(\rbzero.spi_registers.new_texadd[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21492_ (.CLK(clknet_leaf_5_i_clk),
    .D(net1407),
    .Q(\rbzero.spi_registers.new_texadd[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21493_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1772),
    .Q(\rbzero.spi_registers.new_texadd[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(clknet_leaf_7_i_clk),
    .D(net1813),
    .Q(\rbzero.spi_registers.new_texadd[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21495_ (.CLK(clknet_leaf_7_i_clk),
    .D(net1330),
    .Q(\rbzero.spi_registers.new_texadd[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21496_ (.CLK(clknet_leaf_0_i_clk),
    .D(net2270),
    .Q(\rbzero.spi_registers.new_texadd[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21497_ (.CLK(clknet_leaf_1_i_clk),
    .D(net1905),
    .Q(\rbzero.spi_registers.new_texadd[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21498_ (.CLK(clknet_leaf_3_i_clk),
    .D(net1572),
    .Q(\rbzero.spi_registers.new_texadd[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21499_ (.CLK(clknet_leaf_3_i_clk),
    .D(net1333),
    .Q(\rbzero.spi_registers.new_texadd[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21500_ (.CLK(clknet_leaf_3_i_clk),
    .D(net1651),
    .Q(\rbzero.spi_registers.new_texadd[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21501_ (.CLK(clknet_leaf_22_i_clk),
    .D(net1434),
    .Q(\rbzero.spi_registers.new_texadd[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21502_ (.CLK(clknet_leaf_15_i_clk),
    .D(net1268),
    .Q(\rbzero.spi_registers.new_texadd[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21503_ (.CLK(clknet_leaf_13_i_clk),
    .D(net1309),
    .Q(\rbzero.spi_registers.new_texadd[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21504_ (.CLK(clknet_leaf_14_i_clk),
    .D(net1312),
    .Q(\rbzero.spi_registers.new_texadd[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1339),
    .Q(\rbzero.spi_registers.new_texadd[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21506_ (.CLK(clknet_leaf_11_i_clk),
    .D(net1696),
    .Q(\rbzero.spi_registers.new_texadd[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(clknet_leaf_45_i_clk),
    .D(net1348),
    .Q(\rbzero.spi_registers.new_texadd[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(clknet_leaf_45_i_clk),
    .D(net1418),
    .Q(\rbzero.spi_registers.new_texadd[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(clknet_leaf_48_i_clk),
    .D(net1693),
    .Q(\rbzero.spi_registers.new_texadd[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21510_ (.CLK(clknet_leaf_48_i_clk),
    .D(net1802),
    .Q(\rbzero.spi_registers.new_texadd[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21511_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1554),
    .Q(\rbzero.spi_registers.new_texadd[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21512_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1513),
    .Q(\rbzero.spi_registers.new_texadd[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21513_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1491),
    .Q(\rbzero.spi_registers.new_texadd[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21514_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1351),
    .Q(\rbzero.spi_registers.new_texadd[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21515_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1455),
    .Q(\rbzero.spi_registers.new_texadd[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21516_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1464),
    .Q(\rbzero.spi_registers.new_texadd[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21517_ (.CLK(clknet_leaf_5_i_clk),
    .D(net1336),
    .Q(\rbzero.spi_registers.new_texadd[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21518_ (.CLK(clknet_leaf_7_i_clk),
    .D(net1498),
    .Q(\rbzero.spi_registers.new_texadd[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(clknet_leaf_7_i_clk),
    .D(net1327),
    .Q(\rbzero.spi_registers.new_texadd[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1699),
    .Q(\rbzero.spi_registers.new_texadd[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21521_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1747),
    .Q(\rbzero.spi_registers.new_texadd[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21522_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1667),
    .Q(\rbzero.spi_registers.new_texadd[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21523_ (.CLK(clknet_leaf_3_i_clk),
    .D(net2077),
    .Q(\rbzero.spi_registers.new_texadd[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21524_ (.CLK(clknet_leaf_3_i_clk),
    .D(net2416),
    .Q(\rbzero.spi_registers.new_texadd[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(clknet_leaf_20_i_clk),
    .D(net2139),
    .Q(\rbzero.spi_registers.new_texadd[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(clknet_leaf_19_i_clk),
    .D(net1525),
    .Q(\rbzero.spi_registers.new_texadd[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(clknet_leaf_119_i_clk),
    .D(net4999),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _21528_ (.CLK(clknet_leaf_124_i_clk),
    .D(net5282),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21529_ (.CLK(clknet_leaf_124_i_clk),
    .D(net3706),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(clknet_leaf_135_i_clk),
    .D(net5498),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21531_ (.CLK(clknet_leaf_135_i_clk),
    .D(net3710),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21532_ (.CLK(clknet_leaf_130_i_clk),
    .D(net3924),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(clknet_leaf_130_i_clk),
    .D(net3826),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21534_ (.CLK(clknet_leaf_130_i_clk),
    .D(net4946),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21535_ (.CLK(net169),
    .D(net1838),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(net170),
    .D(net2837),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21537_ (.CLK(net171),
    .D(net2897),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(net172),
    .D(net2166),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21539_ (.CLK(net173),
    .D(net1945),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(net174),
    .D(net2317),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21541_ (.CLK(net175),
    .D(net3007),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21542_ (.CLK(net176),
    .D(net2834),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21543_ (.CLK(net177),
    .D(net2074),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(net178),
    .D(net1150),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21545_ (.CLK(net179),
    .D(net2894),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21546_ (.CLK(net180),
    .D(net2913),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(net181),
    .D(net1911),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21548_ (.CLK(net182),
    .D(net2172),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(net183),
    .D(net1723),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21550_ (.CLK(net184),
    .D(net2347),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(net185),
    .D(net1954),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21552_ (.CLK(net186),
    .D(net2919),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21553_ (.CLK(net187),
    .D(net2681),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21554_ (.CLK(net188),
    .D(net635),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(net189),
    .D(net1826),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21556_ (.CLK(net190),
    .D(net2481),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21557_ (.CLK(net191),
    .D(net2856),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21558_ (.CLK(net192),
    .D(net1760),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21559_ (.CLK(net193),
    .D(net1732),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(net194),
    .D(net2609),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(net195),
    .D(net2964),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(net196),
    .D(net2529),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(net197),
    .D(net1899),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(net198),
    .D(net906),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(net199),
    .D(net2458),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21566_ (.CLK(net200),
    .D(net2746),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(net201),
    .D(net1775),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21568_ (.CLK(net202),
    .D(net1714),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(net203),
    .D(net2727),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(net204),
    .D(net2843),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(net205),
    .D(net2213),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21572_ (.CLK(net206),
    .D(net2383),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(net207),
    .D(net1931),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(net208),
    .D(net1054),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(net209),
    .D(net2675),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(net210),
    .D(net2815),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21577_ (.CLK(net211),
    .D(net2656),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21578_ (.CLK(net212),
    .D(net2806),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21579_ (.CLK(net213),
    .D(net1984),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(net214),
    .D(net1199),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21581_ (.CLK(net215),
    .D(net3119),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21582_ (.CLK(net216),
    .D(net2490),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(net217),
    .D(net2574),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21584_ (.CLK(net218),
    .D(net940),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21585_ (.CLK(net219),
    .D(net2541),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21586_ (.CLK(net220),
    .D(net2389),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21587_ (.CLK(net221),
    .D(net2169),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21588_ (.CLK(net222),
    .D(net2989),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21589_ (.CLK(net223),
    .D(net1501),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21590_ (.CLK(net224),
    .D(net2514),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21591_ (.CLK(net225),
    .D(net1821),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(net226),
    .D(net1763),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21593_ (.CLK(net227),
    .D(net2281),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21594_ (.CLK(net228),
    .D(net625),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(net229),
    .D(net2650),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21596_ (.CLK(net230),
    .D(net2362),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21597_ (.CLK(net231),
    .D(net2084),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(net232),
    .D(net1969),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21599_ (.CLK(clknet_leaf_130_i_clk),
    .D(net1816),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21600_ (.CLK(clknet_leaf_130_i_clk),
    .D(net3212),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21601_ (.CLK(clknet_leaf_130_i_clk),
    .D(net3232),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21602_ (.CLK(clknet_leaf_134_i_clk),
    .D(net2508),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21603_ (.CLK(clknet_leaf_134_i_clk),
    .D(net3047),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21604_ (.CLK(clknet_leaf_131_i_clk),
    .D(net1318),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21605_ (.CLK(clknet_leaf_130_i_clk),
    .D(net1581),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21606_ (.CLK(clknet_leaf_131_i_clk),
    .D(net2264),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(clknet_leaf_131_i_clk),
    .D(net3028),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(clknet_leaf_132_i_clk),
    .D(net1858),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21609_ (.CLK(clknet_leaf_132_i_clk),
    .D(net3147),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(clknet_leaf_132_i_clk),
    .D(net3103),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(clknet_leaf_133_i_clk),
    .D(net2871),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(clknet_leaf_133_i_clk),
    .D(net2773),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(clknet_leaf_97_i_clk),
    .D(net1184),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21614_ (.CLK(clknet_leaf_97_i_clk),
    .D(net2809),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(clknet_leaf_97_i_clk),
    .D(net3079),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(clknet_leaf_97_i_clk),
    .D(net3065),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1708),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21618_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3157),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21619_ (.CLK(clknet_leaf_128_i_clk),
    .D(net737),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_128_i_clk),
    .D(net3188),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_128_i_clk),
    .D(net2922),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_128_i_clk),
    .D(net3024),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_101_i_clk),
    .D(net2181),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_101_i_clk),
    .D(net3175),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_128_i_clk),
    .D(net1690),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21626_ (.CLK(clknet_leaf_127_i_clk),
    .D(net1232),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3150),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3344),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21629_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3304),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21630_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3235),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21631_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3258),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21632_ (.CLK(clknet_leaf_129_i_clk),
    .D(net3075),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_124_i_clk),
    .D(net1360),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21634_ (.CLK(clknet_leaf_125_i_clk),
    .D(net3300),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21635_ (.CLK(clknet_leaf_125_i_clk),
    .D(net3097),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21636_ (.CLK(clknet_leaf_125_i_clk),
    .D(net3127),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21637_ (.CLK(clknet_leaf_125_i_clk),
    .D(net2936),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21638_ (.CLK(clknet_leaf_127_i_clk),
    .D(net1153),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3322),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21640_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3216),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21641_ (.CLK(clknet_leaf_116_i_clk),
    .D(net3168),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21642_ (.CLK(clknet_leaf_116_i_clk),
    .D(net3262),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21643_ (.CLK(clknet_leaf_116_i_clk),
    .D(net2976),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(clknet_leaf_117_i_clk),
    .D(net2071),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21645_ (.CLK(clknet_leaf_117_i_clk),
    .D(net3140),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21646_ (.CLK(clknet_leaf_117_i_clk),
    .D(net3136),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21647_ (.CLK(clknet_leaf_126_i_clk),
    .D(net1887),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21648_ (.CLK(clknet_leaf_126_i_clk),
    .D(net2803),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21649_ (.CLK(clknet_leaf_126_i_clk),
    .D(net3229),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21650_ (.CLK(clknet_leaf_117_i_clk),
    .D(net2413),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21651_ (.CLK(clknet_leaf_118_i_clk),
    .D(net3054),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(clknet_leaf_118_i_clk),
    .D(net2544),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(clknet_leaf_121_i_clk),
    .D(net1112),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(clknet_leaf_121_i_clk),
    .D(net3123),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21655_ (.CLK(clknet_leaf_121_i_clk),
    .D(net3314),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(clknet_leaf_121_i_clk),
    .D(net3285),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(clknet_leaf_121_i_clk),
    .D(net2862),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(clknet_leaf_121_i_clk),
    .D(net3062),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21659_ (.CLK(clknet_leaf_120_i_clk),
    .D(net2905),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_24_i_clk),
    .D(net1167),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3288),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(clknet_leaf_23_i_clk),
    .D(net2714),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_23_i_clk),
    .D(net3161),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(clknet_leaf_23_i_clk),
    .D(net2929),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_122_i_clk),
    .D(net2192),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(clknet_leaf_122_i_clk),
    .D(net3011),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21667_ (.CLK(clknet_leaf_121_i_clk),
    .D(net1569),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(clknet_leaf_123_i_clk),
    .D(net589),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21669_ (.CLK(clknet_leaf_123_i_clk),
    .D(net3239),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21670_ (.CLK(clknet_leaf_125_i_clk),
    .D(net2314),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21671_ (.CLK(clknet_leaf_123_i_clk),
    .D(net1262),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21672_ (.CLK(clknet_leaf_123_i_clk),
    .D(net1871),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21673_ (.CLK(clknet_leaf_124_i_clk),
    .D(net1868),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21674_ (.CLK(clknet_leaf_124_i_clk),
    .D(net1810),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21675_ (.CLK(clknet_leaf_124_i_clk),
    .D(net3201),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(clknet_leaf_124_i_clk),
    .D(net3050),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21677_ (.CLK(clknet_leaf_124_i_clk),
    .D(net2891),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(clknet_leaf_124_i_clk),
    .D(net3222),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(clknet_leaf_124_i_clk),
    .D(net3307),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(clknet_leaf_114_i_clk),
    .D(net5748),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(clknet_leaf_113_i_clk),
    .D(net5820),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21682_ (.CLK(clknet_leaf_113_i_clk),
    .D(net5839),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(clknet_leaf_114_i_clk),
    .D(net5889),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(clknet_leaf_114_i_clk),
    .D(net3546),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21685_ (.CLK(clknet_leaf_115_i_clk),
    .D(net4445),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21686_ (.CLK(clknet_leaf_115_i_clk),
    .D(net5853),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21687_ (.CLK(clknet_leaf_115_i_clk),
    .D(net4494),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(clknet_leaf_114_i_clk),
    .D(net5829),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21689_ (.CLK(clknet_leaf_28_i_clk),
    .D(net5871),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21690_ (.CLK(clknet_leaf_28_i_clk),
    .D(net3994),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21691_ (.CLK(clknet_leaf_114_i_clk),
    .D(net4457),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(clknet_leaf_114_i_clk),
    .D(net5901),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21693_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3685),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21694_ (.CLK(clknet_leaf_24_i_clk),
    .D(net4022),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21695_ (.CLK(clknet_leaf_110_i_clk),
    .D(net3442),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21696_ (.CLK(clknet_leaf_115_i_clk),
    .D(net4620),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(clknet_leaf_115_i_clk),
    .D(net5861),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21698_ (.CLK(clknet_leaf_116_i_clk),
    .D(net5753),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21699_ (.CLK(clknet_leaf_116_i_clk),
    .D(net4346),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(clknet_leaf_115_i_clk),
    .D(net4365),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(clknet_leaf_115_i_clk),
    .D(net4330),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21702_ (.CLK(clknet_leaf_118_i_clk),
    .D(net5774),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21703_ (.CLK(clknet_leaf_119_i_clk),
    .D(net4286),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21704_ (.CLK(clknet_leaf_118_i_clk),
    .D(net4904),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21705_ (.CLK(clknet_leaf_118_i_clk),
    .D(net4750),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21706_ (.CLK(clknet_leaf_118_i_clk),
    .D(net4438),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21707_ (.CLK(clknet_leaf_119_i_clk),
    .D(net4377),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21708_ (.CLK(clknet_leaf_119_i_clk),
    .D(net3555),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21709_ (.CLK(clknet_leaf_119_i_clk),
    .D(net3471),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21710_ (.CLK(clknet_leaf_109_i_clk),
    .D(net4628),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21711_ (.CLK(clknet_leaf_109_i_clk),
    .D(net4479),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21712_ (.CLK(clknet_leaf_103_i_clk),
    .D(net4475),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21713_ (.CLK(clknet_leaf_103_i_clk),
    .D(net4465),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21714_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3438),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21715_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3693),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21716_ (.CLK(clknet_leaf_127_i_clk),
    .D(net3610),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21717_ (.CLK(clknet_leaf_103_i_clk),
    .D(net4597),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21718_ (.CLK(clknet_leaf_109_i_clk),
    .D(net3722),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21719_ (.CLK(clknet_leaf_109_i_clk),
    .D(net4516),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21720_ (.CLK(clknet_leaf_109_i_clk),
    .D(net4449),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21721_ (.CLK(clknet_leaf_100_i_clk),
    .D(net3689),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_4 _21722_ (.CLK(clknet_leaf_102_i_clk),
    .D(net4411),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21723_ (.CLK(clknet_leaf_103_i_clk),
    .D(net3506),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21724_ (.CLK(clknet_leaf_103_i_clk),
    .D(net3582),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21725_ (.CLK(clknet_leaf_110_i_clk),
    .D(net3883),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21726_ (.CLK(clknet_leaf_102_i_clk),
    .D(net4469),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21727_ (.CLK(clknet_leaf_102_i_clk),
    .D(net4489),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(clknet_leaf_103_i_clk),
    .D(net3714),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(clknet_leaf_101_i_clk),
    .D(net4419),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(clknet_leaf_109_i_clk),
    .D(net3930),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21731_ (.CLK(clknet_leaf_108_i_clk),
    .D(net4005),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21732_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3568),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21733_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4805),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21734_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4736),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21735_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4504),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21736_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3664),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21737_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3512),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21738_ (.CLK(clknet_leaf_98_i_clk),
    .D(net4701),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21739_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3497),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21740_ (.CLK(clknet_leaf_99_i_clk),
    .D(net4557),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21741_ (.CLK(clknet_leaf_100_i_clk),
    .D(net4606),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21742_ (.CLK(clknet_leaf_100_i_clk),
    .D(net5478),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21743_ (.CLK(clknet_leaf_99_i_clk),
    .D(net4593),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21744_ (.CLK(clknet_leaf_98_i_clk),
    .D(net4827),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21745_ (.CLK(clknet_leaf_131_i_clk),
    .D(net4638),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21746_ (.CLK(clknet_leaf_134_i_clk),
    .D(net3541),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21747_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3622),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21748_ (.CLK(clknet_leaf_132_i_clk),
    .D(net3578),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21749_ (.CLK(clknet_leaf_131_i_clk),
    .D(net4689),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21750_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3681),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21751_ (.CLK(clknet_leaf_132_i_clk),
    .D(net4563),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21752_ (.CLK(clknet_leaf_99_i_clk),
    .D(net4712),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21753_ (.CLK(clknet_leaf_101_i_clk),
    .D(net5047),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21754_ (.CLK(clknet_leaf_124_i_clk),
    .D(net3953),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21755_ (.CLK(clknet_leaf_83_i_clk),
    .D(net5986),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _21756_ (.CLK(clknet_leaf_29_i_clk),
    .D(net5210),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_1 _21757_ (.CLK(clknet_leaf_84_i_clk),
    .D(net4104),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21758_ (.CLK(clknet_leaf_111_i_clk),
    .D(net4026),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21759_ (.CLK(clknet_leaf_111_i_clk),
    .D(net4114),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(clknet_leaf_111_i_clk),
    .D(net7683),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(clknet_leaf_111_i_clk),
    .D(net4130),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21762_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01249_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21763_ (.CLK(clknet_leaf_83_i_clk),
    .D(net4072),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21764_ (.CLK(clknet_leaf_83_i_clk),
    .D(net4093),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21765_ (.CLK(clknet_leaf_83_i_clk),
    .D(net4100),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21766_ (.CLK(clknet_leaf_83_i_clk),
    .D(net3997),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21767_ (.CLK(clknet_leaf_15_i_clk),
    .D(net1342),
    .Q(\rbzero.spi_registers.new_texadd[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21768_ (.CLK(clknet_leaf_10_i_clk),
    .D(net1557),
    .Q(\rbzero.spi_registers.new_texadd[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21769_ (.CLK(clknet_leaf_11_i_clk),
    .D(net1370),
    .Q(\rbzero.spi_registers.new_texadd[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21770_ (.CLK(clknet_leaf_11_i_clk),
    .D(net1306),
    .Q(\rbzero.spi_registers.new_texadd[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21771_ (.CLK(clknet_leaf_45_i_clk),
    .D(net1461),
    .Q(\rbzero.spi_registers.new_texadd[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21772_ (.CLK(clknet_leaf_45_i_clk),
    .D(net1467),
    .Q(\rbzero.spi_registers.new_texadd[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21773_ (.CLK(clknet_leaf_48_i_clk),
    .D(net1265),
    .Q(\rbzero.spi_registers.new_texadd[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(clknet_leaf_48_i_clk),
    .D(net1443),
    .Q(\rbzero.spi_registers.new_texadd[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21775_ (.CLK(clknet_leaf_46_i_clk),
    .D(net1216),
    .Q(\rbzero.spi_registers.new_texadd[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21776_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1324),
    .Q(\rbzero.spi_registers.new_texadd[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21777_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1476),
    .Q(\rbzero.spi_registers.new_texadd[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21778_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1787),
    .Q(\rbzero.spi_registers.new_texadd[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21779_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1202),
    .Q(\rbzero.spi_registers.new_texadd[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(clknet_leaf_3_i_clk),
    .D(net1504),
    .Q(\rbzero.spi_registers.new_texadd[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21781_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1357),
    .Q(\rbzero.spi_registers.new_texadd[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21782_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1687),
    .Q(\rbzero.spi_registers.new_texadd[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21783_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1578),
    .Q(\rbzero.spi_registers.new_texadd[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21784_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1769),
    .Q(\rbzero.spi_registers.new_texadd[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(clknet_leaf_1_i_clk),
    .D(net1364),
    .Q(\rbzero.spi_registers.new_texadd[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21786_ (.CLK(clknet_leaf_1_i_clk),
    .D(net2222),
    .Q(\rbzero.spi_registers.new_texadd[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21787_ (.CLK(clknet_leaf_4_i_clk),
    .D(net1401),
    .Q(\rbzero.spi_registers.new_texadd[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21788_ (.CLK(clknet_leaf_20_i_clk),
    .D(net1592),
    .Q(\rbzero.spi_registers.new_texadd[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21789_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1221),
    .Q(\rbzero.spi_registers.new_texadd[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21790_ (.CLK(clknet_leaf_19_i_clk),
    .D(net1388),
    .Q(\rbzero.spi_registers.new_texadd[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21791_ (.CLK(net233),
    .D(net1413),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21792_ (.CLK(net234),
    .D(net2353),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21793_ (.CLK(net235),
    .D(net2705),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21794_ (.CLK(net236),
    .D(net2932),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21795_ (.CLK(net237),
    .D(net2151),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21796_ (.CLK(net238),
    .D(net662),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(net239),
    .D(net2538),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21798_ (.CLK(net240),
    .D(net2580),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21799_ (.CLK(net241),
    .D(net1829),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21800_ (.CLK(net242),
    .D(net2603),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(net243),
    .D(net2666),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21802_ (.CLK(net244),
    .D(net1227),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21803_ (.CLK(net245),
    .D(net2980),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21804_ (.CLK(net246),
    .D(net2885),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(net247),
    .D(net2308),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(net248),
    .D(net1071),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21807_ (.CLK(net249),
    .D(net2369),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(net250),
    .D(net2559),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(net251),
    .D(net2696),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(net252),
    .D(net3245),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(net253),
    .D(net2109),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(net254),
    .D(net3094),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(net255),
    .D(net2276),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(net256),
    .D(net1662),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21815_ (.CLK(net257),
    .D(net1799),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21816_ (.CLK(net258),
    .D(net1019),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21817_ (.CLK(net259),
    .D(net2241),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(net260),
    .D(net1990),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21819_ (.CLK(net261),
    .D(net2825),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21820_ (.CLK(net262),
    .D(net1890),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(net263),
    .D(net2634),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21822_ (.CLK(net264),
    .D(net2216),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21823_ (.CLK(net265),
    .D(net1951),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21824_ (.CLK(net266),
    .D(net1957),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21825_ (.CLK(net267),
    .D(net1410),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21826_ (.CLK(net268),
    .D(net1187),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21827_ (.CLK(net269),
    .D(net2359),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21828_ (.CLK(net270),
    .D(net2708),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21829_ (.CLK(net271),
    .D(net2335),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21830_ (.CLK(net272),
    .D(net2511),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21831_ (.CLK(net273),
    .D(net2779),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21832_ (.CLK(net274),
    .D(net2556),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21833_ (.CLK(net275),
    .D(net2939),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(net276),
    .D(net1354),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(net277),
    .D(net2002),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(net278),
    .D(net999),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(net279),
    .D(net2737),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(net280),
    .D(net2624),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21839_ (.CLK(net281),
    .D(net2992),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(net282),
    .D(net2669),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21841_ (.CLK(net283),
    .D(net2065),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21842_ (.CLK(net284),
    .D(net1160),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21843_ (.CLK(net285),
    .D(net2547),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21844_ (.CLK(net286),
    .D(net2210),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(net287),
    .D(net2255),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21846_ (.CLK(net288),
    .D(net1528),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21847_ (.CLK(net289),
    .D(net2115),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21848_ (.CLK(net290),
    .D(net3165),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(net291),
    .D(net2868),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(net292),
    .D(net2287),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(net293),
    .D(net2136),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(net294),
    .D(net1300),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21853_ (.CLK(net295),
    .D(net2684),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(net296),
    .D(net2847),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(net297),
    .D(net2699),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(net298),
    .D(net657),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(net299),
    .D(net2859),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(net300),
    .D(net2118),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(net301),
    .D(net1893),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(net302),
    .D(net1975),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(net303),
    .D(net2356),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(net304),
    .D(net2717),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21863_ (.CLK(net305),
    .D(net2672),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(net306),
    .D(net1274),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(net307),
    .D(net1717),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(net308),
    .D(net1132),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(net309),
    .D(net1874),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(net310),
    .D(net2493),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(net311),
    .D(net3031),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(net312),
    .D(net2019),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(net313),
    .D(net1922),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(net314),
    .D(net1271),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21873_ (.CLK(net315),
    .D(net1741),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21874_ (.CLK(net316),
    .D(net2267),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(net317),
    .D(net2112),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(net318),
    .D(net926),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(net319),
    .D(net2484),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21878_ (.CLK(net320),
    .D(net2302),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21879_ (.CLK(net321),
    .D(net2219),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21880_ (.CLK(net322),
    .D(net1784),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(net323),
    .D(net2724),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21882_ (.CLK(net324),
    .D(net3265),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(net325),
    .D(net3091),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(net326),
    .D(net3248),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(net327),
    .D(net3109),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(net328),
    .D(net644),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(net329),
    .D(net2618),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(net330),
    .D(net2733),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(net331),
    .D(net3178),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(net332),
    .D(net2565),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(net333),
    .D(net2606),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(net334),
    .D(net1141),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(net335),
    .D(net1902),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(net336),
    .D(net3072),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21895_ (.CLK(net337),
    .D(net2284),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(net338),
    .D(net1082),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(net339),
    .D(net2455),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21898_ (.CLK(net340),
    .D(net2237),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(net341),
    .D(net2591),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(net342),
    .D(net2037),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(net343),
    .D(net3204),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(net344),
    .D(net2902),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(net345),
    .D(net1966),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(net346),
    .D(net2016),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(net347),
    .D(net2577),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(net348),
    .D(net805),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(net349),
    .D(net2054),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(net350),
    .D(net2693),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21909_ (.CLK(net351),
    .D(net2925),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(net352),
    .D(net2888),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21911_ (.CLK(net353),
    .D(net1807),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(net354),
    .D(net2687),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(net355),
    .D(net2422),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(net356),
    .D(net2293),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21915_ (.CLK(net357),
    .D(net2828),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(net358),
    .D(net1589),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(net359),
    .D(net2478),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(net360),
    .D(net2505),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(net361),
    .D(net1598),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(net362),
    .D(net3106),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(net363),
    .D(net2464),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(net364),
    .D(net2597),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(net365),
    .D(net1181),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(net366),
    .D(net2401),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(net367),
    .D(net2025),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21926_ (.CLK(net368),
    .D(net632),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(net369),
    .D(net2967),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(net370),
    .D(net2740),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(net371),
    .D(net2850),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21930_ (.CLK(net372),
    .D(net3154),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21931_ (.CLK(net373),
    .D(net3251),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(net374),
    .D(net1175),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(net375),
    .D(net2031),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(net376),
    .D(net2087),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(net377),
    .D(net2785),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(net378),
    .D(net1259),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(net379),
    .D(net2640),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(net380),
    .D(net1963),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(net381),
    .D(net2523),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(net382),
    .D(net2404),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(net383),
    .D(net2653),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(net384),
    .D(net2998),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(net385),
    .D(net1654),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21944_ (.CLK(net386),
    .D(net2517),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(net387),
    .D(net1987),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21946_ (.CLK(net388),
    .D(net1085),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21947_ (.CLK(net389),
    .D(net3171),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21948_ (.CLK(net390),
    .D(net2972),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21949_ (.CLK(net391),
    .D(net2568),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21950_ (.CLK(net392),
    .D(net2410),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(net393),
    .D(net1315),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(net394),
    .D(net2461),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(net395),
    .D(net2473),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(net396),
    .D(net2571),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(net397),
    .D(net2431),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(net398),
    .D(net966),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(net399),
    .D(net2178),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21958_ (.CLK(net400),
    .D(net2535),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(net401),
    .D(net1937),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21960_ (.CLK(net402),
    .D(net2434),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(net403),
    .D(net2553),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(net404),
    .D(net2378),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21963_ (.CLK(net405),
    .D(net2752),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(net406),
    .D(net1193),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(net407),
    .D(net2290),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(net408),
    .D(net1129),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21967_ (.CLK(net409),
    .D(net2010),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(net410),
    .D(net1452),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(net411),
    .D(net2520),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(net412),
    .D(net2822),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21971_ (.CLK(net413),
    .D(net3001),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(net414),
    .D(net2419),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(net415),
    .D(net1488),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(net416),
    .D(net2702),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(net417),
    .D(net2246),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(net418),
    .D(net1190),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(net419),
    .D(net1996),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(net420),
    .D(net2051),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(net421),
    .D(net2228),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(net422),
    .D(net2749),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(net423),
    .D(net2812),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(net424),
    .D(net2909),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(net425),
    .D(net1796),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(net426),
    .D(net2795),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(net427),
    .D(net1750),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(net428),
    .D(net592),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(net429),
    .D(net2594),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(net430),
    .D(net2763),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(net431),
    .D(net2320),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(net432),
    .D(net2663),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21991_ (.CLK(net433),
    .D(net2145),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21992_ (.CLK(net434),
    .D(net2124),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(net435),
    .D(net1126),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(net436),
    .D(net1928),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(net437),
    .D(net3358),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(net438),
    .D(net1091),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(net439),
    .D(net2189),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21998_ (.CLK(net440),
    .D(net2730),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(net441),
    .D(net2341),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(net442),
    .D(net2452),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(net443),
    .D(net1522),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(net444),
    .D(net2621),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(net445),
    .D(net2034),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(net446),
    .D(net2637),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(net447),
    .D(net2296),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(net448),
    .D(net768),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(net449),
    .D(net2093),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(net450),
    .D(net2627),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(net451),
    .D(net1847),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(net452),
    .D(net2142),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(net453),
    .D(net1208),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22012_ (.CLK(net454),
    .D(net2392),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22013_ (.CLK(net455),
    .D(net2157),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(net456),
    .D(net2407),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(net457),
    .D(net1835),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(net458),
    .D(net2096),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(net459),
    .D(net1855),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(net460),
    .D(net2757),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(net461),
    .D(net2952),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(net462),
    .D(net1519),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(net463),
    .D(net2103),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22022_ (.CLK(net464),
    .D(net2045),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(net465),
    .D(net2425),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(net466),
    .D(net1850),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(net467),
    .D(net2995),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(net468),
    .D(net1074),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(net469),
    .D(net1896),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(net470),
    .D(net2819),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(net471),
    .D(net2612),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(net472),
    .D(net2583),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(net473),
    .D(net1440),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(net474),
    .D(net2678),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22033_ (.CLK(net475),
    .D(net2446),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(net476),
    .D(net2961),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(net477),
    .D(net2249),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22036_ (.CLK(net478),
    .D(net1144),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(net479),
    .D(net2386),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(net480),
    .D(net2329),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(net481),
    .D(net2203),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(net482),
    .D(net2160),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(net483),
    .D(net2532),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(net484),
    .D(net1844),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(net485),
    .D(net2916),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(net486),
    .D(net2788),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(net487),
    .D(net2305),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22046_ (.CLK(net488),
    .D(net2949),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22047_ (.CLK(net489),
    .D(net1277),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22048_ (.CLK(net490),
    .D(net1531),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22049_ (.CLK(net491),
    .D(net1960),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22050_ (.CLK(net492),
    .D(net1385),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22051_ (.CLK(net493),
    .D(net2326),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22052_ (.CLK(net494),
    .D(net2338),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22053_ (.CLK(net495),
    .D(net1757),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22054_ (.CLK(net496),
    .D(net2526),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22055_ (.CLK(net497),
    .D(net2372),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22056_ (.CLK(net498),
    .D(net1066),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22057_ (.CLK(net499),
    .D(net1117),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22058_ (.CLK(net500),
    .D(net2273),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22059_ (.CLK(net501),
    .D(net2882),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22060_ (.CLK(net502),
    .D(net2769),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22061_ (.CLK(net503),
    .D(net2344),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22062_ (.CLK(net504),
    .D(net2743),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22063_ (.CLK(net505),
    .D(net2022),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22064_ (.CLK(net506),
    .D(net2643),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22065_ (.CLK(net507),
    .D(net1841),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22066_ (.CLK(net508),
    .D(net935),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22067_ (.CLK(net509),
    .D(net1914),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22068_ (.CLK(net510),
    .D(net1993),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22069_ (.CLK(net511),
    .D(net2175),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22070_ (.CLK(net512),
    .D(net2467),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22071_ (.CLK(net513),
    .D(net2721),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22072_ (.CLK(net514),
    .D(net1940),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22073_ (.CLK(net515),
    .D(net2983),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22074_ (.CLK(net516),
    .D(net2154),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22075_ (.CLK(net517),
    .D(net3116),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22076_ (.CLK(net518),
    .D(net977),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22077_ (.CLK(net519),
    .D(net2799),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22078_ (.CLK(net520),
    .D(net2375),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22079_ (.CLK(net521),
    .D(net2252),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22080_ (.CLK(net522),
    .D(net2776),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22081_ (.CLK(net523),
    .D(net1237),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22082_ (.CLK(net524),
    .D(net2562),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22083_ (.CLK(net525),
    .D(net2792),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22084_ (.CLK(net526),
    .D(net2042),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22085_ (.CLK(net527),
    .D(net3242),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22086_ (.CLK(net528),
    .D(net586),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22087_ (.CLK(net149),
    .D(net2261),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22088_ (.CLK(net150),
    .D(net2659),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22089_ (.CLK(net151),
    .D(net2013),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22090_ (.CLK(net152),
    .D(net2501),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22091_ (.CLK(net153),
    .D(net2231),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22092_ (.CLK(net154),
    .D(net2130),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22093_ (.CLK(net155),
    .D(net2986),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22094_ (.CLK(net156),
    .D(net3130),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22095_ (.CLK(net157),
    .D(net2440),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22096_ (.CLK(net158),
    .D(net1042),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22097_ (.CLK(net159),
    .D(net2498),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22098_ (.CLK(net160),
    .D(net2690),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22099_ (.CLK(net161),
    .D(net2782),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22100_ (.CLK(net162),
    .D(net2133),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22101_ (.CLK(net163),
    .D(net2121),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22102_ (.CLK(net164),
    .D(net2853),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22103_ (.CLK(net165),
    .D(net1978),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22104_ (.CLK(net166),
    .D(net2299),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22105_ (.CLK(net167),
    .D(net2350),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22106_ (.CLK(net168),
    .D(net1607),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22107_ (.CLK(net145),
    .D(net2028),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22108_ (.CLK(net146),
    .D(net2550),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22109_ (.CLK(net147),
    .D(net3069),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22110_ (.CLK(net148),
    .D(net2395),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22111_ (.CLK(clknet_leaf_89_i_clk),
    .D(net4924),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22112_ (.CLK(clknet_leaf_87_i_clk),
    .D(net921),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22113_ (.CLK(clknet_leaf_62_i_clk),
    .D(net4970),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _22114_ (.CLK(clknet_leaf_54_i_clk),
    .D(net4986),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _22115_ (.CLK(clknet_leaf_62_i_clk),
    .D(net5386),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22116_ (.CLK(clknet_leaf_55_i_clk),
    .D(net5402),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22117_ (.CLK(clknet_leaf_57_i_clk),
    .D(net5382),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22118_ (.CLK(clknet_leaf_57_i_clk),
    .D(net5406),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22119_ (.CLK(clknet_leaf_57_i_clk),
    .D(net5254),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _22120_ (.CLK(clknet_leaf_55_i_clk),
    .D(net5342),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _22121_ (.CLK(clknet_leaf_54_i_clk),
    .D(net5378),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _22122_ (.CLK(clknet_leaf_54_i_clk),
    .D(net4974),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _22123_ (.CLK(clknet_leaf_54_i_clk),
    .D(net4982),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _22124_ (.CLK(clknet_leaf_54_i_clk),
    .D(net5450),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22125_ (.CLK(clknet_leaf_54_i_clk),
    .D(net5494),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22126_ (.CLK(clknet_leaf_53_i_clk),
    .D(net5490),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22127_ (.CLK(clknet_leaf_53_i_clk),
    .D(net5624),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22128_ (.CLK(clknet_leaf_53_i_clk),
    .D(net5583),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22129_ (.CLK(clknet_leaf_53_i_clk),
    .D(net5694),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22130_ (.CLK(clknet_leaf_53_i_clk),
    .D(net5524),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22131_ (.CLK(clknet_leaf_52_i_clk),
    .D(net5728),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22132_ (.CLK(clknet_leaf_52_i_clk),
    .D(net5741),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22133_ (.CLK(clknet_leaf_56_i_clk),
    .D(net5482),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22134_ (.CLK(clknet_leaf_56_i_clk),
    .D(net5611),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22135_ (.CLK(clknet_leaf_85_i_clk),
    .D(net4087),
    .Q(\rbzero.trace_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22136_ (.CLK(clknet_leaf_85_i_clk),
    .D(net3629),
    .Q(\rbzero.trace_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22137_ (.CLK(clknet_leaf_85_i_clk),
    .D(net3977),
    .Q(\rbzero.trace_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22138_ (.CLK(clknet_leaf_85_i_clk),
    .D(net3873),
    .Q(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22139_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01626_),
    .Q(\reg_gpout[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22140_ (.CLK(clknet_leaf_24_i_clk),
    .D(_01627_),
    .Q(\reg_gpout[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22141_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01628_),
    .Q(\reg_gpout[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22142_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01629_),
    .Q(\reg_gpout[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22143_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01630_),
    .Q(\reg_gpout[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22144_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01631_),
    .Q(\reg_gpout[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22145_ (.CLK(clknet_leaf_56_i_clk),
    .D(net901),
    .Q(reg_hsync));
 sky130_fd_sc_hd__dfxtp_1 _22146_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01633_),
    .Q(reg_vsync));
 sky130_fd_sc_hd__dfxtp_1 _22147_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01634_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22148_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01635_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22149_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01636_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22150_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01637_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22151_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01638_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22152_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01639_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22153_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01640_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22154_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01641_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22155_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01642_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22156_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01643_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22157_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01644_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22158_ (.CLK(clknet_leaf_88_i_clk),
    .D(net4934),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22159_ (.CLK(clknet_leaf_88_i_clk),
    .D(net1094),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22160_ (.CLK(clknet_leaf_96_i_clk),
    .D(net5035),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22161_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4717),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22162_ (.CLK(clknet_leaf_94_i_clk),
    .D(net4889),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22163_ (.CLK(clknet_leaf_94_i_clk),
    .D(net4854),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22164_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4426),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22165_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4602),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22166_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4881),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22167_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4850),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22168_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4942),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22169_ (.CLK(clknet_leaf_91_i_clk),
    .D(net1097),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22170_ (.CLK(clknet_leaf_87_i_clk),
    .D(net4950),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22171_ (.CLK(clknet_leaf_89_i_clk),
    .D(net680),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22172_ (.CLK(clknet_leaf_67_i_clk),
    .D(net4930),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22173_ (.CLK(clknet_4_7__leaf_i_clk),
    .D(net2615),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22174_ (.CLK(clknet_leaf_68_i_clk),
    .D(net4938),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22175_ (.CLK(clknet_leaf_68_i_clk),
    .D(net1100),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03506_ (.A(_03506_),
    .X(clknet_0__03506_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03507_ (.A(_03507_),
    .X(clknet_0__03507_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03508_ (.A(_03508_),
    .X(clknet_0__03508_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03509_ (.A(_03509_),
    .X(clknet_0__03509_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03510_ (.A(_03510_),
    .X(clknet_0__03510_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03511_ (.A(_03511_),
    .X(clknet_0__03511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03512_ (.A(_03512_),
    .X(clknet_0__03512_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03513_ (.A(_03513_),
    .X(clknet_0__03513_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03514_ (.A(_03514_),
    .X(clknet_0__03514_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03840_ (.A(_03840_),
    .X(clknet_0__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03841_ (.A(_03841_),
    .X(clknet_0__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03842_ (.A(_03842_),
    .X(clknet_0__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03843_ (.A(_03843_),
    .X(clknet_0__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03844_ (.A(_03844_),
    .X(clknet_0__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03845_ (.A(_03845_),
    .X(clknet_0__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03846_ (.A(_03846_),
    .X(clknet_0__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03847_ (.A(_03847_),
    .X(clknet_0__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03848_ (.A(_03848_),
    .X(clknet_0__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03849_ (.A(_03849_),
    .X(clknet_0__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03850_ (.A(_03850_),
    .X(clknet_0__03850_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03851_ (.A(_03851_),
    .X(clknet_0__03851_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03852_ (.A(_03852_),
    .X(clknet_0__03852_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03853_ (.A(_03853_),
    .X(clknet_0__03853_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03854_ (.A(_03854_),
    .X(clknet_0__03854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03855_ (.A(_03855_),
    .X(clknet_0__03855_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03856_ (.A(_03856_),
    .X(clknet_0__03856_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03857_ (.A(_03857_),
    .X(clknet_0__03857_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03858_ (.A(_03858_),
    .X(clknet_0__03858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03859_ (.A(_03859_),
    .X(clknet_0__03859_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03860_ (.A(_03860_),
    .X(clknet_0__03860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03861_ (.A(_03861_),
    .X(clknet_0__03861_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03862_ (.A(_03862_),
    .X(clknet_0__03862_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03863_ (.A(_03863_),
    .X(clknet_0__03863_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03864_ (.A(_03864_),
    .X(clknet_0__03864_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03865_ (.A(_03865_),
    .X(clknet_0__03865_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03866_ (.A(_03866_),
    .X(clknet_0__03866_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03867_ (.A(_03867_),
    .X(clknet_0__03867_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03868_ (.A(_03868_),
    .X(clknet_0__03868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03869_ (.A(_03869_),
    .X(clknet_0__03869_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03870_ (.A(_03870_),
    .X(clknet_0__03870_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03871_ (.A(_03871_),
    .X(clknet_0__03871_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03872_ (.A(_03872_),
    .X(clknet_0__03872_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05645_ (.A(_05645_),
    .X(clknet_0__05645_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05688_ (.A(_05688_),
    .X(clknet_0__05688_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05742_ (.A(_05742_),
    .X(clknet_0__05742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05794_ (.A(_05794_),
    .X(clknet_0__05794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05847_ (.A(_05847_),
    .X(clknet_0__05847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05898_ (.A(_05898_),
    .X(clknet_0__05898_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05946_ (.A(_05946_),
    .X(clknet_0__05946_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03506_ (.A(clknet_0__03506_),
    .X(clknet_1_0__leaf__03506_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03507_ (.A(clknet_0__03507_),
    .X(clknet_1_0__leaf__03507_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03508_ (.A(clknet_0__03508_),
    .X(clknet_1_0__leaf__03508_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03509_ (.A(clknet_0__03509_),
    .X(clknet_1_0__leaf__03509_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03510_ (.A(clknet_0__03510_),
    .X(clknet_1_0__leaf__03510_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03511_ (.A(clknet_0__03511_),
    .X(clknet_1_0__leaf__03511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03512_ (.A(clknet_0__03512_),
    .X(clknet_1_0__leaf__03512_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03513_ (.A(clknet_0__03513_),
    .X(clknet_1_0__leaf__03513_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03514_ (.A(clknet_0__03514_),
    .X(clknet_1_0__leaf__03514_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03840_ (.A(clknet_0__03840_),
    .X(clknet_1_0__leaf__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03841_ (.A(clknet_0__03841_),
    .X(clknet_1_0__leaf__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03842_ (.A(clknet_0__03842_),
    .X(clknet_1_0__leaf__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03843_ (.A(clknet_0__03843_),
    .X(clknet_1_0__leaf__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03844_ (.A(clknet_0__03844_),
    .X(clknet_1_0__leaf__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03845_ (.A(clknet_0__03845_),
    .X(clknet_1_0__leaf__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03846_ (.A(clknet_0__03846_),
    .X(clknet_1_0__leaf__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03847_ (.A(clknet_0__03847_),
    .X(clknet_1_0__leaf__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03848_ (.A(clknet_0__03848_),
    .X(clknet_1_0__leaf__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03849_ (.A(clknet_0__03849_),
    .X(clknet_1_0__leaf__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03850_ (.A(clknet_0__03850_),
    .X(clknet_1_0__leaf__03850_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03851_ (.A(clknet_0__03851_),
    .X(clknet_1_0__leaf__03851_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03852_ (.A(clknet_0__03852_),
    .X(clknet_1_0__leaf__03852_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03853_ (.A(clknet_0__03853_),
    .X(clknet_1_0__leaf__03853_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03854_ (.A(clknet_0__03854_),
    .X(clknet_1_0__leaf__03854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03855_ (.A(clknet_0__03855_),
    .X(clknet_1_0__leaf__03855_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03856_ (.A(clknet_0__03856_),
    .X(clknet_1_0__leaf__03856_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03857_ (.A(clknet_0__03857_),
    .X(clknet_1_0__leaf__03857_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03858_ (.A(clknet_0__03858_),
    .X(clknet_1_0__leaf__03858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03859_ (.A(clknet_0__03859_),
    .X(clknet_1_0__leaf__03859_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03860_ (.A(clknet_0__03860_),
    .X(clknet_1_0__leaf__03860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03861_ (.A(clknet_0__03861_),
    .X(clknet_1_0__leaf__03861_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03862_ (.A(clknet_0__03862_),
    .X(clknet_1_0__leaf__03862_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03863_ (.A(clknet_0__03863_),
    .X(clknet_1_0__leaf__03863_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03864_ (.A(clknet_0__03864_),
    .X(clknet_1_0__leaf__03864_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03865_ (.A(clknet_0__03865_),
    .X(clknet_1_0__leaf__03865_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03866_ (.A(clknet_0__03866_),
    .X(clknet_1_0__leaf__03866_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03867_ (.A(clknet_0__03867_),
    .X(clknet_1_0__leaf__03867_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03868_ (.A(clknet_0__03868_),
    .X(clknet_1_0__leaf__03868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03869_ (.A(clknet_0__03869_),
    .X(clknet_1_0__leaf__03869_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03870_ (.A(clknet_0__03870_),
    .X(clknet_1_0__leaf__03870_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03871_ (.A(clknet_0__03871_),
    .X(clknet_1_0__leaf__03871_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03872_ (.A(clknet_0__03872_),
    .X(clknet_1_0__leaf__03872_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05645_ (.A(clknet_0__05645_),
    .X(clknet_1_0__leaf__05645_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05688_ (.A(clknet_0__05688_),
    .X(clknet_1_0__leaf__05688_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05742_ (.A(clknet_0__05742_),
    .X(clknet_1_0__leaf__05742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05794_ (.A(clknet_0__05794_),
    .X(clknet_1_0__leaf__05794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05847_ (.A(clknet_0__05847_),
    .X(clknet_1_0__leaf__05847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05898_ (.A(clknet_0__05898_),
    .X(clknet_1_0__leaf__05898_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05946_ (.A(clknet_0__05946_),
    .X(clknet_1_0__leaf__05946_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03506_ (.A(clknet_0__03506_),
    .X(clknet_1_1__leaf__03506_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03507_ (.A(clknet_0__03507_),
    .X(clknet_1_1__leaf__03507_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03508_ (.A(clknet_0__03508_),
    .X(clknet_1_1__leaf__03508_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03509_ (.A(clknet_0__03509_),
    .X(clknet_1_1__leaf__03509_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03510_ (.A(clknet_0__03510_),
    .X(clknet_1_1__leaf__03510_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03511_ (.A(clknet_0__03511_),
    .X(clknet_1_1__leaf__03511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03512_ (.A(clknet_0__03512_),
    .X(clknet_1_1__leaf__03512_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03513_ (.A(clknet_0__03513_),
    .X(clknet_1_1__leaf__03513_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03514_ (.A(clknet_0__03514_),
    .X(clknet_1_1__leaf__03514_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03840_ (.A(clknet_0__03840_),
    .X(clknet_1_1__leaf__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03841_ (.A(clknet_0__03841_),
    .X(clknet_1_1__leaf__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03842_ (.A(clknet_0__03842_),
    .X(clknet_1_1__leaf__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03843_ (.A(clknet_0__03843_),
    .X(clknet_1_1__leaf__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03844_ (.A(clknet_0__03844_),
    .X(clknet_1_1__leaf__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03845_ (.A(clknet_0__03845_),
    .X(clknet_1_1__leaf__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03846_ (.A(clknet_0__03846_),
    .X(clknet_1_1__leaf__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03847_ (.A(clknet_0__03847_),
    .X(clknet_1_1__leaf__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03848_ (.A(clknet_0__03848_),
    .X(clknet_1_1__leaf__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03849_ (.A(clknet_0__03849_),
    .X(clknet_1_1__leaf__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03850_ (.A(clknet_0__03850_),
    .X(clknet_1_1__leaf__03850_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03851_ (.A(clknet_0__03851_),
    .X(clknet_1_1__leaf__03851_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03852_ (.A(clknet_0__03852_),
    .X(clknet_1_1__leaf__03852_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03853_ (.A(clknet_0__03853_),
    .X(clknet_1_1__leaf__03853_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03854_ (.A(clknet_0__03854_),
    .X(clknet_1_1__leaf__03854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03855_ (.A(clknet_0__03855_),
    .X(clknet_1_1__leaf__03855_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03856_ (.A(clknet_0__03856_),
    .X(clknet_1_1__leaf__03856_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03857_ (.A(clknet_0__03857_),
    .X(clknet_1_1__leaf__03857_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03858_ (.A(clknet_0__03858_),
    .X(clknet_1_1__leaf__03858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03859_ (.A(clknet_0__03859_),
    .X(clknet_1_1__leaf__03859_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03860_ (.A(clknet_0__03860_),
    .X(clknet_1_1__leaf__03860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03861_ (.A(clknet_0__03861_),
    .X(clknet_1_1__leaf__03861_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03862_ (.A(clknet_0__03862_),
    .X(clknet_1_1__leaf__03862_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03863_ (.A(clknet_0__03863_),
    .X(clknet_1_1__leaf__03863_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03864_ (.A(clknet_0__03864_),
    .X(clknet_1_1__leaf__03864_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03865_ (.A(clknet_0__03865_),
    .X(clknet_1_1__leaf__03865_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03866_ (.A(clknet_0__03866_),
    .X(clknet_1_1__leaf__03866_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03867_ (.A(clknet_0__03867_),
    .X(clknet_1_1__leaf__03867_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03868_ (.A(clknet_0__03868_),
    .X(clknet_1_1__leaf__03868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03869_ (.A(clknet_0__03869_),
    .X(clknet_1_1__leaf__03869_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03870_ (.A(clknet_0__03870_),
    .X(clknet_1_1__leaf__03870_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03871_ (.A(clknet_0__03871_),
    .X(clknet_1_1__leaf__03871_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03872_ (.A(clknet_0__03872_),
    .X(clknet_1_1__leaf__03872_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05645_ (.A(clknet_0__05645_),
    .X(clknet_1_1__leaf__05645_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05688_ (.A(clknet_0__05688_),
    .X(clknet_1_1__leaf__05688_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05742_ (.A(clknet_0__05742_),
    .X(clknet_1_1__leaf__05742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05794_ (.A(clknet_0__05794_),
    .X(clknet_1_1__leaf__05794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05847_ (.A(clknet_0__05847_),
    .X(clknet_1_1__leaf__05847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05898_ (.A(clknet_0__05898_),
    .X(clknet_1_1__leaf__05898_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05946_ (.A(clknet_0__05946_),
    .X(clknet_1_1__leaf__05946_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_4_0__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_4_10__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_4_11__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_4_12__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_4_13__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_4_14__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_4_15__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_4_1__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_4_2__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_4_3__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_4_4__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_4_5__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_4_6__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_4_7__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_4_8__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_4_9__leaf_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_100_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_101_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_102_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_103_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_104_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_105_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_106_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_107_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_108_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_109_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_110_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_111_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_112_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_113_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_114_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_115_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_116_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_117_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_118_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_119_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_120_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_121_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_122_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_123_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_124_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_125_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_126_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_127_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_128_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_129_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_130_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_131_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_132_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_133_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_134_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_i_clk (.A(clknet_4_4__leaf_i_clk),
    .X(clknet_leaf_135_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_4_3__leaf_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_4_11__leaf_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_4_1__leaf_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_4_11__leaf_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_4_10__leaf_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_4_10__leaf_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_4_10__leaf_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_4_10__leaf_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_4_10__leaf_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_4_10__leaf_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_4_10__leaf_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_4_9__leaf_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_4_9__leaf_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_4_9__leaf_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_4_9__leaf_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_4_8__leaf_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_4_9__leaf_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_4_8__leaf_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_4_8__leaf_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_4_8__leaf_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_4_8__leaf_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_4_14__leaf_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_4_11__leaf_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_4_11__leaf_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_4_14__leaf_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_4_14__leaf_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_4_11__leaf_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_4_14__leaf_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_4_14__leaf_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_4_14__leaf_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_4_12__leaf_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_4_12__leaf_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_4_13__leaf_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_4_13__leaf_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_4_13__leaf_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_4_13__leaf_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_4_13__leaf_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_4_12__leaf_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_4_12__leaf_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_4_12__leaf_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_4_12__leaf_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_4_13__leaf_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_4_12__leaf_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_4_15__leaf_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_4_6__leaf_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_4_0__leaf_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_4_7__leaf_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_4_5__leaf_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_4_2__leaf_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net4720),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(net6549),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(_01333_),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\rbzero.tex_r1[2] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(net5551),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_01535_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(net6013),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_03347_),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(_00905_),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(net5815),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(_03060_),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net2078),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_00707_),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(net6491),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_02489_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(_00578_),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(net3595),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(_03416_),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_00957_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(net6447),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_03435_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(_00970_),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net4503),
    .X(net629));
 sky130_fd_sc_hd__buf_2 hold1020 (.A(net7696),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(_02977_),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(net5880),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(net5517),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(net5519),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(net6398),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_03466_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(_00998_),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(net6551),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(_03816_),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net6033),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_01255_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(net3120),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_03053_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(_00701_),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(net6020),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(net6022),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_00916_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(net6009),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(net6011),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(_00913_),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net6035),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(net3008),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(_03592_),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_01154_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(net6515),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(net6517),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(_00985_),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(net6559),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(_02998_),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_00651_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(net6495),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_01413_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(net6497),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(_01270_),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(net6660),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(net6662),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_01092_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(net5512),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_03390_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(_00937_),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(net8359),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(net4272),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net6029),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(net6586),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(net6588),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_01403_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(net6079),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(net6081),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(_01275_),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(net6049),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(_03356_),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_00912_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(net6292),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net6031),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(net6294),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(_01406_),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(net6159),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(net6161),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_00594_),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(net6527),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(net6529),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(_00590_),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(net6580),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(net6582),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_01041_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_01593_),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(_06503_),
    .X(net3638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(net8108),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(net4794),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(net5530),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(net5532),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(net6664),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(net5785),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_00720_),
    .X(net1615));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1089 (.A(net5580),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net6815),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(net5582),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(net6730),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(net6732),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(_00684_),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(net3896),
    .X(net1621));
 sky130_fd_sc_hd__buf_4 hold1095 (.A(net3898),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_03389_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(_00936_),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(net6055),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(_03358_),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net4452),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_00914_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(net6565),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(net6567),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(_00975_),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(net6453),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(_02490_),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_00579_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(net5499),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_03369_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(_00921_),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net8102),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(net6573),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(net6575),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_00960_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(net5525),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_03375_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(_00925_),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(net6545),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(_03367_),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_00919_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(net3297),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net4735),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_03032_),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(_00682_),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(net6618),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(net6620),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_00987_),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(net6642),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(net6644),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(_01430_),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(net3561),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(_03417_),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net4967),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_00958_),
    .X(net1657));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1131 (.A(net8155),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(net5515),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(net6698),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(net6700),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(_01301_),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(net7954),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(net4586),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(net6561),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(net6563),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net4969),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_01009_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(net6541),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_03438_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(_00973_),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(net6577),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(_03370_),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_00922_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\rbzero.row_render.size[8] ),
    .X(net3686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(net8112),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(net4800),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net6071),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(net6584),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(_02497_),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_00585_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(net4897),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(net4759),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(net7309),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(net6694),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(_00653_),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(net6569),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(net6571),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net6073),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_01269_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(net6648),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_03546_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(_01112_),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(net6598),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(_03464_),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_00996_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(net6503),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_03461_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(_00993_),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_01373_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(net6622),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(net6624),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_01007_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(net5534),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_03379_),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(_00929_),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(net5825),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(_03067_),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_00714_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(net1751),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net7489),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_03537_),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(_01104_),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(net5811),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(net5813),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_00713_),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(net6537),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(net6539),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(_01055_),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(net6640),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(_04306_),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net4562),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_01352_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(net6602),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(net6604),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(_00589_),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(net6779),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(net6781),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_01036_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(net6002),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_03349_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(_00907_),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net7862),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(net6610),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(_03110_),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_00749_),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(net6672),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(net6674),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(_01046_),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(net5993),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(_03346_),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_00904_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(net5539),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net4971),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_03376_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(_00926_),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(net6590),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(_04297_),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_01360_),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(net6543),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_03393_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(_00940_),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(net6628),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(net6630),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net4973),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_01008_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(net5629),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(net5631),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(_01472_),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\rbzero.pov.spi_buffer[17] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(net1706),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_03012_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(_00664_),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(net6606),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(net6608),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net4979),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_01540_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(net6849),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(net6851),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(_01045_),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(net6745),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(net6747),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_01079_),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(net5569),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_03384_),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(_00934_),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net4981),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(net6676),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(net6678),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_01271_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(net6696),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_03446_),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(_00980_),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(net6941),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(net6943),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_01054_),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(net3905),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net8096),
    .X(net652));
 sky130_fd_sc_hd__buf_2 hold1250 (.A(_03387_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(_03401_),
    .X(net1778));
 sky130_fd_sc_hd__buf_2 hold1252 (.A(_03402_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(_03418_),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_00959_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(net6722),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(net6724),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(_01367_),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(net6600),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(_03827_),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net4425),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_01265_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(net3226),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_03048_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(_00696_),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(net8331),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(_08064_),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(net4333),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(net6358),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(net6360),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(_01470_),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net8297),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(net6656),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(net6658),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_01302_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(net6531),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_03465_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(_00997_),
    .X(net1802));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1276 (.A(net8152),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(net5537),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(net6592),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(net6594),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net7211),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(_01398_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(net1865),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_03599_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(_01161_),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(net6519),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(net6521),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_00981_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(net7311),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(_03518_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(_01086_),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net5641),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_2 hold1290 (.A(net8162),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(net5528),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(net6803),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(net6805),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(_01078_),
    .X(net1821));
 sky130_fd_sc_hd__buf_1 hold1295 (.A(net5595),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(net5597),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(net6801),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(_04436_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(_01042_),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net5643),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(net6636),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(net6638),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_01286_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(net7521),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(_03157_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(net4394),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(net6650),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(net6652),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(_01502_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\rbzero.tex_b0[0] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net4983),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(net5567),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(_01022_),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(net6714),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(net6716),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(_01552_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(net7102),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(_04110_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(_01529_),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(net6839),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(net6841),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net4985),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(_01496_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(net6668),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(net6670),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(_01511_),
    .X(net1850));
 sky130_fd_sc_hd__buf_1 hold1324 (.A(net8147),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(net5564),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(net6734),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(net6736),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_01504_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(net3018),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net6051),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(_03527_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(_01095_),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(net6557),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(_02495_),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_00583_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(net6680),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_02997_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(_00650_),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\rbzero.pov.mosi_buffer[0] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(net1808),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net6053),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(_03598_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(_01160_),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(net7509),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(net6666),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(_01159_),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(net6704),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(_04304_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(_01354_),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(net6706),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(net6708),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_01283_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(_00665_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(net3769),
    .X(net1878));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1352 (.A(_02471_),
    .X(net1879));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1353 (.A(_02473_),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(_03397_),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(_03398_),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(_03399_),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(_00943_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(net6743),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(_03570_),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net7464),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_01134_),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(net6865),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_04356_),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(_01307_),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(net6632),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(net6634),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_01346_),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(net2816),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_04126_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(_01514_),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_03693_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(net6829),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(net6831),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_01050_),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(net6761),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(_04275_),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(_01380_),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(net6726),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(net6728),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(_00984_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(net5749),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net4437),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(_03045_),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(_00694_),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(net6867),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(net6869),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(_01034_),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(net6751),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(_04079_),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(_01554_),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(net7142),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(_03022_),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net5032),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(_00673_),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(net5608),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(net5610),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(net6775),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(net6777),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(_01358_),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(net6646),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(_03443_),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(_00977_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(net6833),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net5034),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(_04163_),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(_01481_),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(net7024),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(net7026),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_01060_),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(net6877),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(_03037_),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(_00686_),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(net6811),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(net6813),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net4991),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_01446_),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(net2718),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_04073_),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(_01559_),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(net4824),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(net4826),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(net6968),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(net6970),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(_01026_),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(net3185),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(net4993),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(_03016_),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(_00667_),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(net5633),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(net5635),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(_01310_),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(net6767),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(net6769),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(_01038_),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(net6765),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(_04351_),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net4996),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_01311_),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(net6927),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(net6929),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(_01536_),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(net6807),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(net6809),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_01425_),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(net7050),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(net7052),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(_01390_),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net4998),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(net6903),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(_04388_),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(_01085_),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(net7002),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(_02999_),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(_00652_),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(net6654),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(_04312_),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_01347_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(net6835),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net8341),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(net6837),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(_01590_),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(net5763),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(net5765),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(_00717_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(net6787),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(net6789),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(_01066_),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(net6783),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(net6785),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net4322),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(_01432_),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(net2238),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(net5593),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(_01305_),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(net6753),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(_04078_),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(_01555_),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(net6795),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(_04181_),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(_01464_),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net4802),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(net6799),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(_03405_),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(_00946_),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(net6763),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(_04339_),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(_01322_),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(net3401),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(_03412_),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(_00953_),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(net5553),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net4804),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(net5555),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(net6771),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(_04192_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(_01454_),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(net7160),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(net7162),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(_01576_),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(net6883),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(net6885),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(_01391_),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net7507),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(net7227),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(net7229),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(_01357_),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(net6871),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(_04083_),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(_01550_),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(net7110),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(_04240_),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(_01412_),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(net6939),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net4711),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(_04035_),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(_01594_),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(net6749),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(_04231_),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(_01420_),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(net7128),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(_04153_),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(_01490_),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(net6923),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(net6925),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net6040),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(_01387_),
    .X(net2037));
 sky130_fd_sc_hd__clkbuf_2 hold1511 (.A(net8161),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(net5542),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(net2789),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(net5599),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(_01571_),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(net7018),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(_04132_),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(_01509_),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(net3792),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(net6042),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(_03111_),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(_00750_),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\rbzero.tex_g1[60] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(net6797),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(_01465_),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(net6755),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(_04259_),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(_01394_),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(net6791),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(_03114_),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_01658_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(_00753_),
    .X(net2057));
 sky130_fd_sc_hd__buf_1 hold1531 (.A(net5617),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(net5619),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(net6006),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(net6008),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(_00909_),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(net6893),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(net6895),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(_01328_),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(net7474),
    .X(net2066));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold154 (.A(net8099),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(_03158_),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(net4385),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(net7177),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(_03567_),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_01131_),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(net6931),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(net6933),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(_01030_),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(net6067),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(net6069),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net4601),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(_01010_),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\rbzero.pov.ready_buffer[14] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(net628),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(_03009_),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_00661_),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(net6945),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(_04389_),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(_01084_),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(net6773),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(_04230_),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(net7418),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_01421_),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(net2973),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(_03041_),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(_00690_),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(net6702),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(_04148_),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(_01494_),
    .X(net2093));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1567 (.A(net7016),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_04139_),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(_01503_),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(net4637),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\rbzero.spi_registers.new_vshift[3] ),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(net1365),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_03392_),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(_00939_),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(net6821),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(net6823),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(_01508_),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(net5612),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_03408_),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(_00949_),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(net5016),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(net6845),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(net6847),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(_01298_),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(net6710),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(net6712),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(_01362_),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(net7100),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(_04326_),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(_01334_),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(net6873),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net5018),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(net6875),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(_01345_),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(net6688),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(net6690),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(_01588_),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(net6962),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(net5545),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(_01479_),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(net7044),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(net7046),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net5012),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_00663_),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(net6879),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(net6881),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(_01579_),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(net6757),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(net6759),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(_01587_),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(net5652),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(net5654),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(_01338_),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net5014),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(net6131),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(net6133),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_01012_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(net6859),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(_04145_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(_01497_),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(net7284),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(net6964),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(_01478_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(net6738),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net5056),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(net6740),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(_00923_),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(net6955),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(net6957),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_01282_),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(net7438),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(net5548),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(_01561_),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(net7298),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(_04142_),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net5058),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(_01500_),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(net6905),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(net6907),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(_01527_),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(net7020),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(_03010_),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(_00662_),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(net7112),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(net7114),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(_01025_),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(net5048),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(net6994),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(net6996),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(_01074_),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(net7118),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(_04443_),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(_01035_),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(net6984),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(_04077_),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_01556_),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(net7104),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net5050),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(_04204_),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(_01444_),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(net3172),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(_03544_),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(_01110_),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(net7495),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(net6793),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(_00754_),
    .X(net2184));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1658 (.A(net8157),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(net5572),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(net8104),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(net7094),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(_04159_),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(_01484_),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(net7174),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(net7176),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(_01152_),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(net5709),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(net5711),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(_00697_),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(net7984),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net4716),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(net4696),
    .X(net2197));
 sky130_fd_sc_hd__buf_1 hold1671 (.A(net5844),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(_02970_),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(net5846),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(net7134),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(_04113_),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(_01526_),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(net7750),
    .X(net2204));
 sky130_fd_sc_hd__clkbuf_4 hold1678 (.A(_02487_),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(net7304),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net5084),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(_00950_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(net7156),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(net7158),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(_01331_),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(net7058),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(net7060),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(_01058_),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(net2631),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(net5590),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(_01309_),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net5086),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(net7070),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(net7072),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(_01366_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(net6682),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(net6684),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(_01273_),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(net6959),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(net6961),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(_00941_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(net6817),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net5004),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(net6819),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(_01466_),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(net6974),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(net6976),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(_01578_),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(net6023),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(_03359_),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(_00915_),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(net7056),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(_04270_),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(net5006),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(_01385_),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\rbzero.tex_b1[27] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(net1988),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(_04359_),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(_01304_),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(net7594),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(net4478),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\rbzero.tex_g1[57] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(net6911),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(_01462_),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(net5028),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(net7008),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(net7010),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(_01522_),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(net5644),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(net5646),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(_01566_),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(net7239),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(_04328_),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(_01332_),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(net6843),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net5030),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(_03368_),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(_00920_),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(net7062),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(_04057_),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(_01574_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(net3025),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(_03525_),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(_01093_),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(net6935),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(_04296_),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(net5076),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(_01361_),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(net6861),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(net6863),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(_00983_),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(net6921),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(_04089_),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(_01545_),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(net6947),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(net6949),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(_01300_),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net5078),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(net5604),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(net5606),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(net6972),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(_04394_),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(_01080_),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(net7166),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(net7168),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(_01382_),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(net7388),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(net5575),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(net5036),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(_01337_),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(net7014),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(_04196_),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(_01452_),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(net7144),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(_04251_),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(_01401_),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(net7148),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(net7150),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(_01492_),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(net5038),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(net6887),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(_04038_),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(_01591_),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(net7315),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(net7317),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(_01365_),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(net2946),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(_04107_),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(_01532_),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(net5672),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(net4975),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(net5674),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(_01292_),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(net7505),
    .X(net2309));
 sky130_fd_sc_hd__clkbuf_2 hold1783 (.A(_03487_),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(_03515_),
    .X(net2311));
 sky130_fd_sc_hd__buf_4 hold1785 (.A(_03516_),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(_03595_),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(_01157_),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(net7022),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(_04452_),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(net4977),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(_01027_),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(net2660),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(_04168_),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(_01476_),
    .X(net2320));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1794 (.A(net5995),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(net5997),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(_00906_),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(net6966),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(_04096_),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(_01538_),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net5068),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(net7066),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(net7068),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(_01525_),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(net3259),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(_03040_),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(_00689_),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(net7400),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(_04346_),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(_01316_),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(net6897),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net5070),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(net6899),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(_01539_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(net6978),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(net6980),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(_01486_),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(net7225),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(net5660),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(_01548_),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(net7331),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(_04441_),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net5040),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(_01037_),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(net6901),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(_04037_),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(_01592_),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(\rbzero.tex_b1[1] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(net5681),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(_01279_),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(net7012),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(_04311_),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(_01348_),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(net5042),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(net7098),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(_04348_),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(_01314_),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(net2647),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(_04391_),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(_01083_),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(\rbzero.pov.ready_buffer[19] ),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(net810),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(_03015_),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(_00666_),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(net5080),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(net7406),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(_04370_),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(_01294_),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(net7323),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(_04092_),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(_01542_),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(net7456),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(net5638),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(_01565_),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\rbzero.tex_g1[44] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net5082),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(net7138),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(_01449_),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(net5665),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(net5667),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(net7247),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(_04417_),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(_01059_),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(net7140),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(_04115_),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(_01524_),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net5052),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(net7203),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(net7205),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(_01073_),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(net7223),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(_04143_),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(_01499_),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(net3066),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(_04032_),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(_01597_),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(net7566),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(net5054),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(_03681_),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(net4285),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(net7048),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(_04241_),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(_01411_),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(net7170),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(net7172),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(_01427_),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(net6917),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(net6919),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(net4987),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(_01501_),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\rbzero.tex_g1[32] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(net6992),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(_01437_),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(net7366),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(_03574_),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(_01137_),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(net6075),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(net6077),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(_01011_),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net4989),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(net7028),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(net7030),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(_01459_),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(net7130),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(net7132),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(_01400_),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(net6913),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(net6915),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(_01510_),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(net4900),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(net5024),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(_03052_),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(_00700_),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(net6718),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(net6720),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(_01442_),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(net7090),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(_04201_),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(_01447_),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(net7276),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(_03112_),
    .X(net2436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(net5026),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(_00751_),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(net7327),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(net7329),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(_01582_),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(net6004),
    .X(net2441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(_03350_),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(_00908_),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(net7199),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(_04120_),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(_01520_),
    .X(net2446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net5064),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(net6937),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(_03366_),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(_00918_),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(net7207),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(_04156_),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(_01487_),
    .X(net2452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(net7032),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(_04271_),
    .X(net2454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(_01384_),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(net6986),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net5066),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(_04425_),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(_01052_),
    .X(net2458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(net7209),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(_04210_),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(_01439_),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(net7350),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(net5663),
    .X(net2463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(_01408_),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(net7191),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(_04076_),
    .X(net2466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net5128),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(_01557_),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(net7537),
    .X(net2468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(_03001_),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(_00654_),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(net7398),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(_04209_),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(_01440_),
    .X(net2473));
 sky130_fd_sc_hd__buf_1 hold1947 (.A(net5621),
    .X(net2474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(net5623),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(net2502),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(net5130),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(_04248_),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(_01404_),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(net7296),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(_04435_),
    .X(net2480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(_01043_),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(net7360),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(_04293_),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(_01364_),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(net6953),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(_03021_),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net5092),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(_00672_),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(net7376),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(net7378),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(_01069_),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(net7193),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(_04303_),
    .X(net2492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(_01355_),
    .X(net2493));
 sky130_fd_sc_hd__buf_1 hold1967 (.A(net5691),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(net5693),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(net6951),
    .X(net2496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(net5094),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(_04046_),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(_01584_),
    .X(net2498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(net7164),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(_04054_),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(_01577_),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(\rbzero.tex_g0[63] ),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(net2476),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(_04247_),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(_01405_),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(net3044),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net5072),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(_03521_),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(_01089_),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(net7038),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(net7040),
    .X(net2510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(_01317_),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(net7241),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(_04397_),
    .X(net2513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(_01077_),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(net7152),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(_04219_),
    .X(net2516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(net5074),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(_01431_),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(net7274),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(_04190_),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(_01456_),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(net7335),
    .X(net2521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(_04224_),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(_01426_),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(net7265),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(_04093_),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(_01541_),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(net5008),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(net7106),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(net7108),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(_01049_),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(net6982),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(_04111_),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(_01528_),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(net7380),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(_04203_),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(_01445_),
    .X(net2535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(net6889),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net5010),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(_04381_),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(_01284_),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(net7362),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(_04403_),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(_01072_),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(net3051),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(_03576_),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(_01139_),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(net7337),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(_04330_),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net5000),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(_01330_),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(net7120),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(_04034_),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(_01595_),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(net7136),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(_04200_),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(_01448_),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(net7195),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(net7197),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(_01319_),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net5002),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(net7382),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(net7384),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(_01295_),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(net6998),
    .X(net2560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(_04062_),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(_01569_),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(net6853),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(net6855),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(_01377_),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(net6990),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net5120),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(_04213_),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(_01436_),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(net7179),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(net7181),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(_01441_),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(net7243),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(net7245),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(_01070_),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(net7290),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2049 (.A(_04261_),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net5122),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2050 (.A(_01392_),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2051 (.A(\rbzero.tex_b1[8] ),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2052 (.A(net6891),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2053 (.A(_01285_),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2054 (.A(net7368),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2055 (.A(net5578),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2056 (.A(_01517_),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2057 (.A(net3213),
    .X(net2584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2058 (.A(_03038_),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2059 (.A(_00687_),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net5096),
    .X(net733));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2060 (.A(net8150),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2061 (.A(net5615),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2062 (.A(net7278),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2063 (.A(_04269_),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2064 (.A(_01386_),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2065 (.A(net7251),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2066 (.A(_04170_),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2067 (.A(_01474_),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2068 (.A(\rbzero.tex_g1[4] ),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2069 (.A(net7352),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net5098),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2070 (.A(_01409_),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2071 (.A(net3815),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2072 (.A(_03411_),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2073 (.A(_00952_),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2074 (.A(net7096),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2075 (.A(_04378_),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2076 (.A(_01287_),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2077 (.A(net7422),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2078 (.A(_04278_),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2079 (.A(_01378_),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(net6124),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2080 (.A(net7201),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2081 (.A(_04430_),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2082 (.A(_01047_),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2083 (.A(net7468),
    .X(net2610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2084 (.A(net7370),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2085 (.A(_01516_),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2086 (.A(net6626),
    .X(net2613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2087 (.A(_04018_),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2088 (.A(_01660_),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2089 (.A(net7189),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(net6126),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2090 (.A(_04282_),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2091 (.A(_01374_),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2092 (.A(net6988),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2093 (.A(_04154_),
    .X(net2620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2094 (.A(_01489_),
    .X(net2621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2095 (.A(net2734),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2096 (.A(net5670),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2097 (.A(_01325_),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2098 (.A(net7221),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2099 (.A(_04147_),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_01106_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2100 (.A(_01495_),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2101 (.A(net3366),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2102 (.A(_03127_),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2103 (.A(net5756),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2104 (.A(\rbzero.tex_b1[31] ),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2105 (.A(net2214),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2106 (.A(_04355_),
    .X(net2633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2107 (.A(_01308_),
    .X(net2634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2108 (.A(net7219),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2109 (.A(_04152_),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net5140),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2110 (.A(_01491_),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2111 (.A(net7292),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2112 (.A(_04226_),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2113 (.A(_01424_),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2114 (.A(net7054),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2115 (.A(_04082_),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2116 (.A(_01551_),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2117 (.A(net3877),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2118 (.A(_03410_),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2119 (.A(_00951_),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net5142),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2120 (.A(\rbzero.tex_b0[61] ),
    .X(net2647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2121 (.A(net2360),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2122 (.A(_04392_),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2123 (.A(_01082_),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2124 (.A(net7249),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2125 (.A(_04222_),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2126 (.A(_01428_),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2127 (.A(net7416),
    .X(net2654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2128 (.A(_04411_),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2129 (.A(_01064_),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(net5156),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2130 (.A(\rbzero.tex_r1[42] ),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2131 (.A(net7064),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2132 (.A(_01575_),
    .X(net2659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2133 (.A(\rbzero.tex_r0[7] ),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2134 (.A(net2318),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2135 (.A(_04167_),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2136 (.A(_01477_),
    .X(net2663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2137 (.A(net7074),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2138 (.A(net7076),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2139 (.A(_01288_),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(net5158),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2140 (.A(net7450),
    .X(net2667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2141 (.A(_04334_),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2142 (.A(_01327_),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2143 (.A(net7253),
    .X(net2670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2144 (.A(net7255),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2145 (.A(_01350_),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2146 (.A(net7390),
    .X(net2673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2147 (.A(_04414_),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2148 (.A(_01062_),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2149 (.A(net7183),
    .X(net2676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(net5100),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2150 (.A(_04121_),
    .X(net2677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2151 (.A(_01519_),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2152 (.A(net7124),
    .X(net2679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2153 (.A(net7126),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2154 (.A(_01040_),
    .X(net2681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2155 (.A(net2844),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2156 (.A(_04319_),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2157 (.A(_01340_),
    .X(net2684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2158 (.A(net7215),
    .X(net2685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2159 (.A(_04254_),
    .X(net2686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net5102),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2160 (.A(_01399_),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2161 (.A(net7122),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2162 (.A(_04045_),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2163 (.A(_01585_),
    .X(net2690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2164 (.A(net7185),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2165 (.A(_04258_),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2166 (.A(_01395_),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2167 (.A(net7305),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2168 (.A(net7307),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2169 (.A(_01296_),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(net8347),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2170 (.A(net5713),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2171 (.A(net5715),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2172 (.A(_01342_),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2173 (.A(net6909),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2174 (.A(_04185_),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2175 (.A(_01461_),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2176 (.A(net5683),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2177 (.A(net5685),
    .X(net2704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2178 (.A(_01280_),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2179 (.A(net7345),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net4336),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2180 (.A(_04347_),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2181 (.A(_01315_),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2182 (.A(net7557),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2183 (.A(_03130_),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2184 (.A(net4316),
    .X(net2711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2185 (.A(net7448),
    .X(net2712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2186 (.A(_03587_),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2187 (.A(_01149_),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2188 (.A(net7313),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2189 (.A(_04310_),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(net6692),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2190 (.A(_01349_),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2191 (.A(\rbzero.tex_r1[25] ),
    .X(net2718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2192 (.A(net1938),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2193 (.A(_04074_),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2194 (.A(_01558_),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2195 (.A(net7231),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2196 (.A(_04289_),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2197 (.A(_01368_),
    .X(net2724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2198 (.A(net7088),
    .X(net2725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2199 (.A(_04420_),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(net4688),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2200 (.A(_01056_),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2201 (.A(net7347),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2202 (.A(_04158_),
    .X(net2729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2203 (.A(_01485_),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2204 (.A(net7233),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2205 (.A(_04281_),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2206 (.A(_01375_),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2207 (.A(\rbzero.tex_b1[47] ),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2208 (.A(net2622),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2209 (.A(_04337_),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(net5020),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2210 (.A(_01324_),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2211 (.A(net7004),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2212 (.A(_04236_),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2213 (.A(_01415_),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2214 (.A(net5729),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2215 (.A(net5731),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2216 (.A(_01549_),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2217 (.A(net7269),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2218 (.A(_04424_),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2219 (.A(_01053_),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net5022),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2220 (.A(net7116),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2221 (.A(_04178_),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2222 (.A(_01467_),
    .X(net2749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2223 (.A(net7078),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2224 (.A(net7080),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2225 (.A(_01450_),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2226 (.A(net5725),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2227 (.A(net5727),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2228 (.A(net7237),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2229 (.A(_04136_),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(net5192),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2230 (.A(_01505_),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2231 (.A(net3439),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2232 (.A(_03042_),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2233 (.A(_00691_),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2234 (.A(net7034),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2235 (.A(net7036),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2236 (.A(_01475_),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2237 (.A(net7553),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2238 (.A(net7420),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2239 (.A(_00649_),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(net5194),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2240 (.A(net2879),
    .X(net2767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2241 (.A(_04087_),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2242 (.A(_01547_),
    .X(net2769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2243 (.A(net7528),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2244 (.A(net1194),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2245 (.A(_03532_),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2246 (.A(_01099_),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2247 (.A(net7294),
    .X(net2774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2248 (.A(_04065_),
    .X(net2775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2249 (.A(_01567_),
    .X(net2776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net5124),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2250 (.A(net7217),
    .X(net2777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2251 (.A(_04344_),
    .X(net2778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2252 (.A(_01318_),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2253 (.A(net7364),
    .X(net2780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2254 (.A(_04044_),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2255 (.A(_01586_),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2256 (.A(net7339),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2257 (.A(_04229_),
    .X(net2784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2258 (.A(_01422_),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2259 (.A(net7286),
    .X(net2786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(net5126),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2260 (.A(net7288),
    .X(net2787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2261 (.A(_01531_),
    .X(net2788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2262 (.A(\rbzero.tex_r1[37] ),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2263 (.A(net2040),
    .X(net2790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2264 (.A(_04061_),
    .X(net2791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2265 (.A(_01570_),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2266 (.A(\rbzero.tex_r0[1] ),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2267 (.A(net5602),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2268 (.A(_01471_),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2269 (.A(net7349),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net8231),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2270 (.A(net975),
    .X(net2797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2271 (.A(_04068_),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2272 (.A(_01564_),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2273 (.A(\rbzero.pov.spi_buffer[48] ),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2274 (.A(net1145),
    .X(net2801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2275 (.A(_03571_),
    .X(net2802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2276 (.A(_01135_),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2277 (.A(net7446),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2278 (.A(_04410_),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2279 (.A(_01065_),
    .X(net2806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(net7926),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2280 (.A(net3076),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2281 (.A(_03534_),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2282 (.A(_01101_),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2283 (.A(net2906),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2284 (.A(_04177_),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2285 (.A(_01468_),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2286 (.A(net7392),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2287 (.A(_04413_),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2288 (.A(_01063_),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2289 (.A(\rbzero.tex_r0[45] ),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(net8191),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2290 (.A(net1894),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2291 (.A(_04125_),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2292 (.A(_01515_),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2293 (.A(net7261),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2294 (.A(net7263),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2295 (.A(_01457_),
    .X(net2822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2296 (.A(net5648),
    .X(net2823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2297 (.A(net5650),
    .X(net2824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2298 (.A(_01306_),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2299 (.A(net7430),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(net7913),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2300 (.A(_04250_),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2301 (.A(_01402_),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2302 (.A(net7559),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2303 (.A(net7466),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2304 (.A(_00702_),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2305 (.A(net7257),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2306 (.A(net7259),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2307 (.A(_01029_),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2308 (.A(net5625),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2309 (.A(net5627),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(net5259),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2310 (.A(_01023_),
    .X(net2837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2311 (.A(net3137),
    .X(net2838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2312 (.A(_03043_),
    .X(net2839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2313 (.A(_00692_),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2314 (.A(net7146),
    .X(net2841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2315 (.A(_04419_),
    .X(net2842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2316 (.A(_01057_),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2317 (.A(\rbzero.tex_b1[63] ),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2318 (.A(net2682),
    .X(net2845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2319 (.A(_04318_),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net5261),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2320 (.A(_01341_),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2321 (.A(\rbzero.tex_g1[11] ),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2322 (.A(net7006),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2323 (.A(_01416_),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2324 (.A(net7235),
    .X(net2851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2325 (.A(_04040_),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2326 (.A(_01589_),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2327 (.A(net7300),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2328 (.A(_04433_),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2329 (.A(_01044_),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(net5116),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2330 (.A(\rbzero.tex_g0[3] ),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2331 (.A(net7213),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2332 (.A(_01344_),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2333 (.A(net3282),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2334 (.A(_03581_),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2335 (.A(_01144_),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2336 (.A(net2926),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2337 (.A(_03064_),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2338 (.A(_00711_),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2339 (.A(net3162),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(net5118),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2340 (.A(_04324_),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2341 (.A(_01336_),
    .X(net2868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2342 (.A(net7541),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2343 (.A(_03531_),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2344 (.A(_01098_),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2345 (.A(net3949),
    .X(net2872));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2346 (.A(_02991_),
    .X(net2873));
 sky130_fd_sc_hd__clkbuf_4 hold2347 (.A(_03047_),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2348 (.A(_03051_),
    .X(net2875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2349 (.A(_00699_),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(net7154),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2350 (.A(net7952),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2351 (.A(net4572),
    .X(net2878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2352 (.A(\rbzero.tex_r1[13] ),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2353 (.A(net2767),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2354 (.A(_04088_),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2355 (.A(_01546_),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2356 (.A(net2977),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2357 (.A(net5587),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2358 (.A(_01291_),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2359 (.A(\rbzero.tex_g0[56] ),
    .X(net2886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net4700),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2360 (.A(net7356),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2361 (.A(_01397_),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2362 (.A(net7424),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2363 (.A(_03602_),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2364 (.A(_01164_),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2365 (.A(net7319),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2366 (.A(_04447_),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2367 (.A(_01032_),
    .X(net2894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2368 (.A(net7374),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2369 (.A(_04455_),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(net5148),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2370 (.A(_01024_),
    .X(net2897));
 sky130_fd_sc_hd__buf_2 hold2371 (.A(net8192),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2372 (.A(net5828),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2373 (.A(net7476),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2374 (.A(net7478),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2375 (.A(_01389_),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2376 (.A(net7454),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2377 (.A(_03584_),
    .X(net2904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2378 (.A(_01146_),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2379 (.A(\rbzero.tex_g1[63] ),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(net5150),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2380 (.A(net2810),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2381 (.A(_04176_),
    .X(net2908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2382 (.A(_01469_),
    .X(net2909));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2383 (.A(net8310),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2384 (.A(net7280),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2385 (.A(net7282),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2386 (.A(_01033_),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2387 (.A(net7414),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2388 (.A(_04109_),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2389 (.A(_01530_),
    .X(net2916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(net6083),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2390 (.A(net7386),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2391 (.A(_04439_),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2392 (.A(_01039_),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2393 (.A(net3055),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2394 (.A(_03542_),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2395 (.A(_01108_),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2396 (.A(net7354),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2397 (.A(_04257_),
    .X(net2924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2398 (.A(_01396_),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2399 (.A(\rbzero.pov.spi_buffer[64] ),
    .X(net2926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(net6085),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2400 (.A(net2863),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2401 (.A(_03589_),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2402 (.A(_01151_),
    .X(net2929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2403 (.A(net7341),
    .X(net2930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2404 (.A(_04384_),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2405 (.A(_01281_),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2406 (.A(\rbzero.pov.spi_buffer[38] ),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2407 (.A(net1102),
    .X(net2934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2408 (.A(_03559_),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2409 (.A(_01124_),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_01493_),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2410 (.A(net7343),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2411 (.A(_04341_),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2412 (.A(_01320_),
    .X(net2939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2413 (.A(net3059),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2414 (.A(net5734),
    .X(net2941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2415 (.A(_00705_),
    .X(net2942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2416 (.A(net7408),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2417 (.A(net7410),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2418 (.A(_00658_),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2419 (.A(\rbzero.tex_r0[63] ),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(net5112),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2420 (.A(net2303),
    .X(net2947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2421 (.A(_04106_),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2422 (.A(_01533_),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2423 (.A(net7325),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2424 (.A(_04135_),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2425 (.A(_01506_),
    .X(net2952));
 sky130_fd_sc_hd__buf_2 hold2426 (.A(net7697),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2427 (.A(net7525),
    .X(net2954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2428 (.A(_00933_),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2429 (.A(net3144),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net5114),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2430 (.A(_03004_),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2431 (.A(_00656_),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2432 (.A(net7402),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2433 (.A(_04119_),
    .X(net2960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2434 (.A(_01521_),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2435 (.A(net7458),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2436 (.A(_04429_),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2437 (.A(_01048_),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2438 (.A(net7042),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2439 (.A(_04237_),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net5144),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2440 (.A(_01414_),
    .X(net2967));
 sky130_fd_sc_hd__buf_1 hold2441 (.A(net5721),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2442 (.A(net5723),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2443 (.A(net7000),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2444 (.A(_04214_),
    .X(net2971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2445 (.A(_01435_),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2446 (.A(\rbzero.pov.spi_buffer[43] ),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2447 (.A(net2088),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2448 (.A(_03566_),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2449 (.A(_01130_),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(net5146),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2450 (.A(\rbzero.tex_b1[13] ),
    .X(net2977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2451 (.A(net2883),
    .X(net2978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2452 (.A(_04374_),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2453 (.A(_01290_),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2454 (.A(net7086),
    .X(net2981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2455 (.A(_04072_),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2456 (.A(_01560_),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2457 (.A(net7267),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2458 (.A(_04050_),
    .X(net2985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2459 (.A(_01580_),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(net5132),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2460 (.A(net7404),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2461 (.A(_04399_),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2462 (.A(_01075_),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2463 (.A(net5717),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2464 (.A(net5719),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2465 (.A(_01326_),
    .X(net2992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2466 (.A(net7440),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2467 (.A(_04129_),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2468 (.A(_01512_),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2469 (.A(net7428),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net5134),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2470 (.A(_04221_),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2471 (.A(_01429_),
    .X(net2998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2472 (.A(net7426),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2473 (.A(_04188_),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2474 (.A(_01458_),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2475 (.A(net7394),
    .X(net3002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2476 (.A(_03407_),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2477 (.A(_00948_),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2478 (.A(net7412),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2479 (.A(_04451_),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(net7082),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2480 (.A(_01028_),
    .X(net3007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2481 (.A(\rbzero.pov.spi_buffer[67] ),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2482 (.A(net1567),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2483 (.A(_03591_),
    .X(net3010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2484 (.A(_01153_),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2485 (.A(net4906),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2486 (.A(net4684),
    .X(net3013));
 sky130_fd_sc_hd__buf_2 hold2487 (.A(net4511),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2488 (.A(net5897),
    .X(net3015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2489 (.A(_03071_),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(net4448),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2490 (.A(_00718_),
    .X(net3017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2491 (.A(\rbzero.pov.spi_buffer[8] ),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2492 (.A(net1856),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2493 (.A(_03002_),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2494 (.A(_00655_),
    .X(net3021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2495 (.A(net7442),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2496 (.A(_03543_),
    .X(net3023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2497 (.A(_01109_),
    .X(net3024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2498 (.A(\rbzero.pov.spi_buffer[7] ),
    .X(net3025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2499 (.A(net2262),
    .X(net3026));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold250 (.A(net8151),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2500 (.A(_03526_),
    .X(net3027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2501 (.A(_01094_),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2502 (.A(net7472),
    .X(net3029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2503 (.A(_04302_),
    .X(net3030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2504 (.A(_01356_),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2505 (.A(net4061),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2506 (.A(_03113_),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2507 (.A(_00752_),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2508 (.A(net3332),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2509 (.A(_03129_),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(net7934),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2510 (.A(net4310),
    .X(net3037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2511 (.A(net6060),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2512 (.A(_03056_),
    .X(net3039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2513 (.A(_00704_),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2514 (.A(net5862),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2515 (.A(_03116_),
    .X(net3042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2516 (.A(_00755_),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2517 (.A(net7527),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2518 (.A(net2506),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2519 (.A(_03522_),
    .X(net3046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(net7092),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2520 (.A(_01090_),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2521 (.A(net3198),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2522 (.A(_03601_),
    .X(net3049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2523 (.A(_01163_),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2524 (.A(\rbzero.pov.spi_buffer[52] ),
    .X(net3051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2525 (.A(net2542),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2526 (.A(_03575_),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2527 (.A(_01138_),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2528 (.A(\rbzero.pov.spi_buffer[21] ),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2529 (.A(net2920),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net4515),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2530 (.A(_03017_),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2531 (.A(_00668_),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2532 (.A(\rbzero.pov.spi_buffer[58] ),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2533 (.A(net2940),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2534 (.A(_03582_),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2535 (.A(_01145_),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2536 (.A(net7539),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2537 (.A(_03536_),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2538 (.A(_01103_),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2539 (.A(\rbzero.tex_r1[63] ),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net4851),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2540 (.A(net2393),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2541 (.A(_04033_),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2542 (.A(_01596_),
    .X(net3069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2543 (.A(net7396),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2544 (.A(_04274_),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2545 (.A(_01381_),
    .X(net3072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2546 (.A(net3255),
    .X(net3073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2547 (.A(_03554_),
    .X(net3074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2548 (.A(_01119_),
    .X(net3075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2549 (.A(\rbzero.pov.spi_buffer[15] ),
    .X(net3076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net4853),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2550 (.A(net2807),
    .X(net3077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2551 (.A(_03535_),
    .X(net3078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2552 (.A(_01102_),
    .X(net3079));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2553 (.A(net7612),
    .X(net3080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2554 (.A(_03029_),
    .X(net3081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2555 (.A(_00679_),
    .X(net3082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2556 (.A(net4831),
    .X(net3083));
 sky130_fd_sc_hd__clkbuf_2 hold2557 (.A(_02949_),
    .X(net3084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2558 (.A(_03373_),
    .X(net3085));
 sky130_fd_sc_hd__buf_4 hold2559 (.A(_03374_),
    .X(net3086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net5176),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2560 (.A(_03382_),
    .X(net3087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2561 (.A(_00932_),
    .X(net3088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2562 (.A(net7432),
    .X(net3089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2563 (.A(net7434),
    .X(net3090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2564 (.A(_01370_),
    .X(net3091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2565 (.A(net7321),
    .X(net3092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2566 (.A(_04365_),
    .X(net3093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2567 (.A(_01299_),
    .X(net3094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2568 (.A(net3124),
    .X(net3095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2569 (.A(_03557_),
    .X(net3096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net5178),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2570 (.A(_01122_),
    .X(net3097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2571 (.A(net5744),
    .X(net3098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2572 (.A(_03059_),
    .X(net3099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2573 (.A(_00706_),
    .X(net3100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2574 (.A(net3110),
    .X(net3101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2575 (.A(_03530_),
    .X(net3102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2576 (.A(_01097_),
    .X(net3103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2577 (.A(\rbzero.tex_g1[1] ),
    .X(net3104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2578 (.A(net5701),
    .X(net3105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2579 (.A(_01407_),
    .X(net3106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(net5152),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2580 (.A(net7485),
    .X(net3107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2581 (.A(net7487),
    .X(net3108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2582 (.A(_01372_),
    .X(net3109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2583 (.A(\rbzero.pov.spi_buffer[10] ),
    .X(net3110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2584 (.A(net3101),
    .X(net3111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2585 (.A(_03005_),
    .X(net3112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2586 (.A(_00657_),
    .X(net3113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2587 (.A(net5695),
    .X(net3114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2588 (.A(net5697),
    .X(net3115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2589 (.A(_01562_),
    .X(net3116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net5154),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2590 (.A(net7503),
    .X(net3117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2591 (.A(_04407_),
    .X(net3118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2592 (.A(_01068_),
    .X(net3119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2593 (.A(\rbzero.pov.spi_buffer[54] ),
    .X(net3120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2594 (.A(net1558),
    .X(net3121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2595 (.A(_03578_),
    .X(net3122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2596 (.A(_01141_),
    .X(net3123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2597 (.A(\rbzero.pov.spi_buffer[36] ),
    .X(net3124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2598 (.A(net3095),
    .X(net3125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2599 (.A(_03558_),
    .X(net3126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net5136),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2600 (.A(_01123_),
    .X(net3127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2601 (.A(net7358),
    .X(net3128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2602 (.A(_04049_),
    .X(net3129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2603 (.A(_01581_),
    .X(net3130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2604 (.A(net7460),
    .X(net3131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2605 (.A(net7462),
    .X(net3132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2606 (.A(_00688_),
    .X(net3133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2607 (.A(net7452),
    .X(net3134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2608 (.A(_03569_),
    .X(net3135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2609 (.A(_01133_),
    .X(net3136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net5138),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2610 (.A(\rbzero.pov.spi_buffer[45] ),
    .X(net3137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2611 (.A(net2838),
    .X(net3138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2612 (.A(_03568_),
    .X(net3139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2613 (.A(_01132_),
    .X(net3140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2614 (.A(net5960),
    .X(net3141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2615 (.A(net5962),
    .X(net3142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2616 (.A(_00597_),
    .X(net3143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2617 (.A(\rbzero.pov.spi_buffer[9] ),
    .X(net3144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2618 (.A(net2956),
    .X(net3145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2619 (.A(_03529_),
    .X(net3146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net4886),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2620 (.A(_01096_),
    .X(net3147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2621 (.A(net3194),
    .X(net3148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2622 (.A(_03548_),
    .X(net3149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2623 (.A(_01114_),
    .X(net3150));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2624 (.A(net4304),
    .X(net3151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2625 (.A(net7491),
    .X(net3152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2626 (.A(net7493),
    .X(net3153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2627 (.A(_01417_),
    .X(net3154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2628 (.A(net7497),
    .X(net3155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2629 (.A(_03538_),
    .X(net3156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(net4888),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2630 (.A(_01105_),
    .X(net3157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2631 (.A(\rbzero.pov.spi_buffer[63] ),
    .X(net3158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2632 (.A(net1471),
    .X(net3159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2633 (.A(_03588_),
    .X(net3160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2634 (.A(_01150_),
    .X(net3161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2635 (.A(\rbzero.tex_b1[58] ),
    .X(net3162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2636 (.A(net2866),
    .X(net3163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2637 (.A(_04325_),
    .X(net3164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2638 (.A(_01335_),
    .X(net3165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2639 (.A(net7533),
    .X(net3166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net7187),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2640 (.A(_03564_),
    .X(net3167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2641 (.A(_01128_),
    .X(net3168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2642 (.A(net7372),
    .X(net3169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2643 (.A(_04215_),
    .X(net3170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2644 (.A(_01434_),
    .X(net3171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2645 (.A(\rbzero.pov.spi_buffer[24] ),
    .X(net3172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2646 (.A(net2179),
    .X(net3173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2647 (.A(_03545_),
    .X(net3174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2648 (.A(_01111_),
    .X(net3175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2649 (.A(net7436),
    .X(net3176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net4605),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2650 (.A(_04280_),
    .X(net3177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2651 (.A(_01376_),
    .X(net3178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2652 (.A(net7555),
    .X(net3179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2653 (.A(net7545),
    .X(net3180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2654 (.A(_00675_),
    .X(net3181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2655 (.A(\rbzero.pov.ready_buffer[22] ),
    .X(net3182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2656 (.A(net7444),
    .X(net3183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2657 (.A(_00669_),
    .X(net3184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2658 (.A(\rbzero.pov.spi_buffer[20] ),
    .X(net3185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2659 (.A(net1946),
    .X(net3186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(net5160),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2660 (.A(_03541_),
    .X(net3187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2661 (.A(_01107_),
    .X(net3188));
 sky130_fd_sc_hd__buf_1 hold2662 (.A(net5738),
    .X(net3189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2663 (.A(net5740),
    .X(net3190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2664 (.A(net3236),
    .X(net3191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2665 (.A(net5792),
    .X(net3192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2666 (.A(_00716_),
    .X(net3193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2667 (.A(\rbzero.pov.spi_buffer[27] ),
    .X(net3194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2668 (.A(net3148),
    .X(net3195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2669 (.A(_03023_),
    .X(net3196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(net5162),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2670 (.A(_00674_),
    .X(net3197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2671 (.A(\rbzero.pov.ss_buffer[0] ),
    .X(net3198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2672 (.A(net3048),
    .X(net3199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2673 (.A(_03600_),
    .X(net3200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2674 (.A(_01162_),
    .X(net3201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2675 (.A(net7499),
    .X(net3202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2676 (.A(_04267_),
    .X(net3203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2677 (.A(_01388_),
    .X(net3204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2678 (.A(net7966),
    .X(net3205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2679 (.A(net4578),
    .X(net3206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(net5104),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2680 (.A(net3301),
    .X(net3207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2681 (.A(_03027_),
    .X(net3208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2682 (.A(_00677_),
    .X(net3209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2683 (.A(net3328),
    .X(net3210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2684 (.A(_03519_),
    .X(net3211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2685 (.A(_01087_),
    .X(net3212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2686 (.A(\rbzero.pov.spi_buffer[40] ),
    .X(net3213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2687 (.A(net2584),
    .X(net3214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2688 (.A(_03563_),
    .X(net3215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2689 (.A(_01127_),
    .X(net3216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(net5106),
    .X(net796));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2690 (.A(net5977),
    .X(net3217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2691 (.A(net5979),
    .X(net3218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2692 (.A(_00924_),
    .X(net3219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2693 (.A(net7501),
    .X(net3220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2694 (.A(_03603_),
    .X(net3221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2695 (.A(_01165_),
    .X(net3222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2696 (.A(net3311),
    .X(net3223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2697 (.A(_03055_),
    .X(net3224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2698 (.A(_00703_),
    .X(net3225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2699 (.A(\rbzero.pov.spi_buffer[49] ),
    .X(net3226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(net5108),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2700 (.A(net1788),
    .X(net3227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2701 (.A(_03573_),
    .X(net3228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2702 (.A(_01136_),
    .X(net3229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2703 (.A(net3350),
    .X(net3230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2704 (.A(_03520_),
    .X(net3231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2705 (.A(_01088_),
    .X(net3232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2706 (.A(net7515),
    .X(net3233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2707 (.A(_03552_),
    .X(net3234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2708 (.A(_01117_),
    .X(net3235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2709 (.A(\rbzero.pov.spi_buffer[69] ),
    .X(net3236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net5110),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2710 (.A(net3191),
    .X(net3237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2711 (.A(_03594_),
    .X(net3238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2712 (.A(_01156_),
    .X(net3239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2713 (.A(\rbzero.tex_r1[39] ),
    .X(net3240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2714 (.A(net5678),
    .X(net3241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2715 (.A(_01572_),
    .X(net3242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2716 (.A(net7529),
    .X(net3243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2717 (.A(_04367_),
    .X(net3244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2718 (.A(_01297_),
    .X(net3245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2719 (.A(net7531),
    .X(net3246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(net5239),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2720 (.A(_04285_),
    .X(net3247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2721 (.A(_01371_),
    .X(net3248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2722 (.A(net7513),
    .X(net3249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2723 (.A(_04233_),
    .X(net3250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2724 (.A(_01418_),
    .X(net3251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2725 (.A(net7470),
    .X(net3252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2726 (.A(_03044_),
    .X(net3253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2727 (.A(_00693_),
    .X(net3254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2728 (.A(\rbzero.pov.spi_buffer[32] ),
    .X(net3255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2729 (.A(net3073),
    .X(net3256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(net5241),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2730 (.A(_03553_),
    .X(net3257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2731 (.A(_01118_),
    .X(net3258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2732 (.A(\rbzero.pov.spi_buffer[42] ),
    .X(net3259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2733 (.A(net2330),
    .X(net3260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2734 (.A(_03565_),
    .X(net3261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2735 (.A(_01129_),
    .X(net3262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2736 (.A(net7483),
    .X(net3263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2737 (.A(_04288_),
    .X(net3264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2738 (.A(_01369_),
    .X(net3265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2739 (.A(net5848),
    .X(net3266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(net5267),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2740 (.A(_03065_),
    .X(net3267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2741 (.A(_00712_),
    .X(net3268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2742 (.A(net7535),
    .X(net3269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2743 (.A(_03062_),
    .X(net3270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2744 (.A(_00709_),
    .X(net3271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2745 (.A(\rbzero.pov.spi_buffer[34] ),
    .X(net3272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2746 (.A(net1358),
    .X(net3273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2747 (.A(_03031_),
    .X(net3274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2748 (.A(_00681_),
    .X(net3275));
 sky130_fd_sc_hd__buf_1 hold2749 (.A(net7549),
    .X(net3276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net5269),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2750 (.A(_03028_),
    .X(net3277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2751 (.A(_00678_),
    .X(net3278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2752 (.A(net5867),
    .X(net3279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2753 (.A(_03068_),
    .X(net3280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2754 (.A(_00715_),
    .X(net3281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2755 (.A(\rbzero.pov.spi_buffer[57] ),
    .X(net3282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2756 (.A(net2860),
    .X(net3283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2757 (.A(_03580_),
    .X(net3284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2758 (.A(_01143_),
    .X(net3285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2759 (.A(net7519),
    .X(net3286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(net6091),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2760 (.A(_03586_),
    .X(net3287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2761 (.A(_01148_),
    .X(net3288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2762 (.A(net7547),
    .X(net3289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2763 (.A(_03020_),
    .X(net3290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2764 (.A(_00671_),
    .X(net3291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2765 (.A(net3341),
    .X(net3292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2766 (.A(_03026_),
    .X(net3293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2767 (.A(_00676_),
    .X(net3294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2768 (.A(net7990),
    .X(net3295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2769 (.A(net4739),
    .X(net3296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(net6093),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2770 (.A(\rbzero.pov.spi_buffer[35] ),
    .X(net3297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2771 (.A(net1646),
    .X(net3298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2772 (.A(_03556_),
    .X(net3299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2773 (.A(_01121_),
    .X(net3300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2774 (.A(\rbzero.pov.spi_buffer[30] ),
    .X(net3301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2775 (.A(net3207),
    .X(net3302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2776 (.A(_03551_),
    .X(net3303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2777 (.A(_01116_),
    .X(net3304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2778 (.A(net7271),
    .X(net3305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2779 (.A(_03604_),
    .X(net3306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_01393_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2780 (.A(_01166_),
    .X(net3307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2781 (.A(net5924),
    .X(net3308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2782 (.A(net5926),
    .X(net3309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2783 (.A(_00625_),
    .X(net3310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2784 (.A(\rbzero.pov.spi_buffer[56] ),
    .X(net3311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2785 (.A(net3223),
    .X(net3312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2786 (.A(_03579_),
    .X(net3313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2787 (.A(_01142_),
    .X(net3314));
 sky130_fd_sc_hd__clkbuf_2 hold2788 (.A(net5858),
    .X(net3315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2789 (.A(net5860),
    .X(net3316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net5243),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 hold2790 (.A(net7780),
    .X(net3317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2791 (.A(net4364),
    .X(net3318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2792 (.A(\rbzero.pov.spi_buffer[39] ),
    .X(net3319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2793 (.A(net1151),
    .X(net3320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2794 (.A(_03562_),
    .X(net3321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2795 (.A(_01126_),
    .X(net3322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2796 (.A(net5770),
    .X(net3323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2797 (.A(_03050_),
    .X(net3324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2798 (.A(_00698_),
    .X(net3325));
 sky130_fd_sc_hd__clkbuf_4 hold2799 (.A(net7689),
    .X(net3326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(net5245),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2800 (.A(net4903),
    .X(net3327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2801 (.A(\rbzero.pov.spi_buffer[0] ),
    .X(net3328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2802 (.A(net3210),
    .X(net3329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2803 (.A(_02994_),
    .X(net3330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2804 (.A(_00647_),
    .X(net3331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2805 (.A(\rbzero.spi_registers.new_other[7] ),
    .X(net3332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2806 (.A(net3035),
    .X(net3333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2807 (.A(_03381_),
    .X(net3334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2808 (.A(_00931_),
    .X(net3335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2809 (.A(net4185),
    .X(net3336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(net5172),
    .X(net808));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2810 (.A(net4187),
    .X(net3337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2811 (.A(net5985),
    .X(net3338));
 sky130_fd_sc_hd__clkbuf_2 hold2812 (.A(net5767),
    .X(net3339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2813 (.A(net4444),
    .X(net3340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2814 (.A(\rbzero.pov.spi_buffer[29] ),
    .X(net3341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2815 (.A(net3292),
    .X(net3342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2816 (.A(_03549_),
    .X(net3343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2817 (.A(_01115_),
    .X(net3344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2818 (.A(net7604),
    .X(net3345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2819 (.A(net7511),
    .X(net3346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net5174),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2820 (.A(_00719_),
    .X(net3347));
 sky130_fd_sc_hd__clkbuf_2 hold2821 (.A(net7764),
    .X(net3348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2822 (.A(net5838),
    .X(net3349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2823 (.A(\rbzero.pov.spi_buffer[1] ),
    .X(net3350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2824 (.A(net3230),
    .X(net3351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2825 (.A(_02995_),
    .X(net3352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2826 (.A(_00648_),
    .X(net3353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2827 (.A(net4926),
    .X(net3354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2828 (.A(net4745),
    .X(net3355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2829 (.A(net7517),
    .X(net3356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net2363),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2830 (.A(_04162_),
    .X(net3357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2831 (.A(_01482_),
    .X(net3358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2832 (.A(net7968),
    .X(net3359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2833 (.A(net4753),
    .X(net3360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2834 (.A(\rbzero.pov.ready_buffer[36] ),
    .X(net3361));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2835 (.A(net1026),
    .X(net3362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2836 (.A(_03033_),
    .X(net3363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2837 (.A(_00683_),
    .X(net3364));
 sky130_fd_sc_hd__buf_2 hold2838 (.A(net4614),
    .X(net3365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2839 (.A(\rbzero.spi_registers.new_other[6] ),
    .X(net3366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(net4556),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2840 (.A(net2628),
    .X(net3367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2841 (.A(_03380_),
    .X(net3368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2842 (.A(_00930_),
    .X(net3369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2843 (.A(net5886),
    .X(net3370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2844 (.A(net5888),
    .X(net3371));
 sky130_fd_sc_hd__buf_2 hold2845 (.A(net7767),
    .X(net3372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2846 (.A(net5752),
    .X(net3373));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2847 (.A(net7728),
    .X(net3374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2848 (.A(_03138_),
    .X(net3375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2849 (.A(_03400_),
    .X(net3376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(net5168),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2850 (.A(_00944_),
    .X(net3377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2851 (.A(net7936),
    .X(net3378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2852 (.A(net4680),
    .X(net3379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2853 (.A(net7994),
    .X(net3380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2854 (.A(net4676),
    .X(net3381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2855 (.A(net8345),
    .X(net3382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2856 (.A(net4544),
    .X(net3383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2857 (.A(net7972),
    .X(net3384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2858 (.A(net4548),
    .X(net3385));
 sky130_fd_sc_hd__clkbuf_1 hold2859 (.A(net8251),
    .X(net3386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(net5170),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2860 (.A(net5747),
    .X(net3387));
 sky130_fd_sc_hd__clkbuf_2 hold2861 (.A(net8313),
    .X(net3388));
 sky130_fd_sc_hd__clkbuf_2 hold2862 (.A(net5914),
    .X(net3389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2863 (.A(net4456),
    .X(net3390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2864 (.A(net8316),
    .X(net3391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2865 (.A(net7986),
    .X(net3392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2866 (.A(net4552),
    .X(net3393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2867 (.A(net3694),
    .X(net3394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2868 (.A(_03075_),
    .X(net3395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2869 (.A(net4064),
    .X(net3396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(net5303),
    .X(net814));
 sky130_fd_sc_hd__buf_2 hold2870 (.A(_03077_),
    .X(net3397));
 sky130_fd_sc_hd__buf_4 hold2871 (.A(_03089_),
    .X(net3398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2872 (.A(_03092_),
    .X(net3399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2873 (.A(_00733_),
    .X(net3400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2874 (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .X(net3401));
 sky130_fd_sc_hd__buf_2 hold2875 (.A(net2003),
    .X(net3402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2876 (.A(_03088_),
    .X(net3403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2877 (.A(_00730_),
    .X(net3404));
 sky130_fd_sc_hd__clkbuf_2 hold2878 (.A(net4338),
    .X(net3405));
 sky130_fd_sc_hd__clkbuf_2 hold2879 (.A(net7906),
    .X(net3406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net5305),
    .X(net815));
 sky130_fd_sc_hd__buf_1 hold2880 (.A(net8171),
    .X(net3407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2881 (.A(net4627),
    .X(net3408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2882 (.A(net4916),
    .X(net3409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2883 (.A(net4509),
    .X(net3410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2884 (.A(net5834),
    .X(net3411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2885 (.A(_03061_),
    .X(net3412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2886 (.A(_00708_),
    .X(net3413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2887 (.A(net7572),
    .X(net3414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2888 (.A(_03672_),
    .X(net3415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2889 (.A(net4345),
    .X(net3416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net7333),
    .X(net816));
 sky130_fd_sc_hd__buf_2 hold2890 (.A(net5928),
    .X(net3417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2891 (.A(_09095_),
    .X(net3418));
 sky130_fd_sc_hd__buf_2 hold2892 (.A(net5903),
    .X(net3419));
 sky130_fd_sc_hd__buf_1 hold2893 (.A(_09210_),
    .X(net3420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2894 (.A(net7992),
    .X(net3421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2895 (.A(net4707),
    .X(net3422));
 sky130_fd_sc_hd__clkbuf_2 hold2896 (.A(net4360),
    .X(net3423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2897 (.A(net4911),
    .X(net3424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2898 (.A(net4692),
    .X(net3425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2899 (.A(net7877),
    .X(net3426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(net4596),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2900 (.A(net7938),
    .X(net3427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2901 (.A(net4899),
    .X(net3428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2902 (.A(net4731),
    .X(net3429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2903 (.A(net8374),
    .X(net3430));
 sky130_fd_sc_hd__clkbuf_4 hold2904 (.A(net7700),
    .X(net3431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2905 (.A(net5900),
    .X(net3432));
 sky130_fd_sc_hd__clkbuf_2 hold2906 (.A(net8206),
    .X(net3433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2907 (.A(net4329),
    .X(net3434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2908 (.A(\rbzero.pov.ready_buffer[37] ),
    .X(net3435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2909 (.A(net7659),
    .X(net3436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(net5247),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2910 (.A(_03717_),
    .X(net3437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2911 (.A(_01201_),
    .X(net3438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2912 (.A(\rbzero.pov.ready_buffer[44] ),
    .X(net3439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2913 (.A(net2758),
    .X(net3440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2914 (.A(_03664_),
    .X(net3441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2915 (.A(net5930),
    .X(net3442));
 sky130_fd_sc_hd__clkbuf_4 hold2916 (.A(net8236),
    .X(net3443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2917 (.A(net5870),
    .X(net3444));
 sky130_fd_sc_hd__clkbuf_4 hold2918 (.A(net8224),
    .X(net3445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2919 (.A(net5773),
    .X(net3446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(net5249),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2920 (.A(net7574),
    .X(net3447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2921 (.A(net7576),
    .X(net3448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2922 (.A(_00617_),
    .X(net3449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2923 (.A(net7852),
    .X(net3450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2924 (.A(net3974),
    .X(net3451));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2925 (.A(_04654_),
    .X(net3452));
 sky130_fd_sc_hd__buf_2 hold2926 (.A(_08378_),
    .X(net3453));
 sky130_fd_sc_hd__clkbuf_2 hold2927 (.A(_08421_),
    .X(net3454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2928 (.A(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(net3455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2929 (.A(net4839),
    .X(net3456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(net5223),
    .X(net820));
 sky130_fd_sc_hd__buf_2 hold2930 (.A(net8213),
    .X(net3457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2931 (.A(net5852),
    .X(net3458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2932 (.A(net7867),
    .X(net3459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2933 (.A(net7870),
    .X(net3460));
 sky130_fd_sc_hd__buf_2 hold2934 (.A(net7770),
    .X(net3461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2935 (.A(net4493),
    .X(net3462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2936 (.A(\rbzero.row_render.size[2] ),
    .X(net3715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2937 (.A(net5776),
    .X(net3464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2938 (.A(net5778),
    .X(net3465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2939 (.A(net8321),
    .X(net3466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(net5225),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2940 (.A(net8382),
    .X(net3467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2941 (.A(net8057),
    .X(net3468));
 sky130_fd_sc_hd__buf_2 hold2942 (.A(\rbzero.debug_overlay.playerY[5] ),
    .X(net3469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2943 (.A(net5761),
    .X(net3470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2944 (.A(_01196_),
    .X(net3471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2945 (.A(net7941),
    .X(net3472));
 sky130_fd_sc_hd__clkbuf_4 hold2946 (.A(net7634),
    .X(net3473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2947 (.A(net4376),
    .X(net3474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2948 (.A(net7916),
    .X(net3475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2949 (.A(net7998),
    .X(net3476));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold295 (.A(net8196),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2950 (.A(net4662),
    .X(net3477));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2951 (.A(net7578),
    .X(net3478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2952 (.A(_03100_),
    .X(net3479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2953 (.A(_00741_),
    .X(net3480));
 sky130_fd_sc_hd__clkbuf_2 hold2954 (.A(net7596),
    .X(net3481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2955 (.A(net7580),
    .X(net3482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2956 (.A(_00742_),
    .X(net3483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2957 (.A(net7831),
    .X(net3484));
 sky130_fd_sc_hd__clkbuf_2 hold2958 (.A(net7693),
    .X(net3485));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2959 (.A(_02967_),
    .X(net3486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(net8023),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2960 (.A(net5865),
    .X(net3487));
 sky130_fd_sc_hd__clkbuf_2 hold2961 (.A(net8319),
    .X(net3488));
 sky130_fd_sc_hd__clkbuf_4 hold2962 (.A(net8219),
    .X(net3489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2963 (.A(net4619),
    .X(net3490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2964 (.A(net8324),
    .X(net3491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2965 (.A(net7903),
    .X(net3492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2966 (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(net3493));
 sky130_fd_sc_hd__clkbuf_4 hold2967 (.A(_02552_),
    .X(net3494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2968 (.A(_03760_),
    .X(net3495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2969 (.A(_03761_),
    .X(net3496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net5211),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2970 (.A(_01226_),
    .X(net3497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2972 (.A(net5795),
    .X(net3499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2973 (.A(net5797),
    .X(net3500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2974 (.A(net8358),
    .X(net3501));
 sky130_fd_sc_hd__clkbuf_2 hold2975 (.A(net1585),
    .X(net3502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2977 (.A(net7626),
    .X(net3504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2978 (.A(_03734_),
    .X(net3505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2979 (.A(_01210_),
    .X(net3506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(net5213),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2980 (.A(net7797),
    .X(net3507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2981 (.A(net8037),
    .X(net3508));
 sky130_fd_sc_hd__clkbuf_4 hold2982 (.A(net7735),
    .X(net3509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2983 (.A(_03757_),
    .X(net3510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2984 (.A(_03758_),
    .X(net3511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2985 (.A(_01224_),
    .X(net3512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2987 (.A(_02569_),
    .X(net3514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2988 (.A(net4786),
    .X(net3515));
 sky130_fd_sc_hd__buf_1 hold2989 (.A(net5204),
    .X(net3516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(net5060),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 hold2990 (.A(net5913),
    .X(net3517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2991 (.A(_00478_),
    .X(net3518));
 sky130_fd_sc_hd__buf_2 hold2992 (.A(net5931),
    .X(net3519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2993 (.A(_03361_),
    .X(net3520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2994 (.A(_03362_),
    .X(net3521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2995 (.A(_00917_),
    .X(net3522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2997 (.A(net5804),
    .X(net3524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2998 (.A(net5806),
    .X(net3525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(net5062),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3000 (.A(net5808),
    .X(net3527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3001 (.A(net5810),
    .X(net3528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3002 (.A(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(net3529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3003 (.A(net4829),
    .X(net3530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3004 (.A(net7919),
    .X(net3531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3005 (.A(net7789),
    .X(net3532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3007 (.A(_02808_),
    .X(net3534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3008 (.A(net4773),
    .X(net3535));
 sky130_fd_sc_hd__clkbuf_4 hold3009 (.A(net8226),
    .X(net3536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(net5180),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3010 (.A(net5819),
    .X(net3537));
 sky130_fd_sc_hd__clkbuf_2 hold3011 (.A(net4527),
    .X(net3538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3012 (.A(_03769_),
    .X(net3539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3013 (.A(_03770_),
    .X(net3540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3014 (.A(_01233_),
    .X(net3541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3015 (.A(net7848),
    .X(net3542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3016 (.A(net7586),
    .X(net3543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3017 (.A(_03622_),
    .X(net3544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3018 (.A(_03623_),
    .X(net3545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3019 (.A(net5905),
    .X(net3546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(net5182),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3020 (.A(net7721),
    .X(net3547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3021 (.A(_03327_),
    .X(net3548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3022 (.A(_03328_),
    .X(net3549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3023 (.A(_00893_),
    .X(net3550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3024 (.A(net8380),
    .X(net3551));
 sky130_fd_sc_hd__clkbuf_4 hold3025 (.A(\rbzero.debug_overlay.playerY[4] ),
    .X(net3552));
 sky130_fd_sc_hd__buf_1 hold3026 (.A(_04685_),
    .X(net3553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3027 (.A(net6062),
    .X(net3554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3028 (.A(_01195_),
    .X(net3555));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3029 (.A(net7588),
    .X(net3556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(net5403),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3030 (.A(net7590),
    .X(net3557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3031 (.A(_00738_),
    .X(net3558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3032 (.A(net4873),
    .X(net3559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3033 (.A(net4672),
    .X(net3560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3034 (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .X(net3561));
 sky130_fd_sc_hd__buf_2 hold3035 (.A(net1655),
    .X(net3562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3036 (.A(_03094_),
    .X(net3563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3037 (.A(_00735_),
    .X(net3564));
 sky130_fd_sc_hd__clkbuf_4 hold3038 (.A(net7737),
    .X(net3565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3039 (.A(_03750_),
    .X(net3566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(net5405),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3040 (.A(_03751_),
    .X(net3567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3041 (.A(_01219_),
    .X(net3568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3042 (.A(net7736),
    .X(net3569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3043 (.A(_03313_),
    .X(net3570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3044 (.A(_03314_),
    .X(net3571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3045 (.A(_00886_),
    .X(net3572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3046 (.A(net8391),
    .X(net3573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3047 (.A(net7880),
    .X(net3574));
 sky130_fd_sc_hd__clkbuf_4 hold3048 (.A(net7739),
    .X(net3575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3049 (.A(_03773_),
    .X(net3576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net5327),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3050 (.A(_03774_),
    .X(net3577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3051 (.A(_01235_),
    .X(net3578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3053 (.A(net7642),
    .X(net3580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3054 (.A(_03736_),
    .X(net3581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3055 (.A(_01211_),
    .X(net3582));
 sky130_fd_sc_hd__clkbuf_2 hold3056 (.A(net7600),
    .X(net3583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3057 (.A(net7598),
    .X(net3584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3058 (.A(_00743_),
    .X(net3585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3059 (.A(net8349),
    .X(net3586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(net5329),
    .X(net833));
 sky130_fd_sc_hd__buf_1 hold3060 (.A(net8343),
    .X(net3587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3061 (.A(_02458_),
    .X(net3588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3062 (.A(_02464_),
    .X(net3589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3063 (.A(_02465_),
    .X(net3590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3064 (.A(_02466_),
    .X(net3591));
 sky130_fd_sc_hd__buf_2 hold3065 (.A(net7620),
    .X(net3592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3066 (.A(_03096_),
    .X(net3593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3067 (.A(_00737_),
    .X(net3594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3068 (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .X(net3595));
 sky130_fd_sc_hd__buf_2 hold3069 (.A(net1541),
    .X(net3596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(net8203),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3070 (.A(_03093_),
    .X(net3597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3071 (.A(_00734_),
    .X(net3598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3072 (.A(net7827),
    .X(net3599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3073 (.A(net8329),
    .X(net3600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3074 (.A(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(net3601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3075 (.A(net6047),
    .X(net3602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3076 (.A(_00637_),
    .X(net3603));
 sky130_fd_sc_hd__buf_2 hold3077 (.A(\rbzero.wall_tracer.rayAddendX[2] ),
    .X(net3604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3078 (.A(net5971),
    .X(net3605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3079 (.A(_00603_),
    .X(net3606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(net8020),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3081 (.A(net7652),
    .X(net3608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3082 (.A(_03721_),
    .X(net3609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3083 (.A(_01203_),
    .X(net3610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3084 (.A(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(net3611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3085 (.A(net5956),
    .X(net3612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3086 (.A(_00639_),
    .X(net3613));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3087 (.A(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(net3614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3088 (.A(_02680_),
    .X(net3615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3089 (.A(net4870),
    .X(net3616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net7084),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3090 (.A(net8327),
    .X(net3617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3091 (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(net3618));
 sky130_fd_sc_hd__clkbuf_4 hold3092 (.A(_02762_),
    .X(net3619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3093 (.A(_03771_),
    .X(net3620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3094 (.A(_03772_),
    .X(net3621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3095 (.A(_01234_),
    .X(net3622));
 sky130_fd_sc_hd__clkbuf_2 hold3096 (.A(net5942),
    .X(net3623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3097 (.A(net5944),
    .X(net3624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3098 (.A(_00935_),
    .X(net3625));
 sky130_fd_sc_hd__buf_1 hold3099 (.A(net8447),
    .X(net3626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_03159_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3100 (.A(net5959),
    .X(net3627));
 sky130_fd_sc_hd__clkbuf_2 hold3101 (.A(_04655_),
    .X(net3628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3102 (.A(_01623_),
    .X(net3629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3103 (.A(net8395),
    .X(net3630));
 sky130_fd_sc_hd__clkbuf_2 hold3104 (.A(\rbzero.spi_registers.spi_buffer[23] ),
    .X(net3631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3105 (.A(net7602),
    .X(net3632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3106 (.A(_00744_),
    .X(net3633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3108 (.A(net5822),
    .X(net3635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3109 (.A(net5824),
    .X(net3636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(net4358),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 hold3110 (.A(net7929),
    .X(net3637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3112 (.A(_02595_),
    .X(net3639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3113 (.A(net4727),
    .X(net3640));
 sky130_fd_sc_hd__buf_2 hold3114 (.A(net6037),
    .X(net3641));
 sky130_fd_sc_hd__buf_1 hold3115 (.A(_04497_),
    .X(net3642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3116 (.A(net5209),
    .X(net3643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3117 (.A(net7718),
    .X(net3644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3118 (.A(_03330_),
    .X(net3645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3119 (.A(_03331_),
    .X(net3646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(net6425),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3120 (.A(_00895_),
    .X(net3647));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3121 (.A(net7608),
    .X(net3648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3122 (.A(net7610),
    .X(net3649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3123 (.A(_00522_),
    .X(net3650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3124 (.A(net7724),
    .X(net3651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3125 (.A(_03321_),
    .X(net3652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3126 (.A(_03322_),
    .X(net3653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3127 (.A(_00890_),
    .X(net3654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3128 (.A(net7948),
    .X(net3655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3129 (.A(net7729),
    .X(net3656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_03262_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3130 (.A(_03324_),
    .X(net3657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3131 (.A(_03325_),
    .X(net3658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3132 (.A(_00891_),
    .X(net3659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3133 (.A(net8254),
    .X(net3660));
 sky130_fd_sc_hd__clkbuf_4 hold3134 (.A(_05151_),
    .X(net3661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3135 (.A(_03755_),
    .X(net3662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3136 (.A(_03756_),
    .X(net3663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3137 (.A(_01223_),
    .X(net3664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3138 (.A(net8367),
    .X(net3665));
 sky130_fd_sc_hd__clkbuf_2 hold3139 (.A(_02388_),
    .X(net3666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(net4196),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3140 (.A(_02397_),
    .X(net3667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3141 (.A(net4896),
    .X(net3668));
 sky130_fd_sc_hd__clkbuf_2 hold3142 (.A(net1680),
    .X(net3669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3143 (.A(net7732),
    .X(net3670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3144 (.A(_03317_),
    .X(net3671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3145 (.A(_03318_),
    .X(net3672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3146 (.A(_00888_),
    .X(net3673));
 sky130_fd_sc_hd__clkbuf_2 hold3147 (.A(net7614),
    .X(net3674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3148 (.A(net7616),
    .X(net3675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3149 (.A(_00739_),
    .X(net3676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(net5088),
    .X(net842));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3150 (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(net3677));
 sky130_fd_sc_hd__clkbuf_4 hold3151 (.A(_02792_),
    .X(net3678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3152 (.A(_03776_),
    .X(net3679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3153 (.A(_03777_),
    .X(net3680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3154 (.A(_01237_),
    .X(net3681));
 sky130_fd_sc_hd__clkbuf_4 hold3155 (.A(net7704),
    .X(net3682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3156 (.A(_06059_),
    .X(net3683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3157 (.A(net7606),
    .X(net3684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3158 (.A(_01180_),
    .X(net3685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(net5090),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3160 (.A(net7639),
    .X(net3687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3161 (.A(_03730_),
    .X(net3688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3162 (.A(_01208_),
    .X(net3689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3163 (.A(net7480),
    .X(net3690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3164 (.A(net7662),
    .X(net3691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3165 (.A(_03719_),
    .X(net3692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3166 (.A(_01202_),
    .X(net3693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3167 (.A(\rbzero.spi_registers.spi_counter[6] ),
    .X(net3694));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3168 (.A(net3394),
    .X(net3695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3169 (.A(_02988_),
    .X(net3696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net5200),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3170 (.A(_02990_),
    .X(net3697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3171 (.A(_00646_),
    .X(net3698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3172 (.A(net7841),
    .X(net3699));
 sky130_fd_sc_hd__buf_1 hold3173 (.A(_02316_),
    .X(net3700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3174 (.A(_02325_),
    .X(net3701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3175 (.A(net8353),
    .X(net3702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3176 (.A(net7684),
    .X(net3703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3177 (.A(_03490_),
    .X(net3704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3178 (.A(_03494_),
    .X(net3705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3179 (.A(_01016_),
    .X(net3706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(net5202),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3180 (.A(net7672),
    .X(net3707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3181 (.A(_03497_),
    .X(net3708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3182 (.A(net7675),
    .X(net3709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3183 (.A(_01018_),
    .X(net3710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3184 (.A(net7582),
    .X(net3711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3185 (.A(net7645),
    .X(net3712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3186 (.A(_03742_),
    .X(net3713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3187 (.A(_01215_),
    .X(net3714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3189 (.A(net5831),
    .X(net3716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(net5355),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3190 (.A(net5833),
    .X(net3717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3191 (.A(net7931),
    .X(net3718));
 sky130_fd_sc_hd__buf_1 hold3192 (.A(\rbzero.debug_overlay.facingX[-1] ),
    .X(net3719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3193 (.A(net7741),
    .X(net3720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3194 (.A(_03725_),
    .X(net3721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3195 (.A(_01205_),
    .X(net3722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3196 (.A(net8333),
    .X(net3723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3197 (.A(net8335),
    .X(net3724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3198 (.A(net7858),
    .X(net3725));
 sky130_fd_sc_hd__buf_1 hold3199 (.A(net7875),
    .X(net3726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(net5357),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3200 (.A(net7809),
    .X(net3727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3201 (.A(net8082),
    .X(net3728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3202 (.A(net4875),
    .X(net3729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3203 (.A(_02330_),
    .X(net3730));
 sky130_fd_sc_hd__buf_1 hold3204 (.A(_02335_),
    .X(net3731));
 sky130_fd_sc_hd__buf_1 hold3205 (.A(_02345_),
    .X(net3732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3206 (.A(_02347_),
    .X(net3733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3207 (.A(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(net3734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3208 (.A(net6016),
    .X(net3735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3209 (.A(_00609_),
    .X(net3736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(net5383),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3210 (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .X(net3737));
 sky130_fd_sc_hd__buf_2 hold3211 (.A(net1334),
    .X(net3738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3212 (.A(_03095_),
    .X(net3739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3213 (.A(_00736_),
    .X(net3740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3215 (.A(net5841),
    .X(net3742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3216 (.A(net5843),
    .X(net3743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3217 (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .X(net3744));
 sky130_fd_sc_hd__buf_2 hold3218 (.A(net1392),
    .X(net3745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3219 (.A(_03091_),
    .X(net3746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(net5385),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3220 (.A(_00732_),
    .X(net3747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3221 (.A(net7840),
    .X(net3748));
 sky130_fd_sc_hd__clkbuf_2 hold3222 (.A(net3699),
    .X(net3749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3223 (.A(net7983),
    .X(net3750));
 sky130_fd_sc_hd__clkbuf_2 hold3224 (.A(net2196),
    .X(net3751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3226 (.A(net5855),
    .X(net3753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3227 (.A(net5857),
    .X(net3754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3228 (.A(net7956),
    .X(net3755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3229 (.A(net4915),
    .X(net3756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net8078),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_2 hold3230 (.A(net3409),
    .X(net3757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3232 (.A(_02891_),
    .X(net3759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3233 (.A(net4809),
    .X(net3760));
 sky130_fd_sc_hd__clkbuf_2 hold3234 (.A(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(net3761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3235 (.A(_02918_),
    .X(net3762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3236 (.A(net4859),
    .X(net3763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3237 (.A(net7950),
    .X(net3764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3238 (.A(net4910),
    .X(net3765));
 sky130_fd_sc_hd__clkbuf_2 hold3239 (.A(net3424),
    .X(net3766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(net4251),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3240 (.A(net4905),
    .X(net3767));
 sky130_fd_sc_hd__clkbuf_2 hold3241 (.A(net3012),
    .X(net3768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3242 (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .X(net3769));
 sky130_fd_sc_hd__clkbuf_4 hold3243 (.A(net1878),
    .X(net3770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3244 (.A(_03106_),
    .X(net3771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3245 (.A(_00746_),
    .X(net3772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3246 (.A(net4082),
    .X(net3773));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3247 (.A(_04484_),
    .X(net3774));
 sky130_fd_sc_hd__clkbuf_2 hold3248 (.A(_07871_),
    .X(net3775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3249 (.A(net8366),
    .X(net3776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(net5227),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_2 hold3250 (.A(net3665),
    .X(net3777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3251 (.A(\rbzero.wall_tracer.rayAddendX[10] ),
    .X(net3778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3252 (.A(net5953),
    .X(net3779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3253 (.A(_00611_),
    .X(net3780));
 sky130_fd_sc_hd__buf_2 hold3254 (.A(net7664),
    .X(net3781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3255 (.A(net7666),
    .X(net3782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3256 (.A(_00521_),
    .X(net3783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3257 (.A(net4898),
    .X(net3784));
 sky130_fd_sc_hd__clkbuf_2 hold3258 (.A(net3428),
    .X(net3785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3259 (.A(net4925),
    .X(net3786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(net5229),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 hold3260 (.A(net3354),
    .X(net3787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3261 (.A(net8416),
    .X(net3788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3262 (.A(net7965),
    .X(net3789));
 sky130_fd_sc_hd__clkbuf_2 hold3263 (.A(net3205),
    .X(net3790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3264 (.A(net7960),
    .X(net3791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3265 (.A(\rbzero.spi_registers.mosi ),
    .X(net3792));
 sky130_fd_sc_hd__clkbuf_2 hold3266 (.A(net2046),
    .X(net3793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3267 (.A(_03105_),
    .X(net3794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3268 (.A(_00745_),
    .X(net3795));
 sky130_fd_sc_hd__buf_1 hold3269 (.A(net7996),
    .X(net3796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(net5379),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3270 (.A(net4920),
    .X(net3797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3271 (.A(_09860_),
    .X(net3798));
 sky130_fd_sc_hd__buf_1 hold3272 (.A(_09869_),
    .X(net3799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3273 (.A(_09870_),
    .X(net3800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3274 (.A(net7958),
    .X(net3801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3275 (.A(net7967),
    .X(net3802));
 sky130_fd_sc_hd__clkbuf_2 hold3276 (.A(net3359),
    .X(net3803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3277 (.A(net7873),
    .X(net3804));
 sky130_fd_sc_hd__buf_1 hold3278 (.A(_09789_),
    .X(net3805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3279 (.A(net7962),
    .X(net3806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(net5381),
    .X(net855));
 sky130_fd_sc_hd__buf_2 hold3280 (.A(net7668),
    .X(net3807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3281 (.A(net7670),
    .X(net3808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3282 (.A(_00616_),
    .X(net3809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3283 (.A(net7989),
    .X(net3810));
 sky130_fd_sc_hd__clkbuf_2 hold3284 (.A(net3295),
    .X(net3811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3286 (.A(net5873),
    .X(net3813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3287 (.A(net5875),
    .X(net3814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3288 (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .X(net3815));
 sky130_fd_sc_hd__buf_2 hold3289 (.A(net2598),
    .X(net3816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(net5299),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3290 (.A(_03087_),
    .X(net3817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3291 (.A(_00729_),
    .X(net3818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3292 (.A(net7991),
    .X(net3819));
 sky130_fd_sc_hd__clkbuf_2 hold3293 (.A(net3421),
    .X(net3820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3294 (.A(net7872),
    .X(net3821));
 sky130_fd_sc_hd__clkbuf_2 hold3295 (.A(net3804),
    .X(net3822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3296 (.A(net7654),
    .X(net3823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3297 (.A(_03503_),
    .X(net3824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3298 (.A(net7657),
    .X(net3825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3299 (.A(_01020_),
    .X(net3826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(net5301),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3301 (.A(net5883),
    .X(net3828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3302 (.A(net5885),
    .X(net3829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3303 (.A(net8337),
    .X(net3830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3304 (.A(net7964),
    .X(net3831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3305 (.A(net8339),
    .X(net3832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3306 (.A(net7982),
    .X(net3833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3307 (.A(net7993),
    .X(net3834));
 sky130_fd_sc_hd__clkbuf_2 hold3308 (.A(net3380),
    .X(net3835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3309 (.A(net7970),
    .X(net3836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(net5215),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3310 (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .X(net3837));
 sky130_fd_sc_hd__buf_2 hold3311 (.A(net1477),
    .X(net3838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3312 (.A(_03090_),
    .X(net3839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3313 (.A(_00731_),
    .X(net3840));
 sky130_fd_sc_hd__buf_1 hold3314 (.A(net8405),
    .X(net3841));
 sky130_fd_sc_hd__buf_1 hold3315 (.A(net7742),
    .X(net3842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3316 (.A(_03421_),
    .X(net3843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3317 (.A(_03422_),
    .X(net3844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3318 (.A(_00962_),
    .X(net3845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3319 (.A(net7971),
    .X(net3846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(net5217),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_2 hold3320 (.A(net3384),
    .X(net3847));
 sky130_fd_sc_hd__buf_2 hold3321 (.A(net5932),
    .X(net3848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3322 (.A(net5934),
    .X(net3849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3323 (.A(_00614_),
    .X(net3850));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3324 (.A(net3939),
    .X(net3851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3325 (.A(net5896),
    .X(net3852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3326 (.A(_00748_),
    .X(net3853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3327 (.A(net7988),
    .X(net3854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3328 (.A(net7974),
    .X(net3855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3329 (.A(net7976),
    .X(net3856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(net5263),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_2 hold3330 (.A(net7707),
    .X(net3857));
 sky130_fd_sc_hd__buf_1 hold3331 (.A(_04663_),
    .X(net3858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3332 (.A(_09723_),
    .X(net3859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3333 (.A(_00473_),
    .X(net3860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3334 (.A(net7980),
    .X(net3861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3335 (.A(net3876),
    .X(net3862));
 sky130_fd_sc_hd__buf_2 hold3336 (.A(net2644),
    .X(net3863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3337 (.A(_03085_),
    .X(net3864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3338 (.A(_00727_),
    .X(net3865));
 sky130_fd_sc_hd__clkbuf_2 hold3339 (.A(net7628),
    .X(net3866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net5265),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3340 (.A(_03099_),
    .X(net3867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3341 (.A(_00740_),
    .X(net3868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3342 (.A(net7978),
    .X(net3869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3343 (.A(net5921),
    .X(net3870));
 sky130_fd_sc_hd__buf_2 hold3344 (.A(_04473_),
    .X(net3871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3345 (.A(_03994_),
    .X(net3872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3346 (.A(_01625_),
    .X(net3873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3347 (.A(net5584),
    .X(net3874));
 sky130_fd_sc_hd__clkbuf_2 hold3348 (.A(net626),
    .X(net3875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3349 (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .X(net3876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net5184),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3350 (.A(net3862),
    .X(net3877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3351 (.A(_03086_),
    .X(net3878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3352 (.A(_00728_),
    .X(net3879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3354 (.A(net7623),
    .X(net3881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3355 (.A(_03738_),
    .X(net3882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3356 (.A(_01212_),
    .X(net3883));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3357 (.A(net7630),
    .X(net3884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3358 (.A(net7632),
    .X(net3885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3359 (.A(_00623_),
    .X(net3886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net5186),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3360 (.A(net4919),
    .X(net3887));
 sky130_fd_sc_hd__clkbuf_2 hold3361 (.A(net3797),
    .X(net3888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3362 (.A(net8351),
    .X(net3889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3364 (.A(net5891),
    .X(net3891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3365 (.A(net5893),
    .X(net3892));
 sky130_fd_sc_hd__buf_2 hold3366 (.A(net5973),
    .X(net3893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3367 (.A(_02710_),
    .X(net3894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3368 (.A(_00612_),
    .X(net3895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3369 (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .X(net3896));
 sky130_fd_sc_hd__buf_1 hold337 (.A(net8195),
    .X(net864));
 sky130_fd_sc_hd__buf_1 hold3370 (.A(net1621),
    .X(net3897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3371 (.A(_02470_),
    .X(net3898));
 sky130_fd_sc_hd__buf_1 hold3372 (.A(net1622),
    .X(net3899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3373 (.A(_03079_),
    .X(net3900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3374 (.A(_00721_),
    .X(net3901));
 sky130_fd_sc_hd__clkbuf_2 hold3375 (.A(net5939),
    .X(net3902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3376 (.A(net5941),
    .X(net3903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3377 (.A(_00910_),
    .X(net3904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3378 (.A(\rbzero.spi_registers.spi_done ),
    .X(net3905));
 sky130_fd_sc_hd__buf_1 hold3379 (.A(net1776),
    .X(net3906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(net8001),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3380 (.A(_03343_),
    .X(net3907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3381 (.A(_00903_),
    .X(net3908));
 sky130_fd_sc_hd__clkbuf_2 hold3382 (.A(net5876),
    .X(net3909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3383 (.A(_02974_),
    .X(net3910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3384 (.A(_02975_),
    .X(net3911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3385 (.A(_00641_),
    .X(net3912));
 sky130_fd_sc_hd__buf_1 hold3386 (.A(net8006),
    .X(net3913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3388 (.A(_02834_),
    .X(net3915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3389 (.A(net4766),
    .X(net3916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net5251),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3390 (.A(net5945),
    .X(net3917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3391 (.A(_05064_),
    .X(net3918));
 sky130_fd_sc_hd__buf_1 hold3392 (.A(_05065_),
    .X(net3919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3393 (.A(_00475_),
    .X(net3920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3394 (.A(net7647),
    .X(net3921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3395 (.A(_03500_),
    .X(net3922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3396 (.A(net7650),
    .X(net3923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3397 (.A(_01019_),
    .X(net3924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3398 (.A(net7997),
    .X(net3925));
 sky130_fd_sc_hd__clkbuf_2 hold3399 (.A(net3476),
    .X(net3926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net5253),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3400 (.A(\rbzero.debug_overlay.facingY[0] ),
    .X(net3927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3401 (.A(_03746_),
    .X(net3928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3402 (.A(_03747_),
    .X(net3929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3403 (.A(_01217_),
    .X(net3930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3404 (.A(net4874),
    .X(net3931));
 sky130_fd_sc_hd__clkbuf_2 hold3405 (.A(net3729),
    .X(net3932));
 sky130_fd_sc_hd__buf_1 hold3406 (.A(net8357),
    .X(net3933));
 sky130_fd_sc_hd__buf_1 hold3407 (.A(net7815),
    .X(net3934));
 sky130_fd_sc_hd__clkbuf_2 hold3408 (.A(net7694),
    .X(net3935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3409 (.A(_02981_),
    .X(net3936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(net5331),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3410 (.A(_02982_),
    .X(net3937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3411 (.A(_00643_),
    .X(net3938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3412 (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .X(net3939));
 sky130_fd_sc_hd__clkbuf_2 hold3413 (.A(net3851),
    .X(net3940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3414 (.A(_03107_),
    .X(net3941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3415 (.A(_00747_),
    .X(net3942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3416 (.A(net8274),
    .X(net3943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3417 (.A(net4872),
    .X(net3944));
 sky130_fd_sc_hd__clkbuf_2 hold3418 (.A(net3559),
    .X(net3945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(net5333),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3420 (.A(_02652_),
    .X(net3947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3421 (.A(net4822),
    .X(net3948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3422 (.A(\rbzero.pov.spi_done ),
    .X(net3949));
 sky130_fd_sc_hd__clkbuf_2 hold3423 (.A(net2872),
    .X(net3950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3424 (.A(_03781_),
    .X(net3951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3425 (.A(_03782_),
    .X(net3952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3426 (.A(_01241_),
    .X(net3953));
 sky130_fd_sc_hd__clkbuf_2 hold3427 (.A(net7677),
    .X(net3954));
 sky130_fd_sc_hd__clkbuf_2 hold3428 (.A(_04597_),
    .X(net3955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3429 (.A(_09724_),
    .X(net3956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(net5231),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3430 (.A(_09726_),
    .X(net3957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3431 (.A(_00474_),
    .X(net3958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3432 (.A(net7686),
    .X(net3959));
 sky130_fd_sc_hd__clkbuf_2 hold3433 (.A(_06081_),
    .X(net3960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3434 (.A(_02731_),
    .X(net3961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3435 (.A(net7688),
    .X(net3962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3436 (.A(_00618_),
    .X(net3963));
 sky130_fd_sc_hd__buf_1 hold3437 (.A(\rbzero.map_rom.f2 ),
    .X(net3964));
 sky130_fd_sc_hd__clkbuf_4 hold3438 (.A(_06107_),
    .X(net3965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3439 (.A(net5919),
    .X(net3966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(net5233),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_1 hold3440 (.A(_04492_),
    .X(net3967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3441 (.A(net5780),
    .X(net3968));
 sky130_fd_sc_hd__buf_1 hold3442 (.A(net6000),
    .X(net3969));
 sky130_fd_sc_hd__buf_1 hold3443 (.A(_03117_),
    .X(net3970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3444 (.A(net7682),
    .X(net3971));
 sky130_fd_sc_hd__clkbuf_1 hold3445 (.A(_04472_),
    .X(net3972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3446 (.A(net8053),
    .X(net3973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3447 (.A(\rbzero.trace_state[2] ),
    .X(net3974));
 sky130_fd_sc_hd__buf_1 hold3448 (.A(net3451),
    .X(net3975));
 sky130_fd_sc_hd__buf_2 hold3449 (.A(_04474_),
    .X(net3976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(net5399),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3450 (.A(_01624_),
    .X(net3977));
 sky130_fd_sc_hd__clkbuf_2 hold3451 (.A(net7745),
    .X(net3978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3452 (.A(_03395_),
    .X(net3979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3453 (.A(_03396_),
    .X(net3980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3454 (.A(_00942_),
    .X(net3981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3455 (.A(net5504),
    .X(net3982));
 sky130_fd_sc_hd__buf_1 hold3456 (.A(_04737_),
    .X(net3983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3457 (.A(_06103_),
    .X(net3984));
 sky130_fd_sc_hd__buf_1 hold3458 (.A(_06114_),
    .X(net3985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3459 (.A(_08101_),
    .X(net3986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net5401),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3460 (.A(_08105_),
    .X(net3987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3461 (.A(_08106_),
    .X(net3988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3462 (.A(_00463_),
    .X(net3989));
 sky130_fd_sc_hd__buf_2 hold3463 (.A(\rbzero.debug_overlay.playerX[1] ),
    .X(net3990));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3464 (.A(_04678_),
    .X(net3991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3465 (.A(_03640_),
    .X(net3992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3466 (.A(net5909),
    .X(net3993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3467 (.A(_01177_),
    .X(net3994));
 sky130_fd_sc_hd__buf_1 hold3468 (.A(net6043),
    .X(net3995));
 sky130_fd_sc_hd__clkbuf_4 hold3469 (.A(_05731_),
    .X(net3996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(net5315),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3470 (.A(net6045),
    .X(net3997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3471 (.A(\rbzero.map_rom.f1 ),
    .X(net3998));
 sky130_fd_sc_hd__clkbuf_4 hold3472 (.A(_06109_),
    .X(net3999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3473 (.A(net7703),
    .X(net4000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3474 (.A(_00621_),
    .X(net4001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3475 (.A(\rbzero.debug_overlay.facingY[10] ),
    .X(net4002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3476 (.A(_03748_),
    .X(net4003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3477 (.A(_03749_),
    .X(net4004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3478 (.A(_01218_),
    .X(net4005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3479 (.A(net4047),
    .X(net4006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(net5317),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_2 hold3480 (.A(_06064_),
    .X(net4007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3481 (.A(_06131_),
    .X(net4008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3482 (.A(_06132_),
    .X(net4009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3483 (.A(_08107_),
    .X(net4010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3484 (.A(_08108_),
    .X(net4011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3485 (.A(_08109_),
    .X(net4012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3486 (.A(_08110_),
    .X(net4013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3487 (.A(_00464_),
    .X(net4014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3488 (.A(net4037),
    .X(net4015));
 sky130_fd_sc_hd__clkbuf_4 hold3489 (.A(net4039),
    .X(net4016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(net7564),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3490 (.A(_03083_),
    .X(net4017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3491 (.A(_00725_),
    .X(net4018));
 sky130_fd_sc_hd__buf_2 hold3492 (.A(\rbzero.debug_overlay.playerX[5] ),
    .X(net4019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3493 (.A(net7692),
    .X(net4020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3494 (.A(_03658_),
    .X(net4021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3495 (.A(_01181_),
    .X(net4022));
 sky130_fd_sc_hd__buf_1 hold3496 (.A(net5980),
    .X(net4023));
 sky130_fd_sc_hd__buf_4 hold3497 (.A(net5982),
    .X(net4024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3498 (.A(_03786_),
    .X(net4025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3499 (.A(_01245_),
    .X(net4026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(net4418),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3500 (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .X(net4027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3501 (.A(net1395),
    .X(net4028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3502 (.A(_02479_),
    .X(net4029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3503 (.A(net1396),
    .X(net4030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3504 (.A(_03081_),
    .X(net4031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3505 (.A(_00723_),
    .X(net4032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3506 (.A(net7711),
    .X(net4033));
 sky130_fd_sc_hd__clkbuf_4 hold3507 (.A(_06071_),
    .X(net4034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3508 (.A(_02736_),
    .X(net4035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3509 (.A(_00619_),
    .X(net4036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(net5283),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3510 (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .X(net4037));
 sky130_fd_sc_hd__buf_1 hold3511 (.A(net4015),
    .X(net4038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3512 (.A(_02485_),
    .X(net4039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3513 (.A(net4016),
    .X(net4040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3514 (.A(_03084_),
    .X(net4041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3515 (.A(_00726_),
    .X(net4042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3516 (.A(net8272),
    .X(net4043));
 sky130_fd_sc_hd__clkbuf_4 hold3517 (.A(_06035_),
    .X(net4044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3518 (.A(net7637),
    .X(net4045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3519 (.A(_00615_),
    .X(net4046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(net5285),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3520 (.A(\rbzero.map_rom.i_col[4] ),
    .X(net4047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3521 (.A(net4006),
    .X(net4048));
 sky130_fd_sc_hd__buf_2 hold3522 (.A(_06060_),
    .X(net4049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3523 (.A(_02746_),
    .X(net4050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3524 (.A(_00622_),
    .X(net4051));
 sky130_fd_sc_hd__clkbuf_2 hold3525 (.A(net4747),
    .X(net4052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3526 (.A(_06067_),
    .X(net4053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3527 (.A(_02713_),
    .X(net4054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3528 (.A(net5938),
    .X(net4055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3529 (.A(_00613_),
    .X(net4056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(net5196),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_4 hold3530 (.A(net7561),
    .X(net4057));
 sky130_fd_sc_hd__clkbuf_2 hold3531 (.A(_05059_),
    .X(net4058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3532 (.A(_09728_),
    .X(net4059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3533 (.A(_00476_),
    .X(net4060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3534 (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .X(net4061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3535 (.A(net3032),
    .X(net4062));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3536 (.A(_02969_),
    .X(net4063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3537 (.A(_03076_),
    .X(net4064));
 sky130_fd_sc_hd__buf_1 hold3538 (.A(net5964),
    .X(net4065));
 sky130_fd_sc_hd__buf_4 hold3539 (.A(_05051_),
    .X(net4066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(net5198),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3540 (.A(_05056_),
    .X(net4067));
 sky130_fd_sc_hd__buf_4 hold3541 (.A(_05295_),
    .X(net4068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3542 (.A(_00458_),
    .X(net4069));
 sky130_fd_sc_hd__clkbuf_1 hold3543 (.A(net4137),
    .X(net4070));
 sky130_fd_sc_hd__clkbuf_4 hold3544 (.A(_05674_),
    .X(net4071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3545 (.A(_01250_),
    .X(net4072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3546 (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .X(net4073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3547 (.A(net1425),
    .X(net4074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3548 (.A(_02483_),
    .X(net4075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3549 (.A(net1426),
    .X(net4076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net5188),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3550 (.A(_03082_),
    .X(net4077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3551 (.A(_00724_),
    .X(net4078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3552 (.A(net5967),
    .X(net4079));
 sky130_fd_sc_hd__buf_4 hold3553 (.A(net5969),
    .X(net4080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3554 (.A(_00482_),
    .X(net4081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3555 (.A(net7749),
    .X(net4082));
 sky130_fd_sc_hd__buf_2 hold3556 (.A(net3773),
    .X(net4083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3557 (.A(_03987_),
    .X(net4084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3558 (.A(_03990_),
    .X(net4085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3559 (.A(_03991_),
    .X(net4086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(net5190),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3560 (.A(_01622_),
    .X(net4087));
 sky130_fd_sc_hd__clkbuf_1 hold3561 (.A(net4144),
    .X(net4088));
 sky130_fd_sc_hd__buf_4 hold3562 (.A(_04025_),
    .X(net4089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3563 (.A(net5950),
    .X(net4090));
 sky130_fd_sc_hd__buf_2 hold3564 (.A(net7715),
    .X(net4091));
 sky130_fd_sc_hd__clkbuf_4 hold3565 (.A(_05675_),
    .X(net4092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3566 (.A(net7717),
    .X(net4093));
 sky130_fd_sc_hd__clkbuf_1 hold3567 (.A(net4159),
    .X(net4094));
 sky130_fd_sc_hd__clkbuf_4 hold3568 (.A(_04672_),
    .X(net4095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3569 (.A(_03118_),
    .X(net4096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(net5375),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_2 hold3570 (.A(_03119_),
    .X(net4097));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3571 (.A(_03803_),
    .X(net4098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3572 (.A(_03808_),
    .X(net4099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3573 (.A(_01252_),
    .X(net4100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3574 (.A(net5999),
    .X(net4101));
 sky130_fd_sc_hd__clkbuf_4 hold3575 (.A(net3969),
    .X(net4102));
 sky130_fd_sc_hd__clkbuf_4 hold3576 (.A(_05677_),
    .X(net4103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3577 (.A(_01244_),
    .X(net4104));
 sky130_fd_sc_hd__buf_2 hold3578 (.A(net5910),
    .X(net4105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3579 (.A(_04683_),
    .X(net4106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(net5377),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3580 (.A(_05068_),
    .X(net4107));
 sky130_fd_sc_hd__clkbuf_2 hold3581 (.A(_05082_),
    .X(net4108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3582 (.A(_00477_),
    .X(net4109));
 sky130_fd_sc_hd__clkbuf_2 hold3583 (.A(net7680),
    .X(net4110));
 sky130_fd_sc_hd__clkbuf_4 hold3584 (.A(_05672_),
    .X(net4111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3585 (.A(_03799_),
    .X(net4112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3586 (.A(_03800_),
    .X(net4113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3587 (.A(_01246_),
    .X(net4114));
 sky130_fd_sc_hd__clkbuf_2 hold3588 (.A(net7709),
    .X(net4115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3589 (.A(_05061_),
    .X(net4116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(net6064),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3590 (.A(_05062_),
    .X(net4117));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3591 (.A(net7563),
    .X(net4118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3592 (.A(_00479_),
    .X(net4119));
 sky130_fd_sc_hd__clkbuf_1 hold3593 (.A(net4131),
    .X(net4120));
 sky130_fd_sc_hd__clkbuf_2 hold3594 (.A(net4146),
    .X(net4121));
 sky130_fd_sc_hd__clkbuf_4 hold3595 (.A(_09718_),
    .X(net4122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3596 (.A(_09719_),
    .X(net4123));
 sky130_fd_sc_hd__buf_2 hold3597 (.A(_09720_),
    .X(net4124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3598 (.A(_00472_),
    .X(net4125));
 sky130_fd_sc_hd__clkbuf_4 hold3599 (.A(net7618),
    .X(net4126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(net6066),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_4 hold3600 (.A(_04712_),
    .X(net4127));
 sky130_fd_sc_hd__clkbuf_4 hold3601 (.A(_05680_),
    .X(net4128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3602 (.A(_03802_),
    .X(net4129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3603 (.A(_01248_),
    .X(net4130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3604 (.A(\gpout0.hpos[8] ),
    .X(net4131));
 sky130_fd_sc_hd__buf_4 hold3605 (.A(net4120),
    .X(net4132));
 sky130_fd_sc_hd__clkbuf_4 hold3606 (.A(_04024_),
    .X(net4133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3607 (.A(_09730_),
    .X(net4134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3608 (.A(_09731_),
    .X(net4135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3609 (.A(_00480_),
    .X(net4136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_00961_),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3610 (.A(net7738),
    .X(net4137));
 sky130_fd_sc_hd__clkbuf_4 hold3611 (.A(net4070),
    .X(net4138));
 sky130_fd_sc_hd__clkbuf_2 hold3612 (.A(_04669_),
    .X(net4139));
 sky130_fd_sc_hd__buf_1 hold3613 (.A(_05174_),
    .X(net4140));
 sky130_fd_sc_hd__clkbuf_4 hold3614 (.A(_05462_),
    .X(net4141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3615 (.A(_08096_),
    .X(net4142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3616 (.A(_00460_),
    .X(net4143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3617 (.A(\gpout0.hpos[9] ),
    .X(net4144));
 sky130_fd_sc_hd__clkbuf_4 hold3618 (.A(net4088),
    .X(net4145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3619 (.A(_05049_),
    .X(net4146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(net7523),
    .X(net889));
 sky130_fd_sc_hd__buf_4 hold3620 (.A(net4121),
    .X(net4147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3621 (.A(_05052_),
    .X(net4148));
 sky130_fd_sc_hd__clkbuf_4 hold3622 (.A(_05379_),
    .X(net4149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3623 (.A(_08095_),
    .X(net4150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3624 (.A(_00459_),
    .X(net4151));
 sky130_fd_sc_hd__buf_1 hold3625 (.A(net5754),
    .X(net4152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3626 (.A(_04717_),
    .X(net4153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3627 (.A(_04726_),
    .X(net4154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3628 (.A(_04752_),
    .X(net4155));
 sky130_fd_sc_hd__clkbuf_4 hold3629 (.A(_05053_),
    .X(net4156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_03131_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3630 (.A(_08094_),
    .X(net4157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3631 (.A(_00457_),
    .X(net4158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3632 (.A(\gpout0.vpos[3] ),
    .X(net4159));
 sky130_fd_sc_hd__clkbuf_4 hold3633 (.A(net4094),
    .X(net4160));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3634 (.A(_05042_),
    .X(net4161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3635 (.A(_05046_),
    .X(net4162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3636 (.A(_05047_),
    .X(net4163));
 sky130_fd_sc_hd__clkbuf_4 hold3637 (.A(_05546_),
    .X(net4164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3638 (.A(_08097_),
    .X(net4165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3639 (.A(_00461_),
    .X(net4166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(net4348),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3640 (.A(net8250),
    .X(net4167));
 sky130_fd_sc_hd__buf_4 hold3641 (.A(net3386),
    .X(net4168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3642 (.A(_05112_),
    .X(net4169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3643 (.A(_05119_),
    .X(net4170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3644 (.A(_05173_),
    .X(net4171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3645 (.A(_05175_),
    .X(net4172));
 sky130_fd_sc_hd__buf_2 hold3646 (.A(_05628_),
    .X(net4173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3647 (.A(_08098_),
    .X(net4174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3648 (.A(_00462_),
    .X(net4175));
 sky130_fd_sc_hd__buf_2 hold3649 (.A(\gpout0.vpos[5] ),
    .X(net4176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(net4847),
    .X(net892));
 sky130_fd_sc_hd__buf_2 hold3650 (.A(_04670_),
    .X(net4177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3651 (.A(_05043_),
    .X(net4178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3652 (.A(_03804_),
    .X(net4179));
 sky130_fd_sc_hd__buf_2 hold3653 (.A(\rbzero.side_hot ),
    .X(net4180));
 sky130_fd_sc_hd__buf_2 hold3654 (.A(_04510_),
    .X(net4181));
 sky130_fd_sc_hd__buf_1 hold3655 (.A(_04511_),
    .X(net4182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3656 (.A(_08111_),
    .X(net4183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3657 (.A(_00465_),
    .X(net4184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3658 (.A(\rbzero.vga_sync.vsync ),
    .X(net4185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3659 (.A(net3336),
    .X(net4186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(net4849),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3660 (.A(_04477_),
    .X(net4187));
 sky130_fd_sc_hd__clkbuf_2 hold3661 (.A(net4283),
    .X(net4188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3662 (.A(_09712_),
    .X(net4189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3663 (.A(_09713_),
    .X(net4190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3664 (.A(net7861),
    .X(net4191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3665 (.A(net7863),
    .X(net4192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3666 (.A(net8296),
    .X(net4193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3667 (.A(net8298),
    .X(net4194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3668 (.A(net8115),
    .X(net4195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3669 (.A(_00850_),
    .X(net4196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(net5407),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3670 (.A(net841),
    .X(net4197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3671 (.A(net8117),
    .X(net4198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3672 (.A(_00832_),
    .X(net4199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3673 (.A(net599),
    .X(net4200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3674 (.A(net7884),
    .X(net4201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3675 (.A(net7886),
    .X(net4202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3676 (.A(net7881),
    .X(net4203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3677 (.A(net7883),
    .X(net4204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3678 (.A(net7890),
    .X(net4205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3679 (.A(net7892),
    .X(net4206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(net5409),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3680 (.A(net8134),
    .X(net4207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3681 (.A(net8136),
    .X(net4208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3682 (.A(net988),
    .X(net4209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3683 (.A(net7887),
    .X(net4210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3684 (.A(net7889),
    .X(net4211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3685 (.A(net7896),
    .X(net4212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3686 (.A(net7898),
    .X(net4213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3687 (.A(net7893),
    .X(net4214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3688 (.A(net7895),
    .X(net4215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3689 (.A(net8301),
    .X(net4216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(net8122),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3690 (.A(net8303),
    .X(net4217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3691 (.A(net7899),
    .X(net4218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3692 (.A(net7901),
    .X(net4219));
 sky130_fd_sc_hd__buf_1 hold3693 (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(net4220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3694 (.A(net8000),
    .X(net4221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3695 (.A(net865),
    .X(net4222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3696 (.A(net7908),
    .X(net4223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3697 (.A(net7910),
    .X(net4224));
 sky130_fd_sc_hd__buf_1 hold3698 (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(net4225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3699 (.A(net8069),
    .X(net4226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(net4294),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3700 (.A(net972),
    .X(net4227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3701 (.A(net7854),
    .X(net4228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3702 (.A(net7856),
    .X(net4229));
 sky130_fd_sc_hd__buf_1 hold3703 (.A(net8144),
    .X(net4230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3704 (.A(_00900_),
    .X(net4231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3705 (.A(net1367),
    .X(net4232));
 sky130_fd_sc_hd__buf_1 hold3706 (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(net4233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3707 (.A(net8003),
    .X(net4234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3708 (.A(net1016),
    .X(net4235));
 sky130_fd_sc_hd__buf_2 hold3709 (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(net4236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(net5275),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3710 (.A(net8139),
    .X(net4237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3711 (.A(net1121),
    .X(net4238));
 sky130_fd_sc_hd__buf_1 hold3712 (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(net4239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3713 (.A(net8019),
    .X(net4240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3714 (.A(net835),
    .X(net4241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3716 (.A(net7912),
    .X(net4243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3717 (.A(net7914),
    .X(net4244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3718 (.A(net8306),
    .X(net4245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3719 (.A(net8308),
    .X(net4246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(net5277),
    .X(net899));
 sky130_fd_sc_hd__buf_1 hold3720 (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(net4247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3721 (.A(net8016),
    .X(net4248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3722 (.A(net970),
    .X(net4249));
 sky130_fd_sc_hd__buf_1 hold3723 (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(net4250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3724 (.A(net8080),
    .X(net4251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3725 (.A(net851),
    .X(net4252));
 sky130_fd_sc_hd__buf_1 hold3726 (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(net4253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3727 (.A(net8013),
    .X(net4254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3728 (.A(net1010),
    .X(net4255));
 sky130_fd_sc_hd__clkbuf_1 hold3729 (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(net4256));
 sky130_fd_sc_hd__buf_1 hold373 (.A(net5656),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3730 (.A(net8022),
    .X(net4257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3731 (.A(net823),
    .X(net4258));
 sky130_fd_sc_hd__clkbuf_2 hold3732 (.A(net8145),
    .X(net4259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3733 (.A(_00495_),
    .X(net4260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3734 (.A(net1155),
    .X(net4261));
 sky130_fd_sc_hd__buf_1 hold3735 (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(net4262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3736 (.A(net8010),
    .X(net4263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3737 (.A(net1039),
    .X(net4264));
 sky130_fd_sc_hd__buf_1 hold3738 (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(net4265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3739 (.A(_00519_),
    .X(net4266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(net5658),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3740 (.A(net1029),
    .X(net4267));
 sky130_fd_sc_hd__buf_2 hold3741 (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(net4268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3742 (.A(net8133),
    .X(net4269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3743 (.A(net1049),
    .X(net4270));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3744 (.A(net8146),
    .X(net4271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3745 (.A(_00497_),
    .X(net4272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3746 (.A(net1586),
    .X(net4273));
 sky130_fd_sc_hd__clkbuf_1 hold3747 (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(net4274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3748 (.A(net8030),
    .X(net4275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3749 (.A(net985),
    .X(net4276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(net5295),
    .X(net902));
 sky130_fd_sc_hd__buf_2 hold3750 (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(net4277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3751 (.A(net8127),
    .X(net4278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3752 (.A(net961),
    .X(net4279));
 sky130_fd_sc_hd__buf_2 hold3753 (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(net4280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3754 (.A(net8142),
    .X(net4281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3755 (.A(net1107),
    .X(net4282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3756 (.A(\rbzero.debug_overlay.playerY[-1] ),
    .X(net4283));
 sky130_fd_sc_hd__buf_1 hold3757 (.A(net4188),
    .X(net4284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3758 (.A(_01190_),
    .X(net4285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3759 (.A(net2398),
    .X(net4286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(net5297),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3761 (.A(net7933),
    .X(net4288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3762 (.A(net778),
    .X(net4289));
 sky130_fd_sc_hd__buf_1 hold3763 (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(net4290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3764 (.A(net8089),
    .X(net4291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3765 (.A(net992),
    .X(net4292));
 sky130_fd_sc_hd__clkbuf_4 hold3766 (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(net4293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3767 (.A(net8124),
    .X(net4294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3768 (.A(net897),
    .X(net4295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(net6095),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3770 (.A(net7921),
    .X(net4297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3771 (.A(net7923),
    .X(net4298));
 sky130_fd_sc_hd__buf_1 hold3772 (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(net4299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3773 (.A(net8121),
    .X(net4300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3774 (.A(net949),
    .X(net4301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3775 (.A(net8309),
    .X(net4302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3776 (.A(net8311),
    .X(net4303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3777 (.A(\rbzero.row_render.size[5] ),
    .X(net4304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3778 (.A(net3151),
    .X(net4305));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3779 (.A(net8156),
    .X(net4306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(net6097),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3780 (.A(_00764_),
    .X(net4307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3781 (.A(net1078),
    .X(net4308));
 sky130_fd_sc_hd__clkbuf_2 hold3782 (.A(net8160),
    .X(net4309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3783 (.A(_00757_),
    .X(net4310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3784 (.A(net3037),
    .X(net4311));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3785 (.A(net8159),
    .X(net4312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3786 (.A(_00897_),
    .X(net4313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3787 (.A(net1035),
    .X(net4314));
 sky130_fd_sc_hd__clkbuf_2 hold3788 (.A(net8158),
    .X(net4315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3789 (.A(_00758_),
    .X(net4316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_01051_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3790 (.A(net2711),
    .X(net4317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3792 (.A(net7925),
    .X(net4319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3793 (.A(net7927),
    .X(net4320));
 sky130_fd_sc_hd__clkbuf_2 hold3794 (.A(net8148),
    .X(net4321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3795 (.A(net8149),
    .X(net4322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3796 (.A(net673),
    .X(net4323));
 sky130_fd_sc_hd__clkbuf_2 hold3797 (.A(net8163),
    .X(net4324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3798 (.A(_00763_),
    .X(net4325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3799 (.A(net1063),
    .X(net4326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(net5164),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3800 (.A(\rbzero.pov.ready_buffer[50] ),
    .X(net4327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3801 (.A(_03676_),
    .X(net4328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3802 (.A(_01188_),
    .X(net4329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3803 (.A(net3434),
    .X(net4330));
 sky130_fd_sc_hd__buf_1 hold3804 (.A(net4250),
    .X(net4331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3805 (.A(_08065_),
    .X(net4332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3806 (.A(_00434_),
    .X(net4333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3807 (.A(net1793),
    .X(net4334));
 sky130_fd_sc_hd__clkbuf_2 hold3808 (.A(net8153),
    .X(net4335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3809 (.A(net8154),
    .X(net4336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(net5166),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3810 (.A(net745),
    .X(net4337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3811 (.A(net3715),
    .X(net4338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3812 (.A(net3405),
    .X(net4339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3813 (.A(net8312),
    .X(net4340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3814 (.A(net8314),
    .X(net4341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3815 (.A(net7905),
    .X(net4342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3816 (.A(net7907),
    .X(net4343));
 sky130_fd_sc_hd__clkbuf_2 hold3817 (.A(net8215),
    .X(net4344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3818 (.A(_01186_),
    .X(net4345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3819 (.A(net3416),
    .X(net4346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(net5307),
    .X(net909));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3820 (.A(net8170),
    .X(net4347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3821 (.A(_00759_),
    .X(net4348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3822 (.A(net891),
    .X(net4349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3823 (.A(net7876),
    .X(net4350));
 sky130_fd_sc_hd__buf_1 hold3824 (.A(net7878),
    .X(net4351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3825 (.A(net7937),
    .X(net4352));
 sky130_fd_sc_hd__buf_1 hold3826 (.A(net7939),
    .X(net4353));
 sky130_fd_sc_hd__clkbuf_2 hold3827 (.A(net8166),
    .X(net4354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3828 (.A(_00767_),
    .X(net4355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3829 (.A(net1291),
    .X(net4356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(net5309),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_2 hold3830 (.A(net8165),
    .X(net4357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3831 (.A(_00777_),
    .X(net4358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3832 (.A(net838),
    .X(net4359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3833 (.A(net3686),
    .X(net4360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3834 (.A(net3423),
    .X(net4361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3835 (.A(net5742),
    .X(net4362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3836 (.A(_03674_),
    .X(net4363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3837 (.A(_01187_),
    .X(net4364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3838 (.A(net3318),
    .X(net4365));
 sky130_fd_sc_hd__clkbuf_2 hold3839 (.A(net8167),
    .X(net4366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(net5291),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3840 (.A(_00774_),
    .X(net4367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3841 (.A(net959),
    .X(net4368));
 sky130_fd_sc_hd__clkbuf_2 hold3842 (.A(net8164),
    .X(net4369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3843 (.A(_00768_),
    .X(net4370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3844 (.A(net1178),
    .X(net4371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3845 (.A(net8373),
    .X(net4372));
 sky130_fd_sc_hd__buf_1 hold3846 (.A(net3430),
    .X(net4373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3847 (.A(net5736),
    .X(net4374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3848 (.A(_03697_),
    .X(net4375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3849 (.A(_01194_),
    .X(net4376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(net5293),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3850 (.A(net3474),
    .X(net4377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3851 (.A(net7851),
    .X(net4378));
 sky130_fd_sc_hd__buf_1 hold3852 (.A(net7853),
    .X(net4379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3853 (.A(net7869),
    .X(net4380));
 sky130_fd_sc_hd__buf_1 hold3854 (.A(net7871),
    .X(net4381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3855 (.A(net7866),
    .X(net4382));
 sky130_fd_sc_hd__buf_1 hold3856 (.A(net7868),
    .X(net4383));
 sky130_fd_sc_hd__clkbuf_2 hold3857 (.A(net8168),
    .X(net4384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3858 (.A(_00776_),
    .X(net4385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3859 (.A(net2068),
    .X(net4386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(net5335),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3860 (.A(net8320),
    .X(net4387));
 sky130_fd_sc_hd__buf_1 hold3861 (.A(net8322),
    .X(net4388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3862 (.A(net8056),
    .X(net4389));
 sky130_fd_sc_hd__buf_1 hold3863 (.A(net8058),
    .X(net4390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3864 (.A(net7940),
    .X(net4391));
 sky130_fd_sc_hd__buf_1 hold3865 (.A(net7942),
    .X(net4392));
 sky130_fd_sc_hd__clkbuf_2 hold3866 (.A(net8169),
    .X(net4393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3867 (.A(_00775_),
    .X(net4394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3868 (.A(net1832),
    .X(net4395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3869 (.A(net8381),
    .X(net4396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(net5337),
    .X(net914));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3870 (.A(net3467),
    .X(net4397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3871 (.A(net7915),
    .X(net4398));
 sky130_fd_sc_hd__buf_1 hold3872 (.A(net7917),
    .X(net4399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3873 (.A(net7830),
    .X(net4400));
 sky130_fd_sc_hd__buf_1 hold3874 (.A(net3484),
    .X(net4401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3875 (.A(net8323),
    .X(net4402));
 sky130_fd_sc_hd__buf_1 hold3876 (.A(net8325),
    .X(net4403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3877 (.A(net7902),
    .X(net4404));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3878 (.A(net7904),
    .X(net4405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3879 (.A(net8318),
    .X(net4406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(net5339),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3880 (.A(net3488),
    .X(net4407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3883 (.A(net7945),
    .X(net4410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3884 (.A(net1058),
    .X(net4411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3885 (.A(net7796),
    .X(net4412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3886 (.A(net7798),
    .X(net4413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3887 (.A(net8036),
    .X(net4414));
 sky130_fd_sc_hd__buf_1 hold3888 (.A(net8038),
    .X(net4415));
 sky130_fd_sc_hd__clkbuf_2 hold3889 (.A(\rbzero.debug_overlay.facingY[-1] ),
    .X(net4416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(net5341),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3890 (.A(_03745_),
    .X(net4417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3891 (.A(_01216_),
    .X(net4418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3892 (.A(net877),
    .X(net4419));
 sky130_fd_sc_hd__clkbuf_2 hold3893 (.A(net8173),
    .X(net4420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3894 (.A(_00769_),
    .X(net4421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3895 (.A(net1205),
    .X(net4422));
 sky130_fd_sc_hd__buf_2 hold3896 (.A(net8252),
    .X(net4423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3897 (.A(_02754_),
    .X(net4424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3898 (.A(net8098),
    .X(net4425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3899 (.A(net653),
    .X(net4426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(net4882),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3900 (.A(net7847),
    .X(net4427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3901 (.A(net3542),
    .X(net4428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3902 (.A(net7918),
    .X(net4429));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3903 (.A(net3531),
    .X(net4430));
 sky130_fd_sc_hd__clkbuf_2 hold3904 (.A(net8175),
    .X(net4431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3905 (.A(_00770_),
    .X(net4432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3906 (.A(net1240),
    .X(net4433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3907 (.A(net7788),
    .X(net4434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3908 (.A(net3532),
    .X(net4435));
 sky130_fd_sc_hd__clkbuf_4 hold3909 (.A(net8235),
    .X(net4436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(net4884),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3910 (.A(_01193_),
    .X(net4437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3911 (.A(net665),
    .X(net4438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3912 (.A(net8379),
    .X(net4439));
 sky130_fd_sc_hd__buf_1 hold3913 (.A(net3551),
    .X(net4440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3914 (.A(net5782),
    .X(net4441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3915 (.A(_03624_),
    .X(net4442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3916 (.A(_03625_),
    .X(net4443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3917 (.A(_01172_),
    .X(net4444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3918 (.A(net3340),
    .X(net4445));
 sky130_fd_sc_hd__buf_2 hold3919 (.A(\rbzero.debug_overlay.facingX[10] ),
    .X(net4446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(net6057),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3920 (.A(_03727_),
    .X(net4447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3921 (.A(_01207_),
    .X(net4448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3922 (.A(net776),
    .X(net4449));
 sky130_fd_sc_hd__clkbuf_4 hold3923 (.A(net7568),
    .X(net4450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3924 (.A(_03142_),
    .X(net4451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3925 (.A(_00766_),
    .X(net4452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3926 (.A(net637),
    .X(net4453));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3927 (.A(\rbzero.pov.ready_buffer[70] ),
    .X(net4454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3928 (.A(_03645_),
    .X(net4455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3929 (.A(_01178_),
    .X(net4456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(net6059),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3930 (.A(net3390),
    .X(net4457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3931 (.A(net7879),
    .X(net4458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3932 (.A(net3574),
    .X(net4459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3933 (.A(net8348),
    .X(net4460));
 sky130_fd_sc_hd__buf_1 hold3934 (.A(net3586),
    .X(net4461));
 sky130_fd_sc_hd__buf_1 hold3935 (.A(\rbzero.debug_overlay.facingX[-6] ),
    .X(net4462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3936 (.A(_03715_),
    .X(net4463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3937 (.A(_01200_),
    .X(net4464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3938 (.A(net1027),
    .X(net4465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_01599_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3940 (.A(net8177),
    .X(net4467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3941 (.A(_01213_),
    .X(net4468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3942 (.A(net1060),
    .X(net4469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3943 (.A(net8390),
    .X(net4470));
 sky130_fd_sc_hd__clkbuf_2 hold3944 (.A(net3573),
    .X(net4471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3946 (.A(net8179),
    .X(net4473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3947 (.A(_01199_),
    .X(net4474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3948 (.A(net1114),
    .X(net4475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(net5255),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3950 (.A(net8184),
    .X(net4477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3951 (.A(_01198_),
    .X(net4478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3952 (.A(net2243),
    .X(net4479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3953 (.A(net7826),
    .X(net4480));
 sky130_fd_sc_hd__buf_1 hold3954 (.A(net3599),
    .X(net4481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3955 (.A(net8328),
    .X(net4482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3956 (.A(net3600),
    .X(net4483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3957 (.A(net8326),
    .X(net4484));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3958 (.A(net3617),
    .X(net4485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(net5257),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3960 (.A(net8186),
    .X(net4487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3961 (.A(_01214_),
    .X(net4488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3962 (.A(net1056),
    .X(net4489));
 sky130_fd_sc_hd__buf_1 hold3963 (.A(\rbzero.pov.ready_buffer[66] ),
    .X(net4490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3964 (.A(_03629_),
    .X(net4491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3965 (.A(_03630_),
    .X(net4492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3966 (.A(_01174_),
    .X(net4493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3967 (.A(net3462),
    .X(net4494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3968 (.A(net8394),
    .X(net4495));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3969 (.A(net3630),
    .X(net4496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(net6106),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3970 (.A(net8330),
    .X(net4497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3971 (.A(net1791),
    .X(net4498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3972 (.A(net7947),
    .X(net4499));
 sky130_fd_sc_hd__clkbuf_2 hold3973 (.A(net3655),
    .X(net4500));
 sky130_fd_sc_hd__clkbuf_4 hold3974 (.A(net8268),
    .X(net4501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3975 (.A(_03754_),
    .X(net4502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3976 (.A(_01222_),
    .X(net4503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3977 (.A(net629),
    .X(net4504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3978 (.A(net7930),
    .X(net4505));
 sky130_fd_sc_hd__clkbuf_2 hold3979 (.A(net3718),
    .X(net4506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(net6108),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3980 (.A(net7981),
    .X(net4507));
 sky130_fd_sc_hd__clkbuf_2 hold3981 (.A(net3833),
    .X(net4508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3982 (.A(_00419_),
    .X(net4509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3983 (.A(net3410),
    .X(net4510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3984 (.A(\rbzero.row_render.size[6] ),
    .X(net4511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3985 (.A(net3014),
    .X(net4512));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3986 (.A(\rbzero.debug_overlay.facingX[0] ),
    .X(net4513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3987 (.A(_03726_),
    .X(net4514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3988 (.A(_01206_),
    .X(net4515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3989 (.A(net780),
    .X(net4516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_01363_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3990 (.A(net7935),
    .X(net4517));
 sky130_fd_sc_hd__clkbuf_2 hold3991 (.A(net3378),
    .X(net4518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3992 (.A(net7808),
    .X(net4519));
 sky130_fd_sc_hd__clkbuf_2 hold3993 (.A(net3727),
    .X(net4520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3994 (.A(net7874),
    .X(net4521));
 sky130_fd_sc_hd__buf_1 hold3995 (.A(net3726),
    .X(net4522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3996 (.A(net8334),
    .X(net4523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3997 (.A(net3724),
    .X(net4524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3998 (.A(net7953),
    .X(net4525));
 sky130_fd_sc_hd__clkbuf_2 hold3999 (.A(net1663),
    .X(net4526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(net5219),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4000 (.A(net7699),
    .X(net4527));
 sky130_fd_sc_hd__buf_4 hold4001 (.A(net3538),
    .X(net4528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4002 (.A(_02760_),
    .X(net4529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4003 (.A(_02761_),
    .X(net4530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4004 (.A(_02766_),
    .X(net4531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4005 (.A(net8130),
    .X(net4532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4006 (.A(net1003),
    .X(net4533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4007 (.A(net7857),
    .X(net4534));
 sky130_fd_sc_hd__clkbuf_2 hold4008 (.A(net3725),
    .X(net4535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4009 (.A(net8332),
    .X(net4536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(net5221),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_2 hold4010 (.A(net3723),
    .X(net4537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4011 (.A(net8081),
    .X(net4538));
 sky130_fd_sc_hd__clkbuf_2 hold4012 (.A(net3728),
    .X(net4539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4013 (.A(net7949),
    .X(net4540));
 sky130_fd_sc_hd__clkbuf_2 hold4014 (.A(net3764),
    .X(net4541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4016 (.A(net8190),
    .X(net4543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4017 (.A(_00413_),
    .X(net4544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4018 (.A(net3383),
    .X(net4545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4019 (.A(net7987),
    .X(net4546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(net5363),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_2 hold4020 (.A(net3854),
    .X(net4547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4021 (.A(_00418_),
    .X(net4548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4022 (.A(net3385),
    .X(net4549));
 sky130_fd_sc_hd__clkbuf_2 hold4023 (.A(net4239),
    .X(net4550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4024 (.A(_08051_),
    .X(net4551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4025 (.A(_00422_),
    .X(net4552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4026 (.A(net3393),
    .X(net4553));
 sky130_fd_sc_hd__buf_2 hold4027 (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(net4554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4028 (.A(_03762_),
    .X(net4555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4029 (.A(_01227_),
    .X(net4556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(net5365),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4030 (.A(net811),
    .X(net4557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4031 (.A(net8340),
    .X(net4558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4032 (.A(net672),
    .X(net4559));
 sky130_fd_sc_hd__buf_2 hold4033 (.A(net8245),
    .X(net4560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4034 (.A(_03778_),
    .X(net4561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4035 (.A(_01238_),
    .X(net4562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4036 (.A(net646),
    .X(net4563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4037 (.A(net7951),
    .X(net4564));
 sky130_fd_sc_hd__clkbuf_2 hold4038 (.A(net2877),
    .X(net4565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4039 (.A(net7955),
    .X(net4566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(net5311),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_2 hold4040 (.A(net3755),
    .X(net4567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4041 (.A(net7957),
    .X(net4568));
 sky130_fd_sc_hd__clkbuf_2 hold4042 (.A(net3801),
    .X(net4569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4044 (.A(_08044_),
    .X(net4571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4045 (.A(_00417_),
    .X(net4572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4046 (.A(net2878),
    .X(net4573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4047 (.A(net7959),
    .X(net4574));
 sky130_fd_sc_hd__clkbuf_2 hold4048 (.A(net3791),
    .X(net4575));
 sky130_fd_sc_hd__clkbuf_2 hold4049 (.A(net4256),
    .X(net4576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(net5313),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4050 (.A(_08053_),
    .X(net4577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4051 (.A(_00423_),
    .X(net4578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4052 (.A(net3206),
    .X(net4579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4053 (.A(net7995),
    .X(net4580));
 sky130_fd_sc_hd__clkbuf_2 hold4054 (.A(net3796),
    .X(net4581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4055 (.A(net8415),
    .X(net4582));
 sky130_fd_sc_hd__clkbuf_2 hold4056 (.A(net3788),
    .X(net4583));
 sky130_fd_sc_hd__clkbuf_2 hold4057 (.A(net4274),
    .X(net4584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4058 (.A(_08054_),
    .X(net4585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4059 (.A(_00424_),
    .X(net4586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(net6087),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4060 (.A(net1664),
    .X(net4587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4061 (.A(net7961),
    .X(net4588));
 sky130_fd_sc_hd__clkbuf_2 hold4062 (.A(net3806),
    .X(net4589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4063 (.A(\rbzero.pov.ready_buffer[0] ),
    .X(net4590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4064 (.A(net1171),
    .X(net4591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4065 (.A(_01230_),
    .X(net4592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4066 (.A(net1172),
    .X(net4593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4068 (.A(net8212),
    .X(net4595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4069 (.A(_01204_),
    .X(net4596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(net6089),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4070 (.A(net817),
    .X(net4597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4071 (.A(net8248),
    .X(net4598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4072 (.A(_02755_),
    .X(net4599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4073 (.A(_04011_),
    .X(net4600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4074 (.A(net8101),
    .X(net4601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4075 (.A(net682),
    .X(net4602));
 sky130_fd_sc_hd__buf_2 hold4076 (.A(net8259),
    .X(net4603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4077 (.A(_03763_),
    .X(net4604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4078 (.A(_01228_),
    .X(net4605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4079 (.A(net792),
    .X(net4606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_01553_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4080 (.A(net8342),
    .X(net4607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4081 (.A(net3587),
    .X(net4608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4082 (.A(net7963),
    .X(net4609));
 sky130_fd_sc_hd__clkbuf_2 hold4083 (.A(net3831),
    .X(net4610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4084 (.A(net8457),
    .X(net4611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4085 (.A(net1154),
    .X(net4612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4086 (.A(_09216_),
    .X(net4613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4087 (.A(\rbzero.row_render.size[7] ),
    .X(net4614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4088 (.A(net3365),
    .X(net4615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4089 (.A(net5703),
    .X(net4616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net5235),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4090 (.A(_03665_),
    .X(net4617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4091 (.A(_03666_),
    .X(net4618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4092 (.A(_01183_),
    .X(net4619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4093 (.A(net3490),
    .X(net4620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4094 (.A(net8336),
    .X(net4621));
 sky130_fd_sc_hd__clkbuf_2 hold4095 (.A(net3830),
    .X(net4622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4096 (.A(net8338),
    .X(net4623));
 sky130_fd_sc_hd__clkbuf_2 hold4097 (.A(net3832),
    .X(net4624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4099 (.A(_03712_),
    .X(net4626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(net5237),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4100 (.A(net8172),
    .X(net4627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4101 (.A(net3408),
    .X(net4628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4102 (.A(net8350),
    .X(net4629));
 sky130_fd_sc_hd__clkbuf_2 hold4103 (.A(net3889),
    .X(net4630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4104 (.A(_09825_),
    .X(net4631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4105 (.A(_09832_),
    .X(net4632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4106 (.A(_09840_),
    .X(net4633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4107 (.A(_09844_),
    .X(net4634));
 sky130_fd_sc_hd__clkbuf_4 hold4108 (.A(net8262),
    .X(net4635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4109 (.A(_03768_),
    .X(net4636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(net6102),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4110 (.A(_01232_),
    .X(net4637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4111 (.A(net684),
    .X(net4638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4112 (.A(net8346),
    .X(net4639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4113 (.A(net744),
    .X(net4640));
 sky130_fd_sc_hd__buf_1 hold4114 (.A(net5936),
    .X(net4641));
 sky130_fd_sc_hd__clkbuf_2 hold4115 (.A(_06037_),
    .X(net4642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4116 (.A(_06096_),
    .X(net4643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4117 (.A(_06102_),
    .X(net4644));
 sky130_fd_sc_hd__buf_1 hold4118 (.A(_06115_),
    .X(net4645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4119 (.A(_06116_),
    .X(net4646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(net6104),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4120 (.A(_06161_),
    .X(net4647));
 sky130_fd_sc_hd__buf_4 hold4121 (.A(_09767_),
    .X(net4648));
 sky130_fd_sc_hd__buf_4 hold4122 (.A(_09822_),
    .X(net4649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4123 (.A(net7969),
    .X(net4650));
 sky130_fd_sc_hd__clkbuf_2 hold4124 (.A(net3836),
    .X(net4651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4125 (.A(net8404),
    .X(net4652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4126 (.A(net3841),
    .X(net4653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4127 (.A(net7973),
    .X(net4654));
 sky130_fd_sc_hd__clkbuf_2 hold4128 (.A(net3855),
    .X(net4655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4129 (.A(net7975),
    .X(net4656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(_01071_),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_2 hold4130 (.A(net3856),
    .X(net4657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4131 (.A(net7979),
    .X(net4658));
 sky130_fd_sc_hd__clkbuf_2 hold4132 (.A(net3861),
    .X(net4659));
 sky130_fd_sc_hd__buf_1 hold4133 (.A(net4265),
    .X(net4660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4134 (.A(_08063_),
    .X(net4661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4135 (.A(_00433_),
    .X(net4662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4136 (.A(net3477),
    .X(net4663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4137 (.A(net7985),
    .X(net4664));
 sky130_fd_sc_hd__clkbuf_2 hold4138 (.A(net3392),
    .X(net4665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4139 (.A(net8344),
    .X(net4666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(net7882),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_2 hold4140 (.A(net3382),
    .X(net4667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4141 (.A(net7977),
    .X(net4668));
 sky130_fd_sc_hd__clkbuf_2 hold4142 (.A(net3869),
    .X(net4669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4144 (.A(net8188),
    .X(net4671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4145 (.A(_00415_),
    .X(net4672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4146 (.A(net3560),
    .X(net4673));
 sky130_fd_sc_hd__buf_4 hold4147 (.A(net4290),
    .X(net4674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4148 (.A(_08062_),
    .X(net4675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4149 (.A(_00432_),
    .X(net4676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(net4878),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4150 (.A(net3381),
    .X(net4677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4152 (.A(net8202),
    .X(net4679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4153 (.A(_00414_),
    .X(net4680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4154 (.A(net3379),
    .X(net4681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4156 (.A(_08048_),
    .X(net4683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4157 (.A(_00420_),
    .X(net4684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4158 (.A(net3013),
    .X(net4685));
 sky130_fd_sc_hd__clkbuf_4 hold4159 (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(net4686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(net4880),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4160 (.A(_03775_),
    .X(net4687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4161 (.A(_01236_),
    .X(net4688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4162 (.A(net747),
    .X(net4689));
 sky130_fd_sc_hd__clkbuf_2 hold4163 (.A(net4220),
    .X(net4690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4164 (.A(_08056_),
    .X(net4691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4165 (.A(_00426_),
    .X(net4692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4166 (.A(net3425),
    .X(net4693));
 sky130_fd_sc_hd__clkbuf_2 hold4167 (.A(net4299),
    .X(net4694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4168 (.A(_08055_),
    .X(net4695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4169 (.A(_00425_),
    .X(net4696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(net5319),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4170 (.A(net2197),
    .X(net4697));
 sky130_fd_sc_hd__buf_2 hold4171 (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(net4698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4172 (.A(_03759_),
    .X(net4699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4173 (.A(_01225_),
    .X(net4700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4174 (.A(net763),
    .X(net4701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4176 (.A(net7805),
    .X(net4703));
 sky130_fd_sc_hd__clkbuf_2 hold4177 (.A(_07868_),
    .X(net4704));
 sky130_fd_sc_hd__buf_4 hold4178 (.A(net4225),
    .X(net4705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4179 (.A(_08061_),
    .X(net4706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(net5321),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4180 (.A(_00431_),
    .X(net4707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4181 (.A(net3422),
    .X(net4708));
 sky130_fd_sc_hd__buf_2 hold4182 (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(net4709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4183 (.A(_03779_),
    .X(net4710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4184 (.A(_01239_),
    .X(net4711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4185 (.A(net677),
    .X(net4712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4186 (.A(net8244),
    .X(net4713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4187 (.A(_02513_),
    .X(net4714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4188 (.A(_04005_),
    .X(net4715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4189 (.A(net8106),
    .X(net4716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(net5367),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4190 (.A(net694),
    .X(net4717));
 sky130_fd_sc_hd__clkbuf_2 hold4191 (.A(net4233),
    .X(net4718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4192 (.A(_08060_),
    .X(net4719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4193 (.A(_00430_),
    .X(net4720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4194 (.A(net627),
    .X(net4721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4195 (.A(net8005),
    .X(net4722));
 sky130_fd_sc_hd__clkbuf_2 hold4196 (.A(net3913),
    .X(net4723));
 sky130_fd_sc_hd__clkbuf_2 hold4197 (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(net4724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4198 (.A(_02581_),
    .X(net4725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4199 (.A(_02584_),
    .X(net4726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(net5369),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4200 (.A(net8077),
    .X(net4727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4201 (.A(net3640),
    .X(net4728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4203 (.A(_08049_),
    .X(net4730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4204 (.A(_00421_),
    .X(net4731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4205 (.A(net3429),
    .X(net4732));
 sky130_fd_sc_hd__buf_2 hold4206 (.A(net8253),
    .X(net4733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4207 (.A(_03753_),
    .X(net4734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4208 (.A(_01221_),
    .X(net4735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4209 (.A(net639),
    .X(net4736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net8119),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_2 hold4210 (.A(net4253),
    .X(net4737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4211 (.A(_08057_),
    .X(net4738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4212 (.A(_00427_),
    .X(net4739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4213 (.A(net3296),
    .X(net4740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4214 (.A(net8356),
    .X(net4741));
 sky130_fd_sc_hd__clkbuf_2 hold4215 (.A(net3933),
    .X(net4742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4217 (.A(net8205),
    .X(net4744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4218 (.A(_00416_),
    .X(net4745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4219 (.A(net3355),
    .X(net4746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(net4300),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4220 (.A(\rbzero.debug_overlay.playerY[1] ),
    .X(net4747));
 sky130_fd_sc_hd__clkbuf_4 hold4221 (.A(net4052),
    .X(net4748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4222 (.A(_01192_),
    .X(net4749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4223 (.A(net618),
    .X(net4750));
 sky130_fd_sc_hd__clkbuf_2 hold4224 (.A(net4247),
    .X(net4751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4225 (.A(_08059_),
    .X(net4752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4226 (.A(_00429_),
    .X(net4753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4227 (.A(net3360),
    .X(net4754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4228 (.A(net7814),
    .X(net4755));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4229 (.A(net3934),
    .X(net4756));
 sky130_fd_sc_hd__buf_1 hold423 (.A(net7885),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_2 hold4230 (.A(net4262),
    .X(net4757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4231 (.A(net8266),
    .X(net4758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4232 (.A(_00428_),
    .X(net4759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4233 (.A(net1681),
    .X(net4760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4234 (.A(net8273),
    .X(net4761));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4235 (.A(net3943),
    .X(net4762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4237 (.A(_02820_),
    .X(net4764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4238 (.A(_02823_),
    .X(net4765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4239 (.A(net8095),
    .X(net4766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(net5391),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4240 (.A(net3916),
    .X(net4767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4241 (.A(net8352),
    .X(net4768));
 sky130_fd_sc_hd__clkbuf_2 hold4242 (.A(net3702),
    .X(net4769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4244 (.A(_02799_),
    .X(net4771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4245 (.A(_02804_),
    .X(net4772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4246 (.A(net8028),
    .X(net4773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4247 (.A(net3535),
    .X(net4774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4248 (.A(net8446),
    .X(net4775));
 sky130_fd_sc_hd__buf_2 hold4249 (.A(net3626),
    .X(net4776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(net5393),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_2 hold4250 (.A(net4660),
    .X(net4777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4251 (.A(_06091_),
    .X(net4778));
 sky130_fd_sc_hd__buf_1 hold4252 (.A(_06093_),
    .X(net4779));
 sky130_fd_sc_hd__buf_1 hold4253 (.A(net5976),
    .X(net4780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4254 (.A(_06160_),
    .X(net4781));
 sky130_fd_sc_hd__clkbuf_2 hold4255 (.A(_02319_),
    .X(net4782));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4257 (.A(_02561_),
    .X(net4784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4258 (.A(_02565_),
    .X(net4785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4259 (.A(net8050),
    .X(net4786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(net5359),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4260 (.A(net3515),
    .X(net4787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4261 (.A(net7928),
    .X(net4788));
 sky130_fd_sc_hd__buf_1 hold4262 (.A(net3637),
    .X(net4789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4264 (.A(_02618_),
    .X(net4791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4265 (.A(_02622_),
    .X(net4792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4266 (.A(_02624_),
    .X(net4793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4267 (.A(net8110),
    .X(net4794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4268 (.A(net1610),
    .X(net4795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(net5361),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4270 (.A(_02857_),
    .X(net4797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4271 (.A(_02861_),
    .X(net4798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4272 (.A(_02863_),
    .X(net4799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4273 (.A(net8114),
    .X(net4800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4274 (.A(net1676),
    .X(net4801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4275 (.A(\rbzero.pov.ready_buffer[12] ),
    .X(net4802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4276 (.A(net674),
    .X(net4803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4277 (.A(_01220_),
    .X(net4804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4278 (.A(net675),
    .X(net4805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(net5347),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4280 (.A(_02883_),
    .X(net4807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4281 (.A(_02884_),
    .X(net4808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4282 (.A(net8063),
    .X(net4809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4283 (.A(net3760),
    .X(net4810));
 sky130_fd_sc_hd__clkbuf_1 hold4284 (.A(net3972),
    .X(net4811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4285 (.A(net8052),
    .X(net4812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4286 (.A(net3973),
    .X(net4813));
 sky130_fd_sc_hd__clkbuf_2 hold4287 (.A(net5894),
    .X(net4814));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4288 (.A(_02474_),
    .X(net4815));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4289 (.A(_03427_),
    .X(net4816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(net5349),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4290 (.A(_00965_),
    .X(net4817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4291 (.A(net1022),
    .X(net4818));
 sky130_fd_sc_hd__buf_1 hold4293 (.A(_02644_),
    .X(net4820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4294 (.A(_02645_),
    .X(net4821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4295 (.A(net8087),
    .X(net4822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4296 (.A(net3948),
    .X(net4823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4297 (.A(\rbzero.pov.ready_buffer[1] ),
    .X(net4824));
 sky130_fd_sc_hd__buf_1 hold4298 (.A(net1941),
    .X(net4825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4299 (.A(_01231_),
    .X(net4826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(net7302),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4300 (.A(net1942),
    .X(net4827));
 sky130_fd_sc_hd__clkbuf_2 hold4301 (.A(net3529),
    .X(net4828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4302 (.A(_00610_),
    .X(net4829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4303 (.A(net3530),
    .X(net4830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4304 (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .X(net4831));
 sky130_fd_sc_hd__buf_1 hold4305 (.A(net3083),
    .X(net4832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4306 (.A(_02472_),
    .X(net4833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4307 (.A(_03386_),
    .X(net4834));
 sky130_fd_sc_hd__buf_1 hold4308 (.A(_03424_),
    .X(net4835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4309 (.A(_00963_),
    .X(net4836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(_03156_),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4310 (.A(net1032),
    .X(net4837));
 sky130_fd_sc_hd__clkbuf_2 hold4311 (.A(net3455),
    .X(net4838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4312 (.A(_00638_),
    .X(net4839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4313 (.A(net3456),
    .X(net4840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4314 (.A(\rbzero.spi_registers.got_new_texadd[2] ),
    .X(net4841));
 sky130_fd_sc_hd__clkbuf_2 hold4315 (.A(net1043),
    .X(net4842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4316 (.A(_03425_),
    .X(net4843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4317 (.A(net1044),
    .X(net4844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4318 (.A(_00964_),
    .X(net4845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4319 (.A(net1045),
    .X(net4846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(net4367),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4320 (.A(\rbzero.wall_tracer.rayAddendY[-6] ),
    .X(net4847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4321 (.A(net892),
    .X(net4848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4322 (.A(_01654_),
    .X(net4849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4323 (.A(net893),
    .X(net4850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4324 (.A(\rbzero.wall_tracer.rayAddendX[-6] ),
    .X(net4851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4325 (.A(net781),
    .X(net4852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4326 (.A(_01650_),
    .X(net4853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4327 (.A(net782),
    .X(net4854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4329 (.A(_02907_),
    .X(net4856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(net8125),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4330 (.A(_02908_),
    .X(net4857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4331 (.A(_02909_),
    .X(net4858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4332 (.A(_00636_),
    .X(net4859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4333 (.A(net3763),
    .X(net4860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4334 (.A(net5958),
    .X(net4861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4335 (.A(net3627),
    .X(net4862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4336 (.A(_04475_),
    .X(net4863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4337 (.A(_06055_),
    .X(net4864));
 sky130_fd_sc_hd__clkbuf_2 hold4338 (.A(_06056_),
    .X(net4865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net4278),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4340 (.A(_02669_),
    .X(net4867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4341 (.A(_02670_),
    .X(net4868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4342 (.A(_02671_),
    .X(net4869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4343 (.A(_00608_),
    .X(net4870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4344 (.A(net3616),
    .X(net4871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4345 (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .X(net4872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4346 (.A(net3944),
    .X(net4873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4347 (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(net4874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4348 (.A(net3931),
    .X(net4875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net5323),
    .X(net962));
 sky130_fd_sc_hd__buf_2 hold4350 (.A(_08462_),
    .X(net4877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4351 (.A(\rbzero.wall_tracer.rayAddendY[-7] ),
    .X(net4878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4352 (.A(net942),
    .X(net4879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4353 (.A(_01653_),
    .X(net4880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4354 (.A(net943),
    .X(net4881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4355 (.A(\rbzero.wall_tracer.rayAddendX[-5] ),
    .X(net4882));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4356 (.A(net917),
    .X(net4883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4357 (.A(_00596_),
    .X(net4884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4358 (.A(net918),
    .X(net4885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4359 (.A(\rbzero.wall_tracer.rayAddendX[-7] ),
    .X(net4886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(net5325),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4360 (.A(net789),
    .X(net4887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4361 (.A(_01649_),
    .X(net4888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4362 (.A(net790),
    .X(net4889));
 sky130_fd_sc_hd__clkbuf_1 hold4363 (.A(net4331),
    .X(net4890));
 sky130_fd_sc_hd__clkbuf_2 hold4364 (.A(net7817),
    .X(net4891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4366 (.A(net8364),
    .X(net4893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4368 (.A(net8402),
    .X(net4895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4369 (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .X(net4896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(net6113),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4370 (.A(net3668),
    .X(net4897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4371 (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .X(net4898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4372 (.A(net3784),
    .X(net4899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4373 (.A(\rbzero.pov.ready_buffer[53] ),
    .X(net4900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4374 (.A(net2426),
    .X(net4901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4375 (.A(_03685_),
    .X(net4902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4376 (.A(_01191_),
    .X(net4903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4377 (.A(net3327),
    .X(net4904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4378 (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .X(net4905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4379 (.A(net3767),
    .X(net4906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(net6115),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_1 hold4380 (.A(net4705),
    .X(net4907));
 sky130_fd_sc_hd__clkbuf_2 hold4381 (.A(_09223_),
    .X(net4908));
 sky130_fd_sc_hd__buf_1 hold4382 (.A(_09602_),
    .X(net4909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4383 (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .X(net4910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4384 (.A(net3765),
    .X(net4911));
 sky130_fd_sc_hd__buf_1 hold4385 (.A(net4674),
    .X(net4912));
 sky130_fd_sc_hd__clkbuf_2 hold4386 (.A(_09343_),
    .X(net4913));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4387 (.A(_10027_),
    .X(net4914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4388 (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .X(net4915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4389 (.A(net3756),
    .X(net4916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_01443_),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 hold4390 (.A(net4694),
    .X(net4917));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4391 (.A(_08130_),
    .X(net4918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4392 (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .X(net4919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4393 (.A(net3887),
    .X(net4920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4394 (.A(\gpout5.clk_div[0] ),
    .X(net4921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4395 (.A(net602),
    .X(net4922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4396 (.A(_01598_),
    .X(net4923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4397 (.A(net603),
    .X(net4924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4398 (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .X(net4925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4399 (.A(net3786),
    .X(net4926));
 sky130_fd_sc_hd__buf_1 hold440 (.A(net8234),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4400 (.A(\gpout3.clk_div[0] ),
    .X(net4927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4401 (.A(net593),
    .X(net4928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4402 (.A(_01659_),
    .X(net4929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4403 (.A(net594),
    .X(net4930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4404 (.A(\gpout0.clk_div[0] ),
    .X(net4931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4405 (.A(net595),
    .X(net4932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4406 (.A(_01645_),
    .X(net4933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4407 (.A(net596),
    .X(net4934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4408 (.A(\gpout4.clk_div[0] ),
    .X(net4935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4409 (.A(net600),
    .X(net4936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net7922),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4410 (.A(_01661_),
    .X(net4937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4411 (.A(net601),
    .X(net4938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4412 (.A(\gpout1.clk_div[0] ),
    .X(net4939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4413 (.A(net604),
    .X(net4940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4414 (.A(_01655_),
    .X(net4941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4415 (.A(net605),
    .X(net4942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4416 (.A(\rbzero.pov.spi_counter[6] ),
    .X(net4943));
 sky130_fd_sc_hd__buf_1 hold4417 (.A(net614),
    .X(net4944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4418 (.A(_01021_),
    .X(net4945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4419 (.A(net615),
    .X(net4946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net8233),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4420 (.A(\gpout2.clk_div[0] ),
    .X(net4947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4421 (.A(net608),
    .X(net4948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4422 (.A(_01657_),
    .X(net4949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4423 (.A(net609),
    .X(net4950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4424 (.A(\rbzero.color_floor[3] ),
    .X(net4951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4425 (.A(net606),
    .X(net4952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4426 (.A(_00894_),
    .X(net4953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4427 (.A(net607),
    .X(net4954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4428 (.A(\rbzero.color_floor[5] ),
    .X(net4955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4429 (.A(net612),
    .X(net4956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(net8017),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4430 (.A(_00896_),
    .X(net4957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4431 (.A(net613),
    .X(net4958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4432 (.A(\rbzero.color_floor[1] ),
    .X(net4959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4433 (.A(net619),
    .X(net4960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4434 (.A(_00892_),
    .X(net4961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4435 (.A(net620),
    .X(net4962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4436 (.A(\rbzero.color_sky[2] ),
    .X(net4963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4437 (.A(net621),
    .X(net4964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4438 (.A(_00887_),
    .X(net4965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4439 (.A(net622),
    .X(net4966));
 sky130_fd_sc_hd__buf_1 hold444 (.A(net8221),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4440 (.A(\rbzero.texV[-11] ),
    .X(net4967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4441 (.A(net640),
    .X(net4968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4442 (.A(_01600_),
    .X(net4969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4443 (.A(net641),
    .X(net4970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4444 (.A(\rbzero.texV[-2] ),
    .X(net4971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4445 (.A(net648),
    .X(net4972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4446 (.A(_01609_),
    .X(net4973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4447 (.A(net649),
    .X(net4974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4448 (.A(\rbzero.spi_registers.texadd3[23] ),
    .X(net4975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4449 (.A(net705),
    .X(net4976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(net8070),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4450 (.A(_00878_),
    .X(net4977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4451 (.A(net706),
    .X(net4978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4452 (.A(\rbzero.texV[-1] ),
    .X(net4979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4453 (.A(net650),
    .X(net4980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4454 (.A(net8198),
    .X(net4981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4455 (.A(net651),
    .X(net4982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4456 (.A(\rbzero.texV[-10] ),
    .X(net4983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4457 (.A(net658),
    .X(net4984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4458 (.A(_01601_),
    .X(net4985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4459 (.A(net659),
    .X(net4986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(net5279),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4460 (.A(\rbzero.spi_registers.texadd3[20] ),
    .X(net4987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4461 (.A(net715),
    .X(net4988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4462 (.A(_00875_),
    .X(net4989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4463 (.A(net716),
    .X(net4990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4464 (.A(\rbzero.spi_registers.texadd3[3] ),
    .X(net4991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4465 (.A(net668),
    .X(net4992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4466 (.A(_00858_),
    .X(net4993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4467 (.A(net669),
    .X(net4994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4469 (.A(\rbzero.pov.ready ),
    .X(net4996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(net5281),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4470 (.A(net670),
    .X(net4997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4471 (.A(_01014_),
    .X(net4998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4472 (.A(net671),
    .X(net4999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4473 (.A(\rbzero.spi_registers.texadd3[13] ),
    .X(net5000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4474 (.A(net729),
    .X(net5001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4475 (.A(_00868_),
    .X(net5002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4476 (.A(net730),
    .X(net5003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4477 (.A(\rbzero.spi_registers.texadd0[3] ),
    .X(net5004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4478 (.A(net697),
    .X(net5005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4479 (.A(_00786_),
    .X(net5006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(net2796),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4480 (.A(net698),
    .X(net5007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4481 (.A(\rbzero.spi_registers.texadd3[11] ),
    .X(net5008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4482 (.A(net727),
    .X(net5009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4483 (.A(_00866_),
    .X(net5010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4484 (.A(net728),
    .X(net5011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4485 (.A(\rbzero.spi_registers.texadd2[20] ),
    .X(net5012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4486 (.A(net687),
    .X(net5013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4487 (.A(_00851_),
    .X(net5014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4488 (.A(net688),
    .X(net5015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4489 (.A(\rbzero.spi_registers.texadd3[0] ),
    .X(net5016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(_04069_),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4490 (.A(net685),
    .X(net5017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4491 (.A(_00855_),
    .X(net5018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4492 (.A(net686),
    .X(net5019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4493 (.A(\rbzero.spi_registers.texadd3[10] ),
    .X(net5020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4494 (.A(net748),
    .X(net5021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4495 (.A(_00865_),
    .X(net5022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4496 (.A(net749),
    .X(net5023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4497 (.A(\rbzero.spi_registers.texadd3[12] ),
    .X(net5024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4498 (.A(net717),
    .X(net5025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4499 (.A(_00867_),
    .X(net5026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_01563_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4500 (.A(net718),
    .X(net5027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4501 (.A(\rbzero.spi_registers.texadd1[7] ),
    .X(net5028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4502 (.A(net699),
    .X(net5029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4503 (.A(_00814_),
    .X(net5030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4504 (.A(net700),
    .X(net5031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4505 (.A(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(net5032));
 sky130_fd_sc_hd__buf_1 hold4506 (.A(net666),
    .X(net5033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4507 (.A(_01647_),
    .X(net5034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4508 (.A(net667),
    .X(net5035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4509 (.A(\rbzero.spi_registers.texadd1[21] ),
    .X(net5036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(net5351),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4510 (.A(net703),
    .X(net5037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4511 (.A(_00828_),
    .X(net5038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4512 (.A(net704),
    .X(net5039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4513 (.A(\rbzero.spi_registers.texadd3[1] ),
    .X(net5040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4514 (.A(net709),
    .X(net5041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4515 (.A(_00856_),
    .X(net5042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4516 (.A(net710),
    .X(net5043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4517 (.A(\rbzero.pov.ready_buffer[10] ),
    .X(net5044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4518 (.A(net610),
    .X(net5045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4519 (.A(_01240_),
    .X(net5046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(net5353),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4520 (.A(net611),
    .X(net5047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4521 (.A(\rbzero.color_sky[4] ),
    .X(net5048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4522 (.A(net691),
    .X(net5049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4523 (.A(_00889_),
    .X(net5050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4524 (.A(net692),
    .X(net5051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4525 (.A(\rbzero.spi_registers.texadd0[1] ),
    .X(net5052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4526 (.A(net713),
    .X(net5053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4527 (.A(_00784_),
    .X(net5054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4528 (.A(net714),
    .X(net5055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4529 (.A(\rbzero.spi_registers.texadd1[20] ),
    .X(net5056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(net5371),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4530 (.A(net689),
    .X(net5057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4531 (.A(_00827_),
    .X(net5058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4532 (.A(net690),
    .X(net5059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4533 (.A(\rbzero.spi_registers.texadd1[9] ),
    .X(net5060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4534 (.A(net826),
    .X(net5061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4535 (.A(_00816_),
    .X(net5062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4536 (.A(net827),
    .X(net5063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4537 (.A(\rbzero.spi_registers.texadd0[16] ),
    .X(net5064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4538 (.A(net719),
    .X(net5065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4539 (.A(_00799_),
    .X(net5066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(net5373),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4540 (.A(net720),
    .X(net5067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4541 (.A(\rbzero.spi_registers.texadd2[21] ),
    .X(net5068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4542 (.A(net707),
    .X(net5069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4543 (.A(_00852_),
    .X(net5070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4544 (.A(net708),
    .X(net5071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4545 (.A(\rbzero.spi_registers.texadd2[8] ),
    .X(net5072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4546 (.A(net725),
    .X(net5073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4547 (.A(_00839_),
    .X(net5074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4548 (.A(net726),
    .X(net5075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4549 (.A(\rbzero.spi_registers.texadd1[8] ),
    .X(net5076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(net5271),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4550 (.A(net701),
    .X(net5077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4551 (.A(_00815_),
    .X(net5078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4552 (.A(net702),
    .X(net5079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4553 (.A(\rbzero.spi_registers.texadd0[4] ),
    .X(net5080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4554 (.A(net711),
    .X(net5081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4555 (.A(_00787_),
    .X(net5082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4556 (.A(net712),
    .X(net5083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4557 (.A(\rbzero.spi_registers.texadd2[11] ),
    .X(net5084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4558 (.A(net695),
    .X(net5085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4559 (.A(_00842_),
    .X(net5086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(net5273),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4560 (.A(net696),
    .X(net5087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4561 (.A(\rbzero.spi_registers.texadd1[23] ),
    .X(net5088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4562 (.A(net842),
    .X(net5089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4563 (.A(_00830_),
    .X(net5090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4564 (.A(net843),
    .X(net5091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4565 (.A(\rbzero.spi_registers.texadd0[0] ),
    .X(net5092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4566 (.A(net723),
    .X(net5093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4567 (.A(_00783_),
    .X(net5094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4568 (.A(net724),
    .X(net5095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4569 (.A(\rbzero.spi_registers.texadd1[4] ),
    .X(net5096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(net8180),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4570 (.A(net733),
    .X(net5097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4571 (.A(_00811_),
    .X(net5098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4572 (.A(net734),
    .X(net5099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4573 (.A(\rbzero.spi_registers.texadd3[14] ),
    .X(net5100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4574 (.A(net742),
    .X(net5101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4575 (.A(_00869_),
    .X(net5102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4576 (.A(net743),
    .X(net5103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4577 (.A(\rbzero.spi_registers.texadd3[8] ),
    .X(net5104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4578 (.A(net795),
    .X(net5105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4579 (.A(_00863_),
    .X(net5106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(net8031),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4580 (.A(net796),
    .X(net5107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4581 (.A(\rbzero.spi_registers.texadd1[17] ),
    .X(net5108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4582 (.A(net797),
    .X(net5109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4583 (.A(_00824_),
    .X(net5110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4584 (.A(net798),
    .X(net5111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4585 (.A(\rbzero.spi_registers.texadd3[4] ),
    .X(net5112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4586 (.A(net769),
    .X(net5113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4587 (.A(_00859_),
    .X(net5114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4588 (.A(net770),
    .X(net5115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4589 (.A(\rbzero.spi_registers.texadd2[6] ),
    .X(net5116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(net6471),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4590 (.A(net760),
    .X(net5117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4591 (.A(_00837_),
    .X(net5118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4592 (.A(net761),
    .X(net5119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4593 (.A(\rbzero.spi_registers.texadd0[14] ),
    .X(net5120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4594 (.A(net731),
    .X(net5121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4595 (.A(_00797_),
    .X(net5122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4596 (.A(net732),
    .X(net5123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4597 (.A(\rbzero.spi_registers.texadd1[2] ),
    .X(net5124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4598 (.A(net752),
    .X(net5125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4599 (.A(_00809_),
    .X(net5126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_03223_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4600 (.A(net753),
    .X(net5127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4601 (.A(\rbzero.spi_registers.texadd2[0] ),
    .X(net5128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4602 (.A(net721),
    .X(net5129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4603 (.A(_00831_),
    .X(net5130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4604 (.A(net722),
    .X(net5131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4605 (.A(\rbzero.spi_registers.texadd2[18] ),
    .X(net5132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4606 (.A(net773),
    .X(net5133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4607 (.A(_00849_),
    .X(net5134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4608 (.A(net774),
    .X(net5135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4609 (.A(\rbzero.spi_registers.texadd2[9] ),
    .X(net5136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(net4208),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4610 (.A(net787),
    .X(net5137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4611 (.A(_00840_),
    .X(net5138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4612 (.A(net788),
    .X(net5139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4613 (.A(\rbzero.spi_registers.texadd1[5] ),
    .X(net5140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4614 (.A(net738),
    .X(net5141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4615 (.A(_00812_),
    .X(net5142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4616 (.A(net739),
    .X(net5143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4617 (.A(\rbzero.spi_registers.texadd1[12] ),
    .X(net5144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4618 (.A(net771),
    .X(net5145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4619 (.A(_00819_),
    .X(net5146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(net5411),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4620 (.A(net772),
    .X(net5147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4621 (.A(\rbzero.spi_registers.texadd0[17] ),
    .X(net5148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4622 (.A(net764),
    .X(net5149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4623 (.A(_00800_),
    .X(net5150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4624 (.A(net765),
    .X(net5151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4625 (.A(\rbzero.spi_registers.texadd3[16] ),
    .X(net5152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4626 (.A(net785),
    .X(net5153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4627 (.A(_00871_),
    .X(net5154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4628 (.A(net786),
    .X(net5155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4629 (.A(\rbzero.mapdxw[0] ),
    .X(net5156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(net5413),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4630 (.A(net740),
    .X(net5157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4631 (.A(_00779_),
    .X(net5158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4632 (.A(net741),
    .X(net5159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4633 (.A(\rbzero.spi_registers.texadd2[2] ),
    .X(net5160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4634 (.A(net793),
    .X(net5161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4635 (.A(_00833_),
    .X(net5162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4636 (.A(net794),
    .X(net5163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4637 (.A(\rbzero.spi_registers.texadd0[18] ),
    .X(net5164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4638 (.A(net907),
    .X(net5165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4639 (.A(_00801_),
    .X(net5166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(net8199),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4640 (.A(net908),
    .X(net5167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4641 (.A(\rbzero.spi_registers.texadd1[13] ),
    .X(net5168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4642 (.A(net812),
    .X(net5169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4643 (.A(_00820_),
    .X(net5170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4644 (.A(net813),
    .X(net5171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4645 (.A(\rbzero.spi_registers.texadd3[17] ),
    .X(net5172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4646 (.A(net808),
    .X(net5173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4647 (.A(_00872_),
    .X(net5174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4648 (.A(net809),
    .X(net5175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4649 (.A(\rbzero.spi_registers.texadd2[15] ),
    .X(net5176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(net8090),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4650 (.A(net783),
    .X(net5177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4651 (.A(_00846_),
    .X(net5178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4652 (.A(net784),
    .X(net5179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4653 (.A(\rbzero.spi_registers.texadd2[16] ),
    .X(net5180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4654 (.A(net828),
    .X(net5181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4655 (.A(_00847_),
    .X(net5182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4656 (.A(net829),
    .X(net5183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4657 (.A(\rbzero.spi_registers.texadd0[5] ),
    .X(net5184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4658 (.A(net862),
    .X(net5185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4659 (.A(_00788_),
    .X(net5186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(net5287),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4660 (.A(net863),
    .X(net5187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4661 (.A(\rbzero.spi_registers.texadd3[18] ),
    .X(net5188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4662 (.A(net882),
    .X(net5189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4663 (.A(_00873_),
    .X(net5190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4664 (.A(net883),
    .X(net5191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4665 (.A(\rbzero.spi_registers.texadd3[2] ),
    .X(net5192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4666 (.A(net750),
    .X(net5193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4667 (.A(_00857_),
    .X(net5194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4668 (.A(net751),
    .X(net5195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4669 (.A(\rbzero.spi_registers.texadd3[19] ),
    .X(net5196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(net5289),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4670 (.A(net880),
    .X(net5197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4671 (.A(_00874_),
    .X(net5198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4672 (.A(net881),
    .X(net5199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4673 (.A(\rbzero.spi_registers.texadd2[4] ),
    .X(net5200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4674 (.A(net844),
    .X(net5201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4675 (.A(_00835_),
    .X(net5202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4676 (.A(net845),
    .X(net5203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4677 (.A(\gpout0.hpos[6] ),
    .X(net5204));
 sky130_fd_sc_hd__buf_2 hold4678 (.A(net3516),
    .X(net5205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4679 (.A(_04501_),
    .X(net5206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(net5395),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4680 (.A(_03790_),
    .X(net5207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4681 (.A(_03791_),
    .X(net5208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4682 (.A(_01243_),
    .X(net5209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4683 (.A(net3643),
    .X(net5210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4684 (.A(\rbzero.spi_registers.texadd0[10] ),
    .X(net5211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4685 (.A(net824),
    .X(net5212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4686 (.A(_00793_),
    .X(net5213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4687 (.A(net825),
    .X(net5214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4688 (.A(\rbzero.spi_registers.texadd2[5] ),
    .X(net5215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4689 (.A(net858),
    .X(net5216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net5397),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4690 (.A(_00836_),
    .X(net5217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4691 (.A(net859),
    .X(net5218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4692 (.A(\rbzero.spi_registers.texadd0[19] ),
    .X(net5219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4693 (.A(net927),
    .X(net5220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4694 (.A(_00802_),
    .X(net5221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4695 (.A(net928),
    .X(net5222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4696 (.A(\rbzero.spi_registers.texadd3[15] ),
    .X(net5223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4697 (.A(net820),
    .X(net5224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4698 (.A(_00870_),
    .X(net5225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4699 (.A(net821),
    .X(net5226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(net6117),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4700 (.A(\rbzero.spi_registers.texadd1[6] ),
    .X(net5227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4701 (.A(net852),
    .X(net5228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4702 (.A(_00813_),
    .X(net5229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4703 (.A(net853),
    .X(net5230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4704 (.A(\rbzero.spi_registers.texadd0[15] ),
    .X(net5231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4705 (.A(net870),
    .X(net5232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4706 (.A(_00798_),
    .X(net5233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4707 (.A(net871),
    .X(net5234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4708 (.A(\rbzero.spi_registers.texadd0[2] ),
    .X(net5235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4709 (.A(net936),
    .X(net5236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(net6119),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4710 (.A(_00785_),
    .X(net5237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4711 (.A(net937),
    .X(net5238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4712 (.A(\rbzero.spi_registers.texadd0[8] ),
    .X(net5239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4713 (.A(net799),
    .X(net5240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4714 (.A(_00791_),
    .X(net5241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4715 (.A(net800),
    .X(net5242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4716 (.A(\rbzero.spi_registers.texadd0[12] ),
    .X(net5243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4717 (.A(net806),
    .X(net5244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4718 (.A(_00795_),
    .X(net5245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4719 (.A(net807),
    .X(net5246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_01323_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4720 (.A(\rbzero.spi_registers.texadd3[21] ),
    .X(net5247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4721 (.A(net818),
    .X(net5248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4722 (.A(_00876_),
    .X(net5249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4723 (.A(net819),
    .X(net5250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4724 (.A(\rbzero.texV[-5] ),
    .X(net5251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4725 (.A(net866),
    .X(net5252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4726 (.A(_01606_),
    .X(net5253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4727 (.A(net867),
    .X(net5254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4728 (.A(\rbzero.spi_registers.texadd0[7] ),
    .X(net5255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4729 (.A(net922),
    .X(net5256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(net5343),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4730 (.A(_00790_),
    .X(net5257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4731 (.A(net923),
    .X(net5258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4732 (.A(\rbzero.spi_registers.texadd2[10] ),
    .X(net5259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4733 (.A(net758),
    .X(net5260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4734 (.A(_00841_),
    .X(net5261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4735 (.A(net759),
    .X(net5262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4736 (.A(\rbzero.spi_registers.texadd1[0] ),
    .X(net5263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4737 (.A(net860),
    .X(net5264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4738 (.A(_00807_),
    .X(net5265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4739 (.A(net861),
    .X(net5266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(net5345),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4740 (.A(\rbzero.spi_registers.texadd2[3] ),
    .X(net5267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4741 (.A(net801),
    .X(net5268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4742 (.A(_00834_),
    .X(net5269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4743 (.A(net802),
    .X(net5270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4744 (.A(\rbzero.spi_registers.texadd3[22] ),
    .X(net5271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4745 (.A(net982),
    .X(net5272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4746 (.A(_00877_),
    .X(net5273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4747 (.A(net983),
    .X(net5274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4748 (.A(\rbzero.spi_registers.texadd2[17] ),
    .X(net5275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4749 (.A(net898),
    .X(net5276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(net8128),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4750 (.A(_00848_),
    .X(net5277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4751 (.A(net899),
    .X(net5278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4752 (.A(\rbzero.pov.spi_counter[0] ),
    .X(net5279));
 sky130_fd_sc_hd__buf_1 hold4753 (.A(net973),
    .X(net5280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4754 (.A(_01015_),
    .X(net5281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4755 (.A(net974),
    .X(net5282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4756 (.A(\rbzero.spi_registers.texadd1[16] ),
    .X(net5283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4757 (.A(net878),
    .X(net5284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4758 (.A(_00823_),
    .X(net5285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4759 (.A(net879),
    .X(net5286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(net4532),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4760 (.A(\rbzero.spi_registers.texadd3[9] ),
    .X(net5287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4761 (.A(net993),
    .X(net5288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4762 (.A(_00864_),
    .X(net5289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4763 (.A(net994),
    .X(net5290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4764 (.A(\rbzero.spi_registers.texadd0[11] ),
    .X(net5291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4765 (.A(net911),
    .X(net5292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4766 (.A(_00794_),
    .X(net5293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4767 (.A(net912),
    .X(net5294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4768 (.A(\rbzero.spi_registers.texadd2[7] ),
    .X(net5295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4769 (.A(net902),
    .X(net5296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(net5415),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4770 (.A(_00838_),
    .X(net5297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4771 (.A(net903),
    .X(net5298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4772 (.A(\rbzero.spi_registers.texadd2[12] ),
    .X(net5299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4773 (.A(net856),
    .X(net5300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4774 (.A(_00843_),
    .X(net5301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4775 (.A(net857),
    .X(net5302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4776 (.A(\rbzero.spi_registers.texadd2[22] ),
    .X(net5303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4777 (.A(net814),
    .X(net5304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4778 (.A(_00853_),
    .X(net5305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4779 (.A(net815),
    .X(net5306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(net5417),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4780 (.A(\rbzero.spi_registers.texadd1[18] ),
    .X(net5307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4781 (.A(net909),
    .X(net5308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4782 (.A(_00825_),
    .X(net5309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4783 (.A(net910),
    .X(net5310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4784 (.A(\rbzero.spi_registers.texadd3[7] ),
    .X(net5311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4785 (.A(net931),
    .X(net5312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4786 (.A(_00862_),
    .X(net5313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4787 (.A(net932),
    .X(net5314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4788 (.A(\rbzero.spi_registers.texadd2[13] ),
    .X(net5315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4789 (.A(net874),
    .X(net5316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(net5427),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4790 (.A(_00844_),
    .X(net5317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4791 (.A(net875),
    .X(net5318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4792 (.A(\rbzero.spi_registers.texadd1[15] ),
    .X(net5319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4793 (.A(net944),
    .X(net5320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4794 (.A(_00822_),
    .X(net5321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4795 (.A(net945),
    .X(net5322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4796 (.A(\rbzero.spi_registers.texadd0[9] ),
    .X(net5323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4797 (.A(net962),
    .X(net5324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4798 (.A(_00792_),
    .X(net5325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4799 (.A(net963),
    .X(net5326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(net5429),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4800 (.A(\rbzero.wall_tracer.mapX[10] ),
    .X(net5327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4801 (.A(net832),
    .X(net5328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4802 (.A(_00527_),
    .X(net5329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4803 (.A(net833),
    .X(net5330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4804 (.A(\rbzero.spi_registers.texadd1[1] ),
    .X(net5331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4805 (.A(net868),
    .X(net5332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4806 (.A(_00808_),
    .X(net5333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4807 (.A(net869),
    .X(net5334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4808 (.A(\rbzero.spi_registers.texadd0[20] ),
    .X(net5335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4809 (.A(net913),
    .X(net5336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(net7891),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4810 (.A(_00803_),
    .X(net5337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4811 (.A(net914),
    .X(net5338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4812 (.A(\rbzero.texV[-4] ),
    .X(net5339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4813 (.A(net915),
    .X(net5340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4814 (.A(_01607_),
    .X(net5341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4815 (.A(net916),
    .X(net5342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4816 (.A(\rbzero.spi_registers.texadd2[23] ),
    .X(net5343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4817 (.A(net1000),
    .X(net5344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4818 (.A(_00854_),
    .X(net5345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4819 (.A(net1001),
    .X(net5346));
 sky130_fd_sc_hd__buf_1 hold482 (.A(net8223),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4820 (.A(\rbzero.spi_registers.texadd0[21] ),
    .X(net5347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4821 (.A(net955),
    .X(net5348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4822 (.A(_00804_),
    .X(net5349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4823 (.A(net956),
    .X(net5350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4824 (.A(\rbzero.spi_registers.texadd1[3] ),
    .X(net5351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4825 (.A(net978),
    .X(net5352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4826 (.A(_00810_),
    .X(net5353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4827 (.A(net979),
    .X(net5354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4828 (.A(\rbzero.color_sky[0] ),
    .X(net5355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4829 (.A(net846),
    .X(net5356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(net8014),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4830 (.A(_00885_),
    .X(net5357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4831 (.A(net847),
    .X(net5358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4832 (.A(\rbzero.spi_registers.texadd3[5] ),
    .X(net5359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4833 (.A(net953),
    .X(net5360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4834 (.A(_00860_),
    .X(net5361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4835 (.A(net954),
    .X(net5362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4836 (.A(\rbzero.spi_registers.texadd0[6] ),
    .X(net5363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4837 (.A(net929),
    .X(net5364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4838 (.A(_00789_),
    .X(net5365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4839 (.A(net930),
    .X(net5366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(net5387),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4840 (.A(\rbzero.spi_registers.texadd1[22] ),
    .X(net5367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4841 (.A(net946),
    .X(net5368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4842 (.A(_00829_),
    .X(net5369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4843 (.A(net947),
    .X(net5370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4844 (.A(\rbzero.spi_registers.texadd0[13] ),
    .X(net5371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4845 (.A(net980),
    .X(net5372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4846 (.A(_00796_),
    .X(net5373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4847 (.A(net981),
    .X(net5374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4848 (.A(\rbzero.texV[-3] ),
    .X(net5375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4849 (.A(net884),
    .X(net5376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(net5389),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4850 (.A(_01608_),
    .X(net5377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4851 (.A(net885),
    .X(net5378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4852 (.A(\rbzero.texV[-7] ),
    .X(net5379));
 sky130_fd_sc_hd__buf_1 hold4853 (.A(net854),
    .X(net5380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4854 (.A(_01604_),
    .X(net5381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4855 (.A(net855),
    .X(net5382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4856 (.A(\rbzero.texV[-9] ),
    .X(net5383));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4857 (.A(net848),
    .X(net5384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4858 (.A(_01602_),
    .X(net5385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4859 (.A(net849),
    .X(net5386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(net5419),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4860 (.A(\rbzero.spi_registers.texadd1[10] ),
    .X(net5387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4861 (.A(net1011),
    .X(net5388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4862 (.A(_00817_),
    .X(net5389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4863 (.A(net1012),
    .X(net5390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4864 (.A(\rbzero.mapdyw[1] ),
    .X(net5391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4865 (.A(net951),
    .X(net5392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4866 (.A(_00782_),
    .X(net5393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4867 (.A(net952),
    .X(net5394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4868 (.A(\rbzero.spi_registers.texadd3[6] ),
    .X(net5395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4869 (.A(net995),
    .X(net5396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(net5421),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4870 (.A(_00861_),
    .X(net5397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4871 (.A(net996),
    .X(net5398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4872 (.A(\rbzero.texV[-8] ),
    .X(net5399));
 sky130_fd_sc_hd__buf_1 hold4873 (.A(net872),
    .X(net5400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4874 (.A(_01603_),
    .X(net5401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4875 (.A(net873),
    .X(net5402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4876 (.A(\rbzero.texV[-6] ),
    .X(net5403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4877 (.A(net830),
    .X(net5404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4878 (.A(_01605_),
    .X(net5405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4879 (.A(net831),
    .X(net5406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(net8228),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4880 (.A(\rbzero.wall_tracer.mapY[10] ),
    .X(net5407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4881 (.A(net894),
    .X(net5408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4882 (.A(_00390_),
    .X(net5409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4883 (.A(net895),
    .X(net5410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4884 (.A(\rbzero.spi_registers.texadd1[19] ),
    .X(net5411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4885 (.A(net989),
    .X(net5412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4886 (.A(_00826_),
    .X(net5413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4887 (.A(net990),
    .X(net5414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4888 (.A(\rbzero.mapdxw[1] ),
    .X(net5415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4889 (.A(net1004),
    .X(net5416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(net8004),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4890 (.A(_00780_),
    .X(net5417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4891 (.A(net1005),
    .X(net5418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4892 (.A(\rbzero.mapdyw[0] ),
    .X(net5419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4893 (.A(net1013),
    .X(net5420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4894 (.A(_00781_),
    .X(net5421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4895 (.A(net1014),
    .X(net5422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4896 (.A(\rbzero.spi_registers.texadd1[11] ),
    .X(net5423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4897 (.A(net1036),
    .X(net5424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4898 (.A(_00818_),
    .X(net5425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4899 (.A(net1037),
    .X(net5426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(net6127),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4900 (.A(\rbzero.wall_tracer.mapY[8] ),
    .X(net5427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4901 (.A(net1006),
    .X(net5428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4902 (.A(_00388_),
    .X(net5429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4903 (.A(net1007),
    .X(net5430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4904 (.A(\rbzero.map_overlay.i_mapdx[5] ),
    .X(net5431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4905 (.A(net1024),
    .X(net5432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4906 (.A(_00772_),
    .X(net5433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4907 (.A(net1025),
    .X(net5434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4908 (.A(\rbzero.spi_registers.texadd0[22] ),
    .X(net5435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4909 (.A(net1087),
    .X(net5436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(net6129),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4910 (.A(_00805_),
    .X(net5437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4911 (.A(net1088),
    .X(net5438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4912 (.A(\rbzero.floor_leak[0] ),
    .X(net5439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4913 (.A(net1050),
    .X(net5440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4914 (.A(_00879_),
    .X(net5441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4915 (.A(net1051),
    .X(net5442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4916 (.A(\rbzero.spi_registers.texadd0[23] ),
    .X(net5443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4917 (.A(net1067),
    .X(net5444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4918 (.A(_00806_),
    .X(net5445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4919 (.A(net1068),
    .X(net5446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_01303_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4920 (.A(\rbzero.texV[0] ),
    .X(net5447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4921 (.A(net1046),
    .X(net5448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4922 (.A(net8182),
    .X(net5449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4923 (.A(net1047),
    .X(net5450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4924 (.A(\rbzero.spi_registers.vshift[5] ),
    .X(net5451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4925 (.A(net1122),
    .X(net5452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4926 (.A(_00902_),
    .X(net5453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4927 (.A(net1123),
    .X(net5454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4928 (.A(\rbzero.spi_registers.texadd2[14] ),
    .X(net5455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4929 (.A(net1118),
    .X(net5456));
 sky130_fd_sc_hd__buf_1 hold493 (.A(net8174),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4930 (.A(_00845_),
    .X(net5457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4931 (.A(net1119),
    .X(net5458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4932 (.A(\rbzero.floor_leak[1] ),
    .X(net5459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4933 (.A(net1136),
    .X(net5460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4934 (.A(_00880_),
    .X(net5461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4935 (.A(net1137),
    .X(net5462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4936 (.A(\rbzero.spi_registers.vshift[4] ),
    .X(net5463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4937 (.A(net1156),
    .X(net5464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4938 (.A(_00901_),
    .X(net5465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4939 (.A(net1157),
    .X(net5466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_03426_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4940 (.A(\rbzero.map_overlay.i_mapdy[5] ),
    .X(net5467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4941 (.A(net1163),
    .X(net5468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4942 (.A(_00778_),
    .X(net5469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4943 (.A(net1164),
    .X(net5470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4944 (.A(\rbzero.wall_tracer.mapX[8] ),
    .X(net5471));
 sky130_fd_sc_hd__buf_1 hold4945 (.A(net1161),
    .X(net5472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4946 (.A(_00525_),
    .X(net5473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4947 (.A(net1162),
    .X(net5474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4948 (.A(\rbzero.pov.ready_buffer[21] ),
    .X(net5475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4949 (.A(net1108),
    .X(net5476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(net4817),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4950 (.A(_01229_),
    .X(net5477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4951 (.A(net1109),
    .X(net5478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4952 (.A(\rbzero.texV[9] ),
    .X(net5479));
 sky130_fd_sc_hd__buf_1 hold4953 (.A(net1228),
    .X(net5480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4954 (.A(_01620_),
    .X(net5481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4955 (.A(net1229),
    .X(net5482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4956 (.A(\rbzero.floor_leak[2] ),
    .X(net5483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4957 (.A(net1209),
    .X(net5484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4958 (.A(_00881_),
    .X(net5485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4959 (.A(net1210),
    .X(net5486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(net7888),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4960 (.A(\rbzero.texV[2] ),
    .X(net5487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4961 (.A(net1217),
    .X(net5488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4962 (.A(_01613_),
    .X(net5489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4963 (.A(net1218),
    .X(net5490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4964 (.A(\rbzero.texV[1] ),
    .X(net5491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4965 (.A(net1233),
    .X(net5492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4966 (.A(_01612_),
    .X(net5493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4967 (.A(net1234),
    .X(net5494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4968 (.A(\rbzero.pov.spi_counter[2] ),
    .X(net5495));
 sky130_fd_sc_hd__buf_1 hold4969 (.A(net1253),
    .X(net5496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(net5431),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4970 (.A(_01017_),
    .X(net5497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4971 (.A(net1254),
    .X(net5498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4972 (.A(\rbzero.spi_registers.new_leak[3] ),
    .X(net5499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4973 (.A(net1634),
    .X(net5500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4974 (.A(_03307_),
    .X(net5501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4975 (.A(_00882_),
    .X(net5502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4976 (.A(net1256),
    .X(net5503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4977 (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .X(net5504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4978 (.A(net3982),
    .X(net5505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4979 (.A(_00771_),
    .X(net5506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net5433),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4980 (.A(net1135),
    .X(net5507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4981 (.A(\rbzero.floor_leak[5] ),
    .X(net5508));
 sky130_fd_sc_hd__buf_1 hold4982 (.A(net1414),
    .X(net5509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4983 (.A(_00884_),
    .X(net5510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4984 (.A(net1415),
    .X(net5511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4985 (.A(\rbzero.spi_registers.new_vshift[1] ),
    .X(net5512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4986 (.A(net1582),
    .X(net5513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4987 (.A(_03337_),
    .X(net5514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4988 (.A(_00898_),
    .X(net5515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4989 (.A(net1659),
    .X(net5516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(net3361),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4990 (.A(\rbzero.floor_leak[4] ),
    .X(net5517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4991 (.A(net1550),
    .X(net5518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4992 (.A(_00883_),
    .X(net5519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4993 (.A(net1551),
    .X(net5520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4994 (.A(\rbzero.texV[6] ),
    .X(net5521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4995 (.A(net1284),
    .X(net5522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4996 (.A(net8230),
    .X(net5523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4997 (.A(net1285),
    .X(net5524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4998 (.A(\rbzero.spi_registers.new_other[0] ),
    .X(net5525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4999 (.A(net1640),
    .X(net5526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net4464),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5000 (.A(_03133_),
    .X(net5527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5001 (.A(_00761_),
    .X(net5528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5002 (.A(net1818),
    .X(net5529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5003 (.A(\rbzero.wall_tracer.mapY[7] ),
    .X(net5530));
 sky130_fd_sc_hd__buf_1 hold5004 (.A(net1611),
    .X(net5531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5005 (.A(_00387_),
    .X(net5532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5006 (.A(net1612),
    .X(net5533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5007 (.A(\rbzero.spi_registers.new_other[4] ),
    .X(net5534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5008 (.A(net1700),
    .X(net5535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5009 (.A(_03137_),
    .X(net5536));
 sky130_fd_sc_hd__buf_1 hold501 (.A(net8066),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5010 (.A(_00765_),
    .X(net5537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5011 (.A(net1804),
    .X(net5538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5012 (.A(\rbzero.spi_registers.new_other[1] ),
    .X(net5539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5013 (.A(net1736),
    .X(net5540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5014 (.A(_03134_),
    .X(net5541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5015 (.A(_00762_),
    .X(net5542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5016 (.A(net2039),
    .X(net5543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5017 (.A(\rbzero.tex_r0[10] ),
    .X(net5544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5018 (.A(_04165_),
    .X(net5545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5019 (.A(net2123),
    .X(net5546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(net4266),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5020 (.A(\rbzero.tex_r1[28] ),
    .X(net5547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5021 (.A(_04071_),
    .X(net5548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5022 (.A(net2153),
    .X(net5549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5023 (.A(\rbzero.tex_r1[1] ),
    .X(net5550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5024 (.A(_04100_),
    .X(net5551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5025 (.A(net1530),
    .X(net5552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5026 (.A(\rbzero.wall_tracer.mapX[6] ),
    .X(net5553));
 sky130_fd_sc_hd__buf_1 hold5027 (.A(net2006),
    .X(net5554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5028 (.A(_00523_),
    .X(net5555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5029 (.A(net2007),
    .X(net5556));
 sky130_fd_sc_hd__buf_1 hold503 (.A(net8194),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5030 (.A(\rbzero.tex_r1[0] ),
    .X(net5557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5031 (.A(net1275),
    .X(net5558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5032 (.A(_04101_),
    .X(net5559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5033 (.A(net1276),
    .X(net5560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5034 (.A(\rbzero.spi_registers.new_vshift[2] ),
    .X(net5561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5035 (.A(net1402),
    .X(net5562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5036 (.A(_03338_),
    .X(net5563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5037 (.A(_00899_),
    .X(net5564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5038 (.A(net1852),
    .X(net5565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5039 (.A(\rbzero.tex_b0[1] ),
    .X(net5566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_03423_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5040 (.A(_04457_),
    .X(net5567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5041 (.A(net1837),
    .X(net5568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5042 (.A(\rbzero.spi_registers.new_other[10] ),
    .X(net5569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5043 (.A(net1764),
    .X(net5570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5044 (.A(_03132_),
    .X(net5571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5045 (.A(_00760_),
    .X(net5572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5046 (.A(net2186),
    .X(net5573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5047 (.A(\rbzero.tex_b1[60] ),
    .X(net5574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5048 (.A(_04323_),
    .X(net5575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5049 (.A(net2286),
    .X(net5576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(net4836),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5050 (.A(\rbzero.tex_r0[48] ),
    .X(net5577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5051 (.A(_04123_),
    .X(net5578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5052 (.A(net2582),
    .X(net5579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5053 (.A(\rbzero.texV[4] ),
    .X(net5580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5054 (.A(net1616),
    .X(net5581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5055 (.A(net8210),
    .X(net5582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5056 (.A(net1617),
    .X(net5583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5057 (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .X(net5584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5058 (.A(net3874),
    .X(net5585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5059 (.A(\rbzero.tex_b1[14] ),
    .X(net5586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(net6612),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5060 (.A(_04373_),
    .X(net5587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5061 (.A(net2884),
    .X(net5588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5062 (.A(\rbzero.tex_b1[32] ),
    .X(net5589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5063 (.A(_04354_),
    .X(net5590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5064 (.A(net2215),
    .X(net5591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5065 (.A(\rbzero.tex_b1[28] ),
    .X(net5592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5066 (.A(_04358_),
    .X(net5593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5067 (.A(net1989),
    .X(net5594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5068 (.A(\rbzero.row_render.texu[4] ),
    .X(net5595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5069 (.A(net1822),
    .X(net5596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_03336_),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5070 (.A(_00498_),
    .X(net5597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5071 (.A(net5676),
    .X(net5598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5072 (.A(_04060_),
    .X(net5599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5073 (.A(net2041),
    .X(net5600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5074 (.A(\rbzero.tex_r0[2] ),
    .X(net5601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5075 (.A(_04174_),
    .X(net5602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5076 (.A(net2794),
    .X(net5603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5077 (.A(\rbzero.wall_tracer.mapY[6] ),
    .X(net5604));
 sky130_fd_sc_hd__buf_1 hold5078 (.A(net2277),
    .X(net5605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5079 (.A(_00386_),
    .X(net5606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(net4313),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5080 (.A(net2278),
    .X(net5607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5081 (.A(\rbzero.texV[10] ),
    .X(net5608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5082 (.A(net1918),
    .X(net5609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5083 (.A(_01621_),
    .X(net5610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5084 (.A(net1919),
    .X(net5611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5085 (.A(\rbzero.spi_registers.new_mapd[4] ),
    .X(net5612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5086 (.A(net2104),
    .X(net5613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5087 (.A(_03155_),
    .X(net5614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5088 (.A(_00773_),
    .X(net5615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5089 (.A(net2588),
    .X(net5616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(net5423),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5090 (.A(\rbzero.wall_tracer.mapY[9] ),
    .X(net5617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5091 (.A(net2058),
    .X(net5618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5092 (.A(_00389_),
    .X(net5619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5093 (.A(net2059),
    .X(net5620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5094 (.A(\rbzero.texV[3] ),
    .X(net5621));
 sky130_fd_sc_hd__buf_1 hold5095 (.A(net2474),
    .X(net5622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5096 (.A(_01614_),
    .X(net5623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5097 (.A(net2475),
    .X(net5624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5098 (.A(\rbzero.tex_b0[2] ),
    .X(net5625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5099 (.A(net2835),
    .X(net5626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(net5425),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5100 (.A(_04456_),
    .X(net5627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5101 (.A(net2836),
    .X(net5628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5102 (.A(\rbzero.tex_r0[3] ),
    .X(net5629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5103 (.A(net1748),
    .X(net5630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5104 (.A(_04173_),
    .X(net5631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5105 (.A(net1749),
    .X(net5632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5106 (.A(\rbzero.tex_b1[33] ),
    .X(net5633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5107 (.A(net1949),
    .X(net5634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5108 (.A(_04352_),
    .X(net5635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5109 (.A(net1950),
    .X(net5636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(net8208),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5110 (.A(\rbzero.tex_r1[32] ),
    .X(net5637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5111 (.A(_04067_),
    .X(net5638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5112 (.A(net2374),
    .X(net5639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5113 (.A(\rbzero.tex_g0[1] ),
    .X(net5640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5114 (.A(_04316_),
    .X(net5641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5115 (.A(net656),
    .X(net5642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5116 (.A(_01343_),
    .X(net5643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5117 (.A(\rbzero.tex_r1[33] ),
    .X(net5644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5118 (.A(net2250),
    .X(net5645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5119 (.A(_04066_),
    .X(net5646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(net8011),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5120 (.A(net2251),
    .X(net5647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5121 (.A(\rbzero.tex_b1[29] ),
    .X(net5648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5122 (.A(net2823),
    .X(net5649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5123 (.A(_04357_),
    .X(net5650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5124 (.A(net2824),
    .X(net5651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5125 (.A(\rbzero.tex_b1[61] ),
    .X(net5652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5126 (.A(net2134),
    .X(net5653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5127 (.A(_04322_),
    .X(net5654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5128 (.A(net2135),
    .X(net5655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5129 (.A(\rbzero.hsync ),
    .X(net5656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(net6139),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5130 (.A(net900),
    .X(net5657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5131 (.A(_01632_),
    .X(net5658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5132 (.A(\rbzero.tex_r1[15] ),
    .X(net5659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5133 (.A(_04085_),
    .X(net5660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5134 (.A(net2343),
    .X(net5661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5135 (.A(net5699),
    .X(net5662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5136 (.A(_04244_),
    .X(net5663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5137 (.A(net2463),
    .X(net5664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5138 (.A(\rbzero.wall_tracer.mapX[7] ),
    .X(net5665));
 sky130_fd_sc_hd__buf_1 hold5139 (.A(net2379),
    .X(net5666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(net6141),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5140 (.A(_00524_),
    .X(net5667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5141 (.A(net2380),
    .X(net5668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5142 (.A(\rbzero.tex_b1[48] ),
    .X(net5669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5143 (.A(_04336_),
    .X(net5670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5144 (.A(net2623),
    .X(net5671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5145 (.A(\rbzero.tex_b1[15] ),
    .X(net5672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5146 (.A(net2306),
    .X(net5673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5147 (.A(_04372_),
    .X(net5674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5148 (.A(net2307),
    .X(net5675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5149 (.A(\rbzero.tex_r1[38] ),
    .X(net5676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_01583_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5150 (.A(net5598),
    .X(net5677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5151 (.A(_04059_),
    .X(net5678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5152 (.A(net3241),
    .X(net5679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5153 (.A(\rbzero.tex_b1[2] ),
    .X(net5680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5154 (.A(_04386_),
    .X(net5681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5155 (.A(net2352),
    .X(net5682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5156 (.A(\rbzero.tex_b1[3] ),
    .X(net5683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5157 (.A(net2703),
    .X(net5684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5158 (.A(_04385_),
    .X(net5685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5159 (.A(net2704),
    .X(net5686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net4841),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5160 (.A(\rbzero.tex_r0[11] ),
    .X(net5687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5161 (.A(net1124),
    .X(net5688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5162 (.A(_04164_),
    .X(net5689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5163 (.A(net1125),
    .X(net5690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5164 (.A(\rbzero.texV[5] ),
    .X(net5691));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold5165 (.A(net2494),
    .X(net5692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5166 (.A(_01616_),
    .X(net5693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5167 (.A(net2495),
    .X(net5694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5168 (.A(\rbzero.tex_r1[29] ),
    .X(net5695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5169 (.A(net3114),
    .X(net5696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(net4843),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5170 (.A(_04070_),
    .X(net5697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5171 (.A(net3115),
    .X(net5698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5172 (.A(\rbzero.tex_g1[2] ),
    .X(net5699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5173 (.A(net5662),
    .X(net5700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5174 (.A(_04245_),
    .X(net5701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5175 (.A(net3105),
    .X(net5702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5176 (.A(\rbzero.pov.ready_buffer[45] ),
    .X(net5703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5177 (.A(net4616),
    .X(net5704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5178 (.A(\rbzero.tex_r0[49] ),
    .X(net5705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5179 (.A(net1438),
    .X(net5706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(net4845),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5180 (.A(_04122_),
    .X(net5707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5181 (.A(net1439),
    .X(net5708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5182 (.A(\rbzero.pov.spi_buffer[50] ),
    .X(net5709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5183 (.A(net2193),
    .X(net5710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5184 (.A(_03049_),
    .X(net5711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5185 (.A(net2194),
    .X(net5712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5186 (.A(\rbzero.tex_g0[0] ),
    .X(net5713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5187 (.A(net2697),
    .X(net5714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5188 (.A(_04317_),
    .X(net5715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5189 (.A(net2698),
    .X(net5716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net5447),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5190 (.A(\rbzero.tex_b1[49] ),
    .X(net5717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5191 (.A(net2990),
    .X(net5718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5192 (.A(_04335_),
    .X(net5719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5193 (.A(net2991),
    .X(net5720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5194 (.A(\rbzero.wall_tracer.mapX[9] ),
    .X(net5721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5195 (.A(net2968),
    .X(net5722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5196 (.A(_00526_),
    .X(net5723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5197 (.A(net2969),
    .X(net5724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5198 (.A(\rbzero.texV[7] ),
    .X(net5725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5199 (.A(net2753),
    .X(net5726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net5449),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5200 (.A(_01618_),
    .X(net5727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5201 (.A(net2754),
    .X(net5728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5202 (.A(\rbzero.tex_r1[16] ),
    .X(net5729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5203 (.A(net2741),
    .X(net5730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5204 (.A(_04084_),
    .X(net5731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5205 (.A(net2742),
    .X(net5732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5206 (.A(net5758),
    .X(net5733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5207 (.A(_03057_),
    .X(net5734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5208 (.A(net2941),
    .X(net5735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5209 (.A(\rbzero.pov.ready_buffer[56] ),
    .X(net5736));
 sky130_fd_sc_hd__buf_1 hold521 (.A(net8131),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5210 (.A(net4374),
    .X(net5737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5211 (.A(\rbzero.texV[8] ),
    .X(net5738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5212 (.A(net3189),
    .X(net5739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5213 (.A(_01619_),
    .X(net5740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5214 (.A(net3190),
    .X(net5741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5215 (.A(\rbzero.pov.ready_buffer[49] ),
    .X(net5742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5216 (.A(net4362),
    .X(net5743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5217 (.A(\rbzero.pov.ready_buffer[59] ),
    .X(net5744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5218 (.A(net3098),
    .X(net5745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5219 (.A(_03612_),
    .X(net5746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(net4269),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5220 (.A(_01167_),
    .X(net5747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5221 (.A(net3387),
    .X(net5748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5222 (.A(\rbzero.pov.ready_buffer[47] ),
    .X(net5749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5223 (.A(net1906),
    .X(net5750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5224 (.A(_03670_),
    .X(net5751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5225 (.A(_01185_),
    .X(net5752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5226 (.A(net3373),
    .X(net5753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5227 (.A(\rbzero.map_overlay.i_otherx[0] ),
    .X(net5754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5228 (.A(net4152),
    .X(net5755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5229 (.A(_00756_),
    .X(net5756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(net5439),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5230 (.A(net2630),
    .X(net5757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5231 (.A(\rbzero.pov.ready_buffer[58] ),
    .X(net5758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5232 (.A(net5733),
    .X(net5759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5233 (.A(_03704_),
    .X(net5760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5234 (.A(_03705_),
    .X(net5761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5235 (.A(net3470),
    .X(net5762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5236 (.A(\rbzero.pov.spi_buffer[70] ),
    .X(net5763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5237 (.A(net1979),
    .X(net5764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5238 (.A(_03070_),
    .X(net5765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5239 (.A(net1980),
    .X(net5766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(net5441),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5240 (.A(\rbzero.debug_overlay.playerX[-4] ),
    .X(net5767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5241 (.A(net3339),
    .X(net5768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5242 (.A(_09327_),
    .X(net5769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5243 (.A(\rbzero.pov.ready_buffer[51] ),
    .X(net5770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5244 (.A(net3323),
    .X(net5771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5245 (.A(_03678_),
    .X(net5772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5246 (.A(_01189_),
    .X(net5773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5247 (.A(net3446),
    .X(net5774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5249 (.A(_02878_),
    .X(net5776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(net6155),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5250 (.A(net3464),
    .X(net5777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5251 (.A(_00633_),
    .X(net5778));
 sky130_fd_sc_hd__clkbuf_1 hold5252 (.A(net3967),
    .X(net5779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5253 (.A(net8218),
    .X(net5780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5254 (.A(net3968),
    .X(net5781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5255 (.A(\rbzero.pov.ready_buffer[64] ),
    .X(net5782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5256 (.A(net4441),
    .X(net5783));
 sky130_fd_sc_hd__buf_1 hold5257 (.A(net7691),
    .X(net5784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5258 (.A(_03073_),
    .X(net5785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5259 (.A(net1614),
    .X(net5786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net6157),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5260 (.A(\rbzero.tex_r1[40] ),
    .X(net5787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5261 (.A(net584),
    .X(net5788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5262 (.A(_04058_),
    .X(net5789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5263 (.A(net585),
    .X(net5790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5264 (.A(net5906),
    .X(net5791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5265 (.A(_03069_),
    .X(net5792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5266 (.A(net3192),
    .X(net5793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5268 (.A(_02819_),
    .X(net5795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5269 (.A(net3499),
    .X(net5796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(_01061_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5270 (.A(_00629_),
    .X(net5797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5271 (.A(\rbzero.spi_registers.spi_counter[5] ),
    .X(net5798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5272 (.A(net1250),
    .X(net5799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5273 (.A(_02986_),
    .X(net5800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5274 (.A(_00645_),
    .X(net5801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5275 (.A(net1252),
    .X(net5802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5277 (.A(_02798_),
    .X(net5804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5278 (.A(net3524),
    .X(net5805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5279 (.A(_00627_),
    .X(net5806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(net7543),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5281 (.A(_02788_),
    .X(net5808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5282 (.A(net3527),
    .X(net5809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5283 (.A(_00626_),
    .X(net5810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5284 (.A(\rbzero.pov.spi_buffer[66] ),
    .X(net5811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5285 (.A(net1709),
    .X(net5812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5286 (.A(_03066_),
    .X(net5813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5287 (.A(net1710),
    .X(net5814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5288 (.A(\rbzero.pov.ready_buffer[60] ),
    .X(net5815));
 sky130_fd_sc_hd__buf_1 hold5289 (.A(net1535),
    .X(net5816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net4488),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5290 (.A(_03616_),
    .X(net5817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5291 (.A(_03617_),
    .X(net5818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5292 (.A(_01168_),
    .X(net5819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5293 (.A(net3537),
    .X(net5820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5295 (.A(_02548_),
    .X(net5822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5296 (.A(net3635),
    .X(net5823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5297 (.A(_00598_),
    .X(net5824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5298 (.A(\rbzero.pov.ready_buffer[67] ),
    .X(net5825));
 sky130_fd_sc_hd__buf_1 hold5299 (.A(net1703),
    .X(net5826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\rbzero.pov.ready_buffer[23] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5300 (.A(_03633_),
    .X(net5827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5301 (.A(_01175_),
    .X(net5828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5302 (.A(net2899),
    .X(net5829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5304 (.A(_02558_),
    .X(net5831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5305 (.A(net3716),
    .X(net5832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5306 (.A(_00599_),
    .X(net5833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5307 (.A(\rbzero.pov.ready_buffer[61] ),
    .X(net5834));
 sky130_fd_sc_hd__buf_1 hold5308 (.A(net3411),
    .X(net5835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5309 (.A(_03618_),
    .X(net5836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net7946),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5310 (.A(_03619_),
    .X(net5837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5311 (.A(_01169_),
    .X(net5838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5312 (.A(net3349),
    .X(net5839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5314 (.A(_02903_),
    .X(net5841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5315 (.A(net3742),
    .X(net5842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5316 (.A(_00635_),
    .X(net5843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5317 (.A(\rbzero.spi_registers.spi_counter[0] ),
    .X(net5844));
 sky130_fd_sc_hd__clkbuf_2 hold5318 (.A(net2198),
    .X(net5845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5319 (.A(_00640_),
    .X(net5846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(net7551),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5320 (.A(net2200),
    .X(net5847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5321 (.A(\rbzero.pov.ready_buffer[65] ),
    .X(net5848));
 sky130_fd_sc_hd__buf_1 hold5322 (.A(net3266),
    .X(net5849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5323 (.A(_03626_),
    .X(net5850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5324 (.A(_03627_),
    .X(net5851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5325 (.A(_01173_),
    .X(net5852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5326 (.A(net3458),
    .X(net5853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5328 (.A(_02844_),
    .X(net5855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5329 (.A(net3753),
    .X(net5856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(net4468),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5330 (.A(_00631_),
    .X(net5857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5331 (.A(\rbzero.debug_overlay.playerY[-7] ),
    .X(net5858));
 sky130_fd_sc_hd__clkbuf_2 hold5332 (.A(net3315),
    .X(net5859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5333 (.A(_01184_),
    .X(net5860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5334 (.A(net3316),
    .X(net5861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5335 (.A(\rbzero.spi_registers.sclk_buffer[2] ),
    .X(net5862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5336 (.A(net3041),
    .X(net5863));
 sky130_fd_sc_hd__buf_1 hold5337 (.A(_02972_),
    .X(net5864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5338 (.A(_00644_),
    .X(net5865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5339 (.A(net3487),
    .X(net5866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net6493),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5340 (.A(\rbzero.pov.ready_buffer[68] ),
    .X(net5867));
 sky130_fd_sc_hd__buf_1 hold5341 (.A(net3279),
    .X(net5868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5342 (.A(_03637_),
    .X(net5869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5343 (.A(_01176_),
    .X(net5870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5344 (.A(net3444),
    .X(net5871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5346 (.A(_02639_),
    .X(net5873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5347 (.A(net3813),
    .X(net5874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5348 (.A(_00605_),
    .X(net5875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5349 (.A(\rbzero.spi_registers.spi_counter[1] ),
    .X(net5876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_03135_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5350 (.A(net3909),
    .X(net5877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5351 (.A(_02971_),
    .X(net5878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5352 (.A(_02976_),
    .X(net5879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5353 (.A(_00642_),
    .X(net5880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5354 (.A(net1549),
    .X(net5881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5356 (.A(_02580_),
    .X(net5883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5357 (.A(net3828),
    .X(net5884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5358 (.A(_00601_),
    .X(net5885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5359 (.A(\rbzero.debug_overlay.playerX[-6] ),
    .X(net5886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(net4325),
    .X(net1063));
 sky130_fd_sc_hd__buf_2 hold5360 (.A(net3370),
    .X(net5887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5361 (.A(_01170_),
    .X(net5888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5362 (.A(net3371),
    .X(net5889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5364 (.A(_02665_),
    .X(net5891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5365 (.A(net3891),
    .X(net5892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5366 (.A(_00607_),
    .X(net5893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5367 (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .X(net5894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5368 (.A(net4814),
    .X(net5895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5369 (.A(_03108_),
    .X(net5896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(net6143),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5370 (.A(\rbzero.pov.ready_buffer[71] ),
    .X(net5897));
 sky130_fd_sc_hd__buf_1 hold5371 (.A(net3015),
    .X(net5898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5372 (.A(_03649_),
    .X(net5899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5373 (.A(_01179_),
    .X(net5900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5374 (.A(net3432),
    .X(net5901));
 sky130_fd_sc_hd__clkbuf_4 hold5375 (.A(_06757_),
    .X(net5902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5376 (.A(\rbzero.debug_overlay.playerX[-5] ),
    .X(net5903));
 sky130_fd_sc_hd__buf_1 hold5377 (.A(net3419),
    .X(net5904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5378 (.A(_01171_),
    .X(net5905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5379 (.A(\rbzero.pov.ready_buffer[69] ),
    .X(net5906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(net6145),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5380 (.A(net5791),
    .X(net5907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5381 (.A(_03639_),
    .X(net5908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5382 (.A(_03641_),
    .X(net5909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5383 (.A(\gpout0.hpos[5] ),
    .X(net5910));
 sky130_fd_sc_hd__buf_1 hold5384 (.A(net4105),
    .X(net5911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5385 (.A(_05067_),
    .X(net5912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5386 (.A(_05069_),
    .X(net5913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5387 (.A(\rbzero.debug_overlay.playerX[2] ),
    .X(net5914));
 sky130_fd_sc_hd__buf_1 hold5388 (.A(net3389),
    .X(net5915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5389 (.A(_04686_),
    .X(net5916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_01543_),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5390 (.A(_02738_),
    .X(net5917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5391 (.A(_02739_),
    .X(net5918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5392 (.A(_00620_),
    .X(net5919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5393 (.A(net3966),
    .X(net5920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5394 (.A(\rbzero.trace_state[3] ),
    .X(net5921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5395 (.A(net3870),
    .X(net5922));
 sky130_fd_sc_hd__buf_1 hold5396 (.A(_03989_),
    .X(net5923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5397 (.A(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(net5924));
 sky130_fd_sc_hd__buf_1 hold5398 (.A(net3308),
    .X(net5925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5399 (.A(_02778_),
    .X(net5926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(net5443),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5400 (.A(net3309),
    .X(net5927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5401 (.A(\rbzero.debug_overlay.playerY[-9] ),
    .X(net5928));
 sky130_fd_sc_hd__clkbuf_2 hold5402 (.A(net3417),
    .X(net5929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5403 (.A(_01182_),
    .X(net5930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5404 (.A(\rbzero.spi_registers.got_new_floor ),
    .X(net5931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5405 (.A(\rbzero.map_rom.b6 ),
    .X(net5932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5406 (.A(net3848),
    .X(net5933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5407 (.A(_02718_),
    .X(net5934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5408 (.A(net3849),
    .X(net5935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5409 (.A(\rbzero.map_rom.c6 ),
    .X(net5936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(net5445),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5410 (.A(net4641),
    .X(net5937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5411 (.A(_02714_),
    .X(net5938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5412 (.A(\rbzero.spi_registers.got_new_sky ),
    .X(net5939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5413 (.A(net3902),
    .X(net5940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5414 (.A(_03353_),
    .X(net5941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5415 (.A(\rbzero.spi_registers.got_new_other ),
    .X(net5942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5416 (.A(net3623),
    .X(net5943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5417 (.A(_03385_),
    .X(net5944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5418 (.A(\gpout0.hpos[3] ),
    .X(net5945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5419 (.A(net3917),
    .X(net5946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(net6183),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5420 (.A(_04462_),
    .X(net5947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5421 (.A(_05185_),
    .X(net5948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5422 (.A(_09729_),
    .X(net5949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5423 (.A(_00481_),
    .X(net5950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5424 (.A(net4090),
    .X(net5951));
 sky130_fd_sc_hd__clkbuf_2 hold5425 (.A(net3778),
    .X(net5952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5426 (.A(_02708_),
    .X(net5953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5427 (.A(net3779),
    .X(net5954));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold5428 (.A(net3611),
    .X(net5955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5429 (.A(_02946_),
    .X(net5956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(net6185),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5430 (.A(net3612),
    .X(net5957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5431 (.A(\rbzero.trace_state[0] ),
    .X(net5958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5432 (.A(net4861),
    .X(net5959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5433 (.A(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(net5960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5434 (.A(net3141),
    .X(net5961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5435 (.A(_02538_),
    .X(net5962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5436 (.A(net3142),
    .X(net5963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5437 (.A(\gpout0.vpos[8] ),
    .X(net5964));
 sky130_fd_sc_hd__buf_2 hold5438 (.A(net4065),
    .X(net5965));
 sky130_fd_sc_hd__buf_1 hold5439 (.A(_05730_),
    .X(net5966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_01293_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5440 (.A(\rbzero.row_render.side ),
    .X(net5967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5441 (.A(net4079),
    .X(net5968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5442 (.A(_05013_),
    .X(net5969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5444 (.A(_02605_),
    .X(net5971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5445 (.A(net3605),
    .X(net5972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5446 (.A(\rbzero.map_rom.d6 ),
    .X(net5973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5447 (.A(net3893),
    .X(net5974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5448 (.A(_06145_),
    .X(net5975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5449 (.A(_06159_),
    .X(net5976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(net6171),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5450 (.A(\rbzero.spi_registers.got_new_leak ),
    .X(net5977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5451 (.A(net3217),
    .X(net5978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5452 (.A(_03372_),
    .X(net5979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5453 (.A(\gpout0.vpos[1] ),
    .X(net5980));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold5454 (.A(net4023),
    .X(net5981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5455 (.A(_05678_),
    .X(net5982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5456 (.A(_03784_),
    .X(net5983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5457 (.A(_03785_),
    .X(net5984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5458 (.A(_01242_),
    .X(net5985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5459 (.A(net3338),
    .X(net5986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(net6173),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5460 (.A(\rbzero.pov.spi_buffer[68] ),
    .X(net5987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5461 (.A(net587),
    .X(net5988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5462 (.A(_03593_),
    .X(net5989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5463 (.A(\rbzero.tex_r0[4] ),
    .X(net5990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5464 (.A(net590),
    .X(net5991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5465 (.A(_04172_),
    .X(net5992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5466 (.A(\rbzero.spi_registers.new_sky[0] ),
    .X(net5993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5467 (.A(net1733),
    .X(net5994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5468 (.A(\rbzero.spi_registers.new_sky[2] ),
    .X(net5995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5469 (.A(net2321),
    .X(net5996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_01513_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5470 (.A(_03348_),
    .X(net5997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5471 (.A(net2322),
    .X(net5998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5472 (.A(\gpout0.vpos[0] ),
    .X(net5999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5473 (.A(net4101),
    .X(net6000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5474 (.A(_03795_),
    .X(net6001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5475 (.A(\rbzero.spi_registers.new_sky[3] ),
    .X(net6002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5476 (.A(net1724),
    .X(net6003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5477 (.A(\rbzero.spi_registers.new_sky[4] ),
    .X(net6004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5478 (.A(net2441),
    .X(net6005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5479 (.A(\rbzero.spi_registers.new_sky[5] ),
    .X(net6006));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold548 (.A(net7897),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5480 (.A(net2060),
    .X(net6007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5481 (.A(_03351_),
    .X(net6008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5482 (.A(\rbzero.spi_registers.new_floor[2] ),
    .X(net6009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5483 (.A(net1564),
    .X(net6010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5484 (.A(_03357_),
    .X(net6011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5485 (.A(net1565),
    .X(net6012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5486 (.A(\rbzero.spi_registers.new_sky[1] ),
    .X(net6013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5487 (.A(net1532),
    .X(net6014));
 sky130_fd_sc_hd__clkbuf_2 hold5488 (.A(net3734),
    .X(net6015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5489 (.A(_02694_),
    .X(net6016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(net6485),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5490 (.A(net3735),
    .X(net6017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5491 (.A(\rbzero.spi_registers.new_floor[0] ),
    .X(net6018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5492 (.A(net1480),
    .X(net6019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5493 (.A(\rbzero.spi_registers.new_floor[5] ),
    .X(net6020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5494 (.A(net1561),
    .X(net6021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5495 (.A(_03360_),
    .X(net6022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5496 (.A(\rbzero.spi_registers.new_floor[4] ),
    .X(net6023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5497 (.A(net2232),
    .X(net6024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5498 (.A(\rbzero.tex_b0[60] ),
    .X(net6025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5499 (.A(net623),
    .X(net6026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_03136_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5500 (.A(_04393_),
    .X(net6027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5501 (.A(net624),
    .X(net6028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5502 (.A(\rbzero.tex_b0[20] ),
    .X(net6029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5503 (.A(net633),
    .X(net6030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5504 (.A(_04437_),
    .X(net6031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5505 (.A(net634),
    .X(net6032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5506 (.A(\rbzero.tex_g1[8] ),
    .X(net6033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5507 (.A(net630),
    .X(net6034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5508 (.A(_04239_),
    .X(net6035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5509 (.A(net631),
    .X(net6036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(net4307),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5510 (.A(\gpout0.hpos[0] ),
    .X(net6037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5511 (.A(net3641),
    .X(net6038));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold5512 (.A(_04020_),
    .X(net6039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5513 (.A(\gpout2.clk_div[1] ),
    .X(net6040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5514 (.A(net678),
    .X(net6041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5515 (.A(_04017_),
    .X(net6042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5516 (.A(\gpout0.vpos[9] ),
    .X(net6043));
 sky130_fd_sc_hd__buf_2 hold5517 (.A(net3995),
    .X(net6044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5518 (.A(_01253_),
    .X(net6045));
 sky130_fd_sc_hd__clkbuf_2 hold5519 (.A(net3601),
    .X(net6046));
 sky130_fd_sc_hd__buf_1 hold552 (.A(net8302),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5520 (.A(_02932_),
    .X(net6047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5521 (.A(net3602),
    .X(net6048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5522 (.A(\rbzero.spi_registers.new_floor[1] ),
    .X(net6049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5523 (.A(net1593),
    .X(net6050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5524 (.A(\rbzero.tex_b1[6] ),
    .X(net6051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5525 (.A(net660),
    .X(net6052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5526 (.A(_04382_),
    .X(net6053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5527 (.A(net661),
    .X(net6054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5528 (.A(\rbzero.spi_registers.new_floor[3] ),
    .X(net6055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5529 (.A(net1625),
    .X(net6056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(net6163),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5530 (.A(\gpout5.clk_div[1] ),
    .X(net6057));
 sky130_fd_sc_hd__clkbuf_2 hold5531 (.A(net919),
    .X(net6058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5532 (.A(_03873_),
    .X(net6059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5533 (.A(\rbzero.pov.ready_buffer[57] ),
    .X(net6060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5534 (.A(net3038),
    .X(net6061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5535 (.A(_03702_),
    .X(net6062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5536 (.A(net3554),
    .X(net6063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5537 (.A(\rbzero.spi_registers.got_new_mapd ),
    .X(net6064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5538 (.A(net886),
    .X(net6065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5539 (.A(_03420_),
    .X(net6066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(net6165),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5540 (.A(\rbzero.spi_registers.new_texadd[1][20] ),
    .X(net6067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5541 (.A(net2075),
    .X(net6068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5542 (.A(_03479_),
    .X(net6069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5543 (.A(net2076),
    .X(net6070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5544 (.A(\rbzero.tex_g0[32] ),
    .X(net6071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5545 (.A(net642),
    .X(net6072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5546 (.A(_04283_),
    .X(net6073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5547 (.A(net643),
    .X(net6074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5548 (.A(\rbzero.spi_registers.new_texadd[1][21] ),
    .X(net6075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5549 (.A(net2414),
    .X(net6076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_01383_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5550 (.A(_03480_),
    .X(net6077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5551 (.A(net2415),
    .X(net6078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5552 (.A(\rbzero.spi_registers.new_texadd[3][21] ),
    .X(net6079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5553 (.A(net1590),
    .X(net6080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5554 (.A(_03837_),
    .X(net6081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5555 (.A(net1591),
    .X(net6082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5556 (.A(\rbzero.tex_r0[24] ),
    .X(net6083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5557 (.A(net766),
    .X(net6084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5558 (.A(_04150_),
    .X(net6085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5559 (.A(net767),
    .X(net6086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(net6167),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5560 (.A(\rbzero.tex_r1[20] ),
    .X(net6087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5561 (.A(net933),
    .X(net6088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5562 (.A(_04080_),
    .X(net6089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5563 (.A(net934),
    .X(net6090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5564 (.A(\rbzero.tex_g0[52] ),
    .X(net6091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5565 (.A(net803),
    .X(net6092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5566 (.A(_04260_),
    .X(net6093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5567 (.A(net804),
    .X(net6094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5568 (.A(\rbzero.tex_b0[30] ),
    .X(net6095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5569 (.A(net904),
    .X(net6096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(net6169),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5570 (.A(_04426_),
    .X(net6097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5571 (.A(net905),
    .X(net6098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5572 (.A(\gpout1.clk_div[1] ),
    .X(net6099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5573 (.A(net1095),
    .X(net6100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5574 (.A(_04016_),
    .X(net6101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5575 (.A(\rbzero.tex_b0[50] ),
    .X(net6102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5576 (.A(net938),
    .X(net6103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5577 (.A(_04404_),
    .X(net6104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5578 (.A(net939),
    .X(net6105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5579 (.A(\rbzero.tex_g0[22] ),
    .X(net6106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_01433_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5580 (.A(net924),
    .X(net6107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5581 (.A(_04294_),
    .X(net6108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5582 (.A(net925),
    .X(net6109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5583 (.A(\gpout4.clk_div[1] ),
    .X(net6110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5584 (.A(net1098),
    .X(net6111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5585 (.A(_04019_),
    .X(net6112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5586 (.A(\rbzero.tex_g1[38] ),
    .X(net6113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5587 (.A(net964),
    .X(net6114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5588 (.A(_04206_),
    .X(net6115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5589 (.A(net965),
    .X(net6116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net7894),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5590 (.A(\rbzero.tex_b1[46] ),
    .X(net6117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5591 (.A(net997),
    .X(net6118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5592 (.A(_04338_),
    .X(net6119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5593 (.A(net998),
    .X(net6120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5594 (.A(\gpout0.clk_div[1] ),
    .X(net6121));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold5595 (.A(net1092),
    .X(net6122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5596 (.A(_04003_),
    .X(net6123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5597 (.A(\rbzero.pov.spi_buffer[19] ),
    .X(net6124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5598 (.A(net735),
    .X(net6125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5599 (.A(_03540_),
    .X(net6126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(net5435),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5600 (.A(\rbzero.tex_b1[26] ),
    .X(net6127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5601 (.A(net1017),
    .X(net6128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5602 (.A(_04360_),
    .X(net6129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5603 (.A(net1018),
    .X(net6130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5604 (.A(\rbzero.spi_registers.new_texadd[1][22] ),
    .X(net6131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5605 (.A(net2137),
    .X(net6132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5606 (.A(_03481_),
    .X(net6133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5607 (.A(net2138),
    .X(net6134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5608 (.A(\rbzero.spi_registers.new_texadd[3][20] ),
    .X(net6135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5609 (.A(net1399),
    .X(net6136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(net5437),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5610 (.A(_03836_),
    .X(net6137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5611 (.A(net1400),
    .X(net6138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5612 (.A(\rbzero.tex_r1[50] ),
    .X(net6139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5613 (.A(net1040),
    .X(net6140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5614 (.A(_04047_),
    .X(net6141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5615 (.A(net1041),
    .X(net6142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5616 (.A(\rbzero.tex_r1[10] ),
    .X(net6143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5617 (.A(net1064),
    .X(net6144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5618 (.A(_04091_),
    .X(net6145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5619 (.A(net1065),
    .X(net6146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(net6151),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5620 (.A(\rbzero.spi_registers.new_texadd[2][21] ),
    .X(net6147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5621 (.A(net1505),
    .X(net6148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5622 (.A(_02505_),
    .X(net6149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5623 (.A(net1506),
    .X(net6150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5624 (.A(\rbzero.tex_r0[14] ),
    .X(net6151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5625 (.A(net1089),
    .X(net6152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5626 (.A(_04161_),
    .X(net6153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5627 (.A(net1090),
    .X(net6154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5628 (.A(\rbzero.tex_b0[40] ),
    .X(net6155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5629 (.A(net1052),
    .X(net6156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(net6153),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5630 (.A(_04415_),
    .X(net6157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5631 (.A(net1053),
    .X(net6158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5632 (.A(\rbzero.spi_registers.new_texadd[2][22] ),
    .X(net6159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5633 (.A(net1599),
    .X(net6160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5634 (.A(_02506_),
    .X(net6161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5635 (.A(net1600),
    .X(net6162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5636 (.A(\rbzero.tex_g0[42] ),
    .X(net6163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5637 (.A(net1080),
    .X(net6164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5638 (.A(_04272_),
    .X(net6165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5639 (.A(net1081),
    .X(net6166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_01483_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5640 (.A(\rbzero.tex_g1[28] ),
    .X(net6167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5641 (.A(net1083),
    .X(net6168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5642 (.A(_04217_),
    .X(net6169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5643 (.A(net1084),
    .X(net6170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5644 (.A(\rbzero.tex_r0[44] ),
    .X(net6171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5645 (.A(net1072),
    .X(net6172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5646 (.A(_04128_),
    .X(net6173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5647 (.A(net1073),
    .X(net6174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5648 (.A(\rbzero.spi_registers.new_texadd[3][23] ),
    .X(net6175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5649 (.A(net1386),
    .X(net6176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(net6121),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5650 (.A(_03839_),
    .X(net6177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5651 (.A(net1387),
    .X(net6178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5652 (.A(\rbzero.spi_registers.new_texadd[3][22] ),
    .X(net6179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5653 (.A(net1219),
    .X(net6180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5654 (.A(_03838_),
    .X(net6181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5655 (.A(net1220),
    .X(net6182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5656 (.A(\rbzero.tex_b1[16] ),
    .X(net6183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5657 (.A(net1069),
    .X(net6184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5658 (.A(_04371_),
    .X(net6185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5659 (.A(\rbzero.tex_r0[54] ),
    .X(net6186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(net6123),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5660 (.A(net1142),
    .X(net6187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5661 (.A(_04117_),
    .X(net6188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5662 (.A(net1143),
    .X(net6189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5663 (.A(\rbzero.spi_registers.new_texadd[2][20] ),
    .X(net6190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5664 (.A(net1343),
    .X(net6191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5665 (.A(_02504_),
    .X(net6192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5666 (.A(net1344),
    .X(net6193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5667 (.A(\rbzero.tex_r1[11] ),
    .X(net6194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5668 (.A(net1115),
    .X(net6195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5669 (.A(\rbzero.tex_g0[12] ),
    .X(net6196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(_01646_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5670 (.A(net1130),
    .X(net6197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5671 (.A(_04305_),
    .X(net6198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5672 (.A(net1131),
    .X(net6199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5673 (.A(\rbzero.pov.spi_buffer[53] ),
    .X(net6200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5674 (.A(net1110),
    .X(net6201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5675 (.A(\rbzero.tex_g1[48] ),
    .X(net6202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5676 (.A(net1127),
    .X(net6203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5677 (.A(_04195_),
    .X(net6204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5678 (.A(net1128),
    .X(net6205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5679 (.A(\rbzero.spi_registers.new_texadd[1][23] ),
    .X(net6206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(net6099),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5680 (.A(net1523),
    .X(net6207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5681 (.A(_03482_),
    .X(net6208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5682 (.A(net1524),
    .X(net6209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5683 (.A(\rbzero.tex_g1[14] ),
    .X(net6210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5684 (.A(net1173),
    .X(net6211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5685 (.A(_04232_),
    .X(net6212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5686 (.A(net1174),
    .X(net6213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5687 (.A(\rbzero.tex_b0[10] ),
    .X(net6214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5688 (.A(net1148),
    .X(net6215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5689 (.A(_04448_),
    .X(net6216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(net6101),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5690 (.A(net1149),
    .X(net6217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5691 (.A(\rbzero.tex_b1[36] ),
    .X(net6218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5692 (.A(net1185),
    .X(net6219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5693 (.A(_04349_),
    .X(net6220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5694 (.A(net1186),
    .X(net6221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5695 (.A(\rbzero.tex_g1[5] ),
    .X(net6222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5696 (.A(net1179),
    .X(net6223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5697 (.A(_04242_),
    .X(net6224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5698 (.A(net1180),
    .X(net6225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5699 (.A(\rbzero.tex_g1[58] ),
    .X(net6226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net5787),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_01656_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5700 (.A(net1188),
    .X(net6227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5701 (.A(_04183_),
    .X(net6228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5702 (.A(net1189),
    .X(net6229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5703 (.A(\rbzero.pov.spi_buffer[13] ),
    .X(net6230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5704 (.A(net1168),
    .X(net6231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5705 (.A(_03008_),
    .X(net6232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5706 (.A(net1169),
    .X(net6233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5707 (.A(\rbzero.tex_g0[38] ),
    .X(net6234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5708 (.A(net1139),
    .X(net6235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5709 (.A(_04277_),
    .X(net6236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(net6110),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5710 (.A(net1140),
    .X(net6237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5711 (.A(net6579),
    .X(net6238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5712 (.A(net1165),
    .X(net6239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5713 (.A(_03585_),
    .X(net6240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5714 (.A(net1166),
    .X(net6241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5715 (.A(\rbzero.tex_g1[46] ),
    .X(net6242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5716 (.A(net1191),
    .X(net6243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5717 (.A(_04197_),
    .X(net6244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5718 (.A(net1192),
    .X(net6245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5719 (.A(\rbzero.pov.spi_buffer[14] ),
    .X(net6246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(net6112),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5720 (.A(net1182),
    .X(net6247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5721 (.A(\rbzero.tex_b1[52] ),
    .X(net6248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5722 (.A(net1158),
    .X(net6249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5723 (.A(_04332_),
    .X(net6250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5724 (.A(net1159),
    .X(net6251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5725 (.A(\rbzero.spi_registers.new_texadd[0][2] ),
    .X(net6252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5726 (.A(net1211),
    .X(net6253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5727 (.A(_03433_),
    .X(net6254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5728 (.A(net1212),
    .X(net6255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5729 (.A(\rbzero.spi_registers.new_texadd[3][12] ),
    .X(net6256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(_01662_),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5730 (.A(net1200),
    .X(net6257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5731 (.A(\rbzero.tex_r1[35] ),
    .X(net6258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5732 (.A(net1235),
    .X(net6259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5733 (.A(_04063_),
    .X(net6260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5734 (.A(net1236),
    .X(net6261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5735 (.A(\rbzero.spi_registers.new_texadd[0][3] ),
    .X(net6262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5736 (.A(net1247),
    .X(net6263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5737 (.A(\rbzero.spi_registers.new_texadd[3][8] ),
    .X(net6264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5738 (.A(net1214),
    .X(net6265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5739 (.A(\rbzero.tex_b1[0] ),
    .X(net6266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(net7900),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5740 (.A(net1411),
    .X(net6267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5741 (.A(_04387_),
    .X(net6268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5742 (.A(net1412),
    .X(net6269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5743 (.A(\rbzero.tex_b1[12] ),
    .X(net6270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5744 (.A(net1225),
    .X(net6271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5745 (.A(_04376_),
    .X(net6272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5746 (.A(net1226),
    .X(net6273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5747 (.A(\rbzero.spi_registers.new_texadd[3][0] ),
    .X(net6274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5748 (.A(net1340),
    .X(net6275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5749 (.A(\rbzero.tex_r0[29] ),
    .X(net6276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(net2933),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5750 (.A(net1206),
    .X(net6277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5751 (.A(_04144_),
    .X(net6278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5752 (.A(net1207),
    .X(net6279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5753 (.A(\rbzero.spi_registers.new_texadd[0][8] ),
    .X(net6280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5754 (.A(net1278),
    .X(net6281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5755 (.A(\rbzero.spi_registers.new_texadd[3][6] ),
    .X(net6282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5756 (.A(net1263),
    .X(net6283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5757 (.A(\rbzero.spi_registers.new_texadd[0][1] ),
    .X(net6284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5758 (.A(net1377),
    .X(net6285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5759 (.A(\rbzero.spi_registers.new_mapd[9] ),
    .X(net6286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(net7482),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5760 (.A(net1292),
    .X(net6287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5761 (.A(_03413_),
    .X(net6288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5762 (.A(net1293),
    .X(net6289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5763 (.A(\rbzero.spi_registers.new_texadd[2][3] ),
    .X(net6290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5764 (.A(net1281),
    .X(net6291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5765 (.A(\rbzero.tex_g1[0] ),
    .X(net6292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5766 (.A(net1596),
    .X(net6293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5767 (.A(_04246_),
    .X(net6294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5768 (.A(net1597),
    .X(net6295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5769 (.A(\rbzero.spi_registers.new_texadd[0][6] ),
    .X(net6296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(_00685_),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5770 (.A(net1295),
    .X(net6297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5771 (.A(\rbzero.spi_registers.new_texadd[2][4] ),
    .X(net6298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5772 (.A(net1241),
    .X(net6299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5773 (.A(\rbzero.spi_registers.new_texadd[0][16] ),
    .X(net6300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5774 (.A(net1328),
    .X(net6301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5775 (.A(_03448_),
    .X(net6302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5776 (.A(net1329),
    .X(net6303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5777 (.A(\rbzero.spi_registers.new_texadd[0][0] ),
    .X(net6304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5778 (.A(net1301),
    .X(net6305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5779 (.A(\rbzero.spi_registers.new_texadd[2][10] ),
    .X(net6306));
 sky130_fd_sc_hd__buf_1 hold578 (.A(net7909),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5780 (.A(net1435),
    .X(net6307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5781 (.A(\rbzero.spi_registers.new_texadd[3][9] ),
    .X(net6308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5782 (.A(net1322),
    .X(net6309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5783 (.A(_03824_),
    .X(net6310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5784 (.A(net1323),
    .X(net6311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5785 (.A(\rbzero.spi_registers.new_texadd[1][1] ),
    .X(net6312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5786 (.A(net1310),
    .X(net6313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5787 (.A(\rbzero.spi_registers.new_texadd[0][10] ),
    .X(net6314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5788 (.A(net1468),
    .X(net6315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5789 (.A(\rbzero.spi_registers.new_texadd[3][18] ),
    .X(net6316));
 sky130_fd_sc_hd__buf_1 hold579 (.A(net8140),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5790 (.A(net1362),
    .X(net6317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5791 (.A(_03834_),
    .X(net6318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5792 (.A(net1363),
    .X(net6319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5793 (.A(\rbzero.spi_registers.new_texadd[0][23] ),
    .X(net6320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5794 (.A(net1266),
    .X(net6321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5795 (.A(_03455_),
    .X(net6322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5796 (.A(net1267),
    .X(net6323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5797 (.A(\rbzero.spi_registers.new_texadd[1][11] ),
    .X(net6324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5798 (.A(net1349),
    .X(net6325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5799 (.A(\rbzero.pov.spi_buffer[71] ),
    .X(net6326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net5789),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(net4281),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5800 (.A(net1260),
    .X(net6327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5801 (.A(_03596_),
    .X(net6328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5802 (.A(net1261),
    .X(net6329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5803 (.A(\rbzero.spi_registers.new_texadd[2][23] ),
    .X(net6330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5804 (.A(net1389),
    .X(net6331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5805 (.A(_02507_),
    .X(net6332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5806 (.A(net1390),
    .X(net6333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5807 (.A(\rbzero.spi_registers.new_texadd[2][2] ),
    .X(net6334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5808 (.A(net1422),
    .X(net6335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5809 (.A(_02482_),
    .X(net6336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(net5475),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5810 (.A(net1423),
    .X(net6337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5811 (.A(\rbzero.spi_registers.new_texadd[2][14] ),
    .X(net6338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5812 (.A(net1380),
    .X(net6339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5813 (.A(\rbzero.spi_registers.new_texadd[1][2] ),
    .X(net6340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5814 (.A(net1337),
    .X(net6341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5815 (.A(_03460_),
    .X(net6342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5816 (.A(net1338),
    .X(net6343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5817 (.A(\rbzero.tex_b1[62] ),
    .X(net6344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5818 (.A(net1298),
    .X(net6345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5819 (.A(\rbzero.spi_registers.new_texadd[1][16] ),
    .X(net6346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(net5477),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5820 (.A(net1325),
    .X(net6347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5821 (.A(_03475_),
    .X(net6348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5822 (.A(net1326),
    .X(net6349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5823 (.A(\rbzero.spi_registers.new_texadd[1][9] ),
    .X(net6350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5824 (.A(net1511),
    .X(net6351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5825 (.A(_03467_),
    .X(net6352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5826 (.A(net1512),
    .X(net6353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5827 (.A(\rbzero.spi_registers.new_texadd[2][0] ),
    .X(net6354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5828 (.A(net1286),
    .X(net6355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5829 (.A(\rbzero.pov.spi_buffer[26] ),
    .X(net6356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net6200),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5830 (.A(net1230),
    .X(net6357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5831 (.A(\rbzero.tex_r0[0] ),
    .X(net6358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5832 (.A(net1794),
    .X(net6359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5833 (.A(_04175_),
    .X(net6360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5834 (.A(net1795),
    .X(net6361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5835 (.A(\rbzero.spi_registers.new_texadd[2][9] ),
    .X(net6362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5836 (.A(net1514),
    .X(net6363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5837 (.A(_02492_),
    .X(net6364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5838 (.A(net1515),
    .X(net6365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5839 (.A(\rbzero.spi_registers.new_texadd[0][5] ),
    .X(net6366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_03577_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5840 (.A(net1374),
    .X(net6367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5841 (.A(_03436_),
    .X(net6368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5842 (.A(\rbzero.spi_registers.new_texadd[1][12] ),
    .X(net6369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5843 (.A(net1453),
    .X(net6370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5844 (.A(\rbzero.spi_registers.new_texadd[3][14] ),
    .X(net6371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5845 (.A(net1355),
    .X(net6372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5846 (.A(\rbzero.spi_registers.new_texadd[3][2] ),
    .X(net6373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5847 (.A(net1368),
    .X(net6374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5848 (.A(_03817_),
    .X(net6375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5849 (.A(net1369),
    .X(net6376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(_01140_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5850 (.A(\rbzero.spi_registers.new_texadd[3][7] ),
    .X(net6377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5851 (.A(net1441),
    .X(net6378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5852 (.A(\rbzero.spi_registers.new_texadd[2][15] ),
    .X(net6379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5853 (.A(net1444),
    .X(net6380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5854 (.A(_02499_),
    .X(net6381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5855 (.A(net1445),
    .X(net6382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5856 (.A(\rbzero.spi_registers.new_texadd[2][16] ),
    .X(net6383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5857 (.A(net1371),
    .X(net6384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5858 (.A(_02500_),
    .X(net6385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5859 (.A(net1372),
    .X(net6386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(net7592),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5860 (.A(\rbzero.spi_registers.new_texadd[0][13] ),
    .X(net6387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5861 (.A(net1405),
    .X(net6388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5862 (.A(\rbzero.spi_registers.new_texadd[2][5] ),
    .X(net6389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5863 (.A(net1419),
    .X(net6390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5864 (.A(_02488_),
    .X(net6391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5865 (.A(\rbzero.spi_registers.new_texadd[2][1] ),
    .X(net6392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5866 (.A(net597),
    .X(net6393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5867 (.A(\rbzero.spi_registers.new_mapd[2] ),
    .X(net6394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5868 (.A(net1319),
    .X(net6395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5869 (.A(_03406_),
    .X(net6396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(net4474),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5870 (.A(net1320),
    .X(net6397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5871 (.A(\rbzero.spi_registers.new_texadd[1][8] ),
    .X(net6398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5872 (.A(net1552),
    .X(net6399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5873 (.A(\rbzero.spi_registers.new_texadd[0][20] ),
    .X(net6400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5874 (.A(net1331),
    .X(net6401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5875 (.A(_03452_),
    .X(net6402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5876 (.A(net1332),
    .X(net6403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5877 (.A(\rbzero.spi_registers.new_texadd[2][8] ),
    .X(net6404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5878 (.A(net1508),
    .X(net6405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5879 (.A(\rbzero.spi_registers.new_texadd[2][12] ),
    .X(net6406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(net6194),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5880 (.A(net1456),
    .X(net6407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5881 (.A(\rbzero.spi_registers.new_texadd[3][3] ),
    .X(net6408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5882 (.A(net1304),
    .X(net6409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5883 (.A(\rbzero.spi_registers.new_mapd[0] ),
    .X(net6410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5884 (.A(net1429),
    .X(net6411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5885 (.A(\rbzero.pov.spi_buffer[4] ),
    .X(net6412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5886 (.A(net1316),
    .X(net6413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5887 (.A(_03523_),
    .X(net6414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5888 (.A(net1317),
    .X(net6415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5889 (.A(\rbzero.spi_registers.new_texadd[1][10] ),
    .X(net6416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_04090_),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5890 (.A(net1489),
    .X(net6417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5891 (.A(\rbzero.spi_registers.new_texadd[1][5] ),
    .X(net6418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5892 (.A(net1416),
    .X(net6419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5893 (.A(_03463_),
    .X(net6420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5894 (.A(\rbzero.spi_registers.new_texadd[1][15] ),
    .X(net6421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5895 (.A(net1496),
    .X(net6422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5896 (.A(_03474_),
    .X(net6423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5897 (.A(net1497),
    .X(net6424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5898 (.A(\rbzero.spi_registers.new_texadd[2][19] ),
    .X(net6425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5899 (.A(net839),
    .X(net6426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_01573_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_01544_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5900 (.A(_02503_),
    .X(net6427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5901 (.A(net1448),
    .X(net6428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5902 (.A(net8276),
    .X(net6429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5903 (.A(net1432),
    .X(net6430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5904 (.A(_03454_),
    .X(net6431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5905 (.A(net1433),
    .X(net6432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5906 (.A(\rbzero.spi_registers.new_texadd[0][12] ),
    .X(net6433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5907 (.A(net1483),
    .X(net6434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5908 (.A(\rbzero.pov.spi_buffer[33] ),
    .X(net6435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5909 (.A(net1244),
    .X(net6436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net5455),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5910 (.A(_03030_),
    .X(net6437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5911 (.A(net1245),
    .X(net6438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5912 (.A(\rbzero.spi_registers.new_texadd[1][4] ),
    .X(net6439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5913 (.A(net1346),
    .X(net6440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5914 (.A(\rbzero.tex_b1[44] ),
    .X(net6441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5915 (.A(net1352),
    .X(net6442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5916 (.A(_04340_),
    .X(net6443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5917 (.A(net1353),
    .X(net6444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5918 (.A(\rbzero.spi_registers.new_texadd[3][10] ),
    .X(net6445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5919 (.A(net1474),
    .X(net6446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(net5457),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5920 (.A(\rbzero.spi_registers.new_texadd[0][4] ),
    .X(net6447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5921 (.A(net1544),
    .X(net6448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5922 (.A(\rbzero.spi_registers.new_texadd[3][5] ),
    .X(net6449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5923 (.A(net1465),
    .X(net6450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5924 (.A(_03820_),
    .X(net6451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5925 (.A(net1466),
    .X(net6452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5926 (.A(\rbzero.spi_registers.new_texadd[2][7] ),
    .X(net6453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5927 (.A(net1631),
    .X(net6454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5928 (.A(\rbzero.tex_g1[33] ),
    .X(net6455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5929 (.A(net1313),
    .X(net6456));
 sky130_fd_sc_hd__buf_1 hold593 (.A(net8137),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5930 (.A(_04211_),
    .X(net6457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5931 (.A(net1314),
    .X(net6458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5932 (.A(\rbzero.tex_b0[46] ),
    .X(net6459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5933 (.A(net1197),
    .X(net6460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5934 (.A(_04408_),
    .X(net6461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5935 (.A(net1198),
    .X(net6462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5936 (.A(\rbzero.spi_registers.new_mapd[11] ),
    .X(net6463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5937 (.A(net1176),
    .X(net6464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5938 (.A(\rbzero.tex_g1[50] ),
    .X(net6465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5939 (.A(net1450),
    .X(net6466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(net4237),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5940 (.A(_04191_),
    .X(net6467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5941 (.A(net1451),
    .X(net6468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5942 (.A(\rbzero.spi_registers.new_texadd[3][13] ),
    .X(net6469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5943 (.A(net1502),
    .X(net6470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5944 (.A(\rbzero.spi_registers.new_texadd[1][14] ),
    .X(net6471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5945 (.A(net986),
    .X(net6472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5946 (.A(\rbzero.spi_registers.new_texadd[1][0] ),
    .X(net6473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5947 (.A(net1307),
    .X(net6474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5948 (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .X(net6475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5949 (.A(net1492),
    .X(net6476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(net5451),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5950 (.A(\rbzero.tex_g1[18] ),
    .X(net6477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5951 (.A(net1257),
    .X(net6478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5952 (.A(_04228_),
    .X(net6479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5953 (.A(net1258),
    .X(net6480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5954 (.A(\rbzero.spi_registers.new_mapd[10] ),
    .X(net6481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5955 (.A(net1289),
    .X(net6482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5956 (.A(\rbzero.spi_registers.new_texadd[1][13] ),
    .X(net6483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5957 (.A(net1462),
    .X(net6484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5958 (.A(\rbzero.spi_registers.new_other[3] ),
    .X(net6485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5959 (.A(net1076),
    .X(net6486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(net5453),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5960 (.A(\rbzero.tex_r0[19] ),
    .X(net6487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5961 (.A(net1520),
    .X(net6488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5962 (.A(_04155_),
    .X(net6489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5963 (.A(net1521),
    .X(net6490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5964 (.A(\rbzero.spi_registers.new_texadd[2][6] ),
    .X(net6491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5965 (.A(net1538),
    .X(net6492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5966 (.A(\rbzero.spi_registers.new_other[2] ),
    .X(net6493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5967 (.A(net1061),
    .X(net6494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5968 (.A(\rbzero.spi_registers.new_texadd[3][16] ),
    .X(net6495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5969 (.A(net1576),
    .X(net6496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(net5687),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5970 (.A(_03832_),
    .X(net6497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5971 (.A(net1577),
    .X(net6498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5972 (.A(\rbzero.tex_g0[10] ),
    .X(net6499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5973 (.A(net1272),
    .X(net6500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5974 (.A(_04307_),
    .X(net6501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5975 (.A(net1273),
    .X(net6502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5976 (.A(\rbzero.spi_registers.new_texadd[1][3] ),
    .X(net6503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5977 (.A(net1694),
    .X(net6504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5978 (.A(\rbzero.tex_g0[18] ),
    .X(net6505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5979 (.A(net1269),
    .X(net6506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(net5689),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5980 (.A(_04299_),
    .X(net6507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5981 (.A(net1270),
    .X(net6508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5982 (.A(\rbzero.spi_registers.new_texadd[3][4] ),
    .X(net6509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5983 (.A(net1459),
    .X(net6510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5984 (.A(\rbzero.pov.spi_buffer[23] ),
    .X(net6511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5985 (.A(net1222),
    .X(net6512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5986 (.A(_03019_),
    .X(net6513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5987 (.A(net1223),
    .X(net6514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5988 (.A(\rbzero.spi_registers.new_texadd[0][19] ),
    .X(net6515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5989 (.A(net1570),
    .X(net6516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(_01480_),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5990 (.A(_03451_),
    .X(net6517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5991 (.A(net1571),
    .X(net6518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5992 (.A(\rbzero.spi_registers.new_texadd[0][15] ),
    .X(net6519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5993 (.A(net1811),
    .X(net6520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5994 (.A(_03447_),
    .X(net6521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5995 (.A(net1812),
    .X(net6522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5996 (.A(\rbzero.tex_b1[35] ),
    .X(net6523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5997 (.A(net1408),
    .X(net6524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5998 (.A(_04350_),
    .X(net6525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5999 (.A(net1409),
    .X(net6526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net5987),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(net6202),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6000 (.A(\rbzero.spi_registers.new_texadd[2][18] ),
    .X(net6527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6001 (.A(net1602),
    .X(net6528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6002 (.A(_02502_),
    .X(net6529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6003 (.A(net1603),
    .X(net6530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6004 (.A(\rbzero.spi_registers.new_texadd[1][7] ),
    .X(net6531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6005 (.A(net1800),
    .X(net6532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6006 (.A(\rbzero.tex_b0[55] ),
    .X(net6533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6007 (.A(net1499),
    .X(net6534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6008 (.A(_04398_),
    .X(net6535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6009 (.A(net1500),
    .X(net6536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(net6204),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6010 (.A(\rbzero.tex_b0[34] ),
    .X(net6537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6011 (.A(net1712),
    .X(net6538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6012 (.A(_04421_),
    .X(net6539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6013 (.A(net1713),
    .X(net6540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6014 (.A(\rbzero.spi_registers.new_texadd[0][7] ),
    .X(net6541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6015 (.A(net1668),
    .X(net6542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6016 (.A(\rbzero.spi_registers.new_vshift[4] ),
    .X(net6543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6017 (.A(net1742),
    .X(net6544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6018 (.A(\rbzero.spi_registers.new_leak[1] ),
    .X(net6545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6019 (.A(net1643),
    .X(net6546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_01453_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6020 (.A(\rbzero.tex_b1[56] ),
    .X(net6547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6021 (.A(net1526),
    .X(net6548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6022 (.A(_04327_),
    .X(net6549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6023 (.A(net1527),
    .X(net6550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6024 (.A(\rbzero.spi_registers.new_texadd[3][1] ),
    .X(net6551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6025 (.A(net1555),
    .X(net6552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6026 (.A(\rbzero.tex_r1[4] ),
    .X(net6553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6027 (.A(net1383),
    .X(net6554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6028 (.A(_04098_),
    .X(net6555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6029 (.A(net1384),
    .X(net6556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(net6196),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6030 (.A(\rbzero.spi_registers.new_texadd[2][11] ),
    .X(net6557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6031 (.A(net1859),
    .X(net6558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6032 (.A(\rbzero.pov.ready_buffer[4] ),
    .X(net6559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6033 (.A(net1573),
    .X(net6560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6034 (.A(\rbzero.spi_registers.new_texadd[1][19] ),
    .X(net6561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6035 (.A(net1665),
    .X(net6562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6036 (.A(_03478_),
    .X(net6563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6037 (.A(net1666),
    .X(net6564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6038 (.A(\rbzero.spi_registers.new_texadd[0][9] ),
    .X(net6565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6039 (.A(net1628),
    .X(net6566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(net6198),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6040 (.A(_03440_),
    .X(net6567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6041 (.A(net1629),
    .X(net6568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6042 (.A(\rbzero.spi_registers.new_texadd[3][15] ),
    .X(net6569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6043 (.A(net1685),
    .X(net6570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6044 (.A(_03831_),
    .X(net6571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6045 (.A(net1686),
    .X(net6572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6046 (.A(\rbzero.spi_registers.new_mapd[15] ),
    .X(net6573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6047 (.A(net1637),
    .X(net6574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6048 (.A(_03419_),
    .X(net6575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6049 (.A(net1638),
    .X(net6576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_01353_),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6050 (.A(\rbzero.spi_registers.new_leak[4] ),
    .X(net6577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6051 (.A(net1671),
    .X(net6578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6052 (.A(\rbzero.pov.spi_buffer[60] ),
    .X(net6579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6053 (.A(\rbzero.tex_r1[60] ),
    .X(net6580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6054 (.A(net1605),
    .X(net6581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6055 (.A(_04036_),
    .X(net6582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6056 (.A(net1606),
    .X(net6583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6057 (.A(\rbzero.spi_registers.new_texadd[2][13] ),
    .X(net6584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6058 (.A(net1677),
    .X(net6585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6059 (.A(\rbzero.tex_g0[62] ),
    .X(net6586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net6857),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6060 (.A(net1587),
    .X(net6587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6061 (.A(_04249_),
    .X(net6588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6062 (.A(net1588),
    .X(net6589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6063 (.A(\rbzero.tex_g0[19] ),
    .X(net6590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6064 (.A(net1739),
    .X(net6591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6065 (.A(\rbzero.tex_g0[57] ),
    .X(net6592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6066 (.A(net1805),
    .X(net6593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6067 (.A(_04255_),
    .X(net6594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6068 (.A(net1806),
    .X(net6595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6069 (.A(\rbzero.spi_registers.new_mapd[12] ),
    .X(net6596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_03153_),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6070 (.A(net1203),
    .X(net6597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6071 (.A(\rbzero.spi_registers.new_texadd[1][6] ),
    .X(net6598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6072 (.A(net1691),
    .X(net6599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6073 (.A(\rbzero.spi_registers.new_texadd[3][11] ),
    .X(net6600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6074 (.A(net1785),
    .X(net6601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6075 (.A(\rbzero.spi_registers.new_texadd[2][17] ),
    .X(net6602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6076 (.A(net1718),
    .X(net6603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6077 (.A(_02501_),
    .X(net6604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6078 (.A(net1719),
    .X(net6605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6079 (.A(\rbzero.tex_r1[7] ),
    .X(net6606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(net5506),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6080 (.A(net1755),
    .X(net6607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6081 (.A(_04094_),
    .X(net6608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6082 (.A(net1756),
    .X(net6609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6083 (.A(\rbzero.spi_registers.mosi_buffer[0] ),
    .X(net6610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6084 (.A(net1727),
    .X(net6611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6085 (.A(\rbzero.spi_registers.new_vshift[0] ),
    .X(net6612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6086 (.A(net1033),
    .X(net6613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6087 (.A(\rbzero.tex_g1[55] ),
    .X(net6614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6088 (.A(net1486),
    .X(net6615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6089 (.A(_04186_),
    .X(net6616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(net5459),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6090 (.A(net1487),
    .X(net6617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6091 (.A(\rbzero.spi_registers.new_texadd[0][21] ),
    .X(net6618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6092 (.A(net1649),
    .X(net6619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6093 (.A(_03453_),
    .X(net6620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6094 (.A(net1650),
    .X(net6621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6095 (.A(\rbzero.spi_registers.new_texadd[1][17] ),
    .X(net6622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6096 (.A(net1697),
    .X(net6623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6097 (.A(_03476_),
    .X(net6624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6098 (.A(net1698),
    .X(net6625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6099 (.A(\gpout3.clk_div[1] ),
    .X(net6626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net5989),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(net5461),
    .X(net1137));
 sky130_fd_sc_hd__buf_1 hold6100 (.A(net2613),
    .X(net6627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6101 (.A(\rbzero.spi_registers.new_texadd[1][18] ),
    .X(net6628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6102 (.A(net1745),
    .X(net6629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6103 (.A(_03477_),
    .X(net6630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6104 (.A(net1746),
    .X(net6631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6105 (.A(\rbzero.tex_g0[5] ),
    .X(net6632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6106 (.A(net1891),
    .X(net6633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6107 (.A(_04313_),
    .X(net6634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6108 (.A(net1892),
    .X(net6635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6109 (.A(\rbzero.tex_b1[9] ),
    .X(net6636));
 sky130_fd_sc_hd__buf_1 hold611 (.A(net7855),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6110 (.A(net1827),
    .X(net6637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6111 (.A(_04379_),
    .X(net6638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6112 (.A(net1828),
    .X(net6639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6113 (.A(\rbzero.tex_g0[11] ),
    .X(net6640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6114 (.A(net1715),
    .X(net6641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6115 (.A(\rbzero.tex_g1[25] ),
    .X(net6642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6116 (.A(net1652),
    .X(net6643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6117 (.A(_04220_),
    .X(net6644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6118 (.A(net1653),
    .X(net6645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6119 (.A(\rbzero.spi_registers.new_texadd[0][11] ),
    .X(net6646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(net6234),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6120 (.A(net1923),
    .X(net6647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6121 (.A(\rbzero.pov.spi_buffer[25] ),
    .X(net6648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6122 (.A(net1688),
    .X(net6649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6123 (.A(\rbzero.tex_r0[33] ),
    .X(net6650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6124 (.A(net1833),
    .X(net6651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6125 (.A(_04140_),
    .X(net6652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6126 (.A(net1834),
    .X(net6653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6127 (.A(\rbzero.tex_g0[6] ),
    .X(net6654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6128 (.A(net1973),
    .X(net6655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6129 (.A(\rbzero.tex_b1[25] ),
    .X(net6656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(net6236),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6130 (.A(net1797),
    .X(net6657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6131 (.A(_04361_),
    .X(net6658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6132 (.A(net1798),
    .X(net6659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6133 (.A(\rbzero.pov.spi_buffer[5] ),
    .X(net6660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6134 (.A(net1579),
    .X(net6661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6135 (.A(_03524_),
    .X(net6662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6136 (.A(net1580),
    .X(net6663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6137 (.A(\rbzero.pov.spi_buffer[73] ),
    .X(net6664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6138 (.A(net1613),
    .X(net6665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6139 (.A(_03597_),
    .X(net6666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_01379_),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6140 (.A(net1870),
    .X(net6667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6141 (.A(\rbzero.tex_r0[42] ),
    .X(net6668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6142 (.A(net1848),
    .X(net6669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6143 (.A(_04130_),
    .X(net6670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6144 (.A(net1849),
    .X(net6671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6145 (.A(\rbzero.tex_b0[25] ),
    .X(net6672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6146 (.A(net1730),
    .X(net6673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6147 (.A(_04431_),
    .X(net6674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6148 (.A(net1731),
    .X(net6675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6149 (.A(\rbzero.spi_registers.new_texadd[3][17] ),
    .X(net6676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(net6186),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6150 (.A(net1767),
    .X(net6677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6151 (.A(_03833_),
    .X(net6678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6152 (.A(net1768),
    .X(net6679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6153 (.A(\rbzero.pov.ready_buffer[3] ),
    .X(net6680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6154 (.A(net1862),
    .X(net6681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6155 (.A(\rbzero.spi_registers.new_texadd[3][19] ),
    .X(net6682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6156 (.A(net2220),
    .X(net6683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6157 (.A(_03835_),
    .X(net6684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6158 (.A(net2221),
    .X(net6685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6159 (.A(\rbzero.pov.ready_buffer[54] ),
    .X(net6686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(net6188),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6160 (.A(net616),
    .X(net6687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6161 (.A(\rbzero.tex_r1[55] ),
    .X(net6688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6162 (.A(net2119),
    .X(net6689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6163 (.A(_04041_),
    .X(net6690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6164 (.A(net2120),
    .X(net6691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6165 (.A(\rbzero.pov.ready_buffer[6] ),
    .X(net6692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6166 (.A(net746),
    .X(net6693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6167 (.A(_03000_),
    .X(net6694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6168 (.A(net1683),
    .X(net6695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6169 (.A(\rbzero.spi_registers.new_texadd[0][14] ),
    .X(net6696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(_01523_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6170 (.A(net1770),
    .X(net6697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6171 (.A(\rbzero.tex_b1[24] ),
    .X(net6698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6172 (.A(net1660),
    .X(net6699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6173 (.A(_04362_),
    .X(net6700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6174 (.A(net1661),
    .X(net6701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6175 (.A(\rbzero.tex_r0[25] ),
    .X(net6702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6176 (.A(net2091),
    .X(net6703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6177 (.A(\rbzero.tex_g0[13] ),
    .X(net6704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6178 (.A(net1872),
    .X(net6705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6179 (.A(\rbzero.pov.ready_buffer[18] ),
    .X(net6706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(net2800),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6180 (.A(net1875),
    .X(net6707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6181 (.A(_03013_),
    .X(net6708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6182 (.A(net1876),
    .X(net6709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6183 (.A(\rbzero.tex_g0[21] ),
    .X(net6710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6184 (.A(net2110),
    .X(net6711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6185 (.A(_04295_),
    .X(net6712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6186 (.A(net2111),
    .X(net6713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6187 (.A(\rbzero.tex_r1[19] ),
    .X(net6714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6188 (.A(net1839),
    .X(net6715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6189 (.A(_04081_),
    .X(net6716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(_03046_),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6190 (.A(net1840),
    .X(net6717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6191 (.A(\rbzero.tex_g1[37] ),
    .X(net6718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6192 (.A(net2429),
    .X(net6719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6193 (.A(_04207_),
    .X(net6720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6194 (.A(net2430),
    .X(net6721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6195 (.A(\rbzero.tex_g0[26] ),
    .X(net6722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6196 (.A(net1782),
    .X(net6723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6197 (.A(_04290_),
    .X(net6724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6198 (.A(net1783),
    .X(net6725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6199 (.A(\rbzero.spi_registers.new_texadd[0][18] ),
    .X(net6726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_01155_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_00695_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6200 (.A(net1903),
    .X(net6727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6201 (.A(_03450_),
    .X(net6728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6202 (.A(net1904),
    .X(net6729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6203 (.A(\rbzero.pov.spi_buffer[37] ),
    .X(net6730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6204 (.A(net1618),
    .X(net6731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6205 (.A(_03034_),
    .X(net6732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6206 (.A(net1619),
    .X(net6733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6207 (.A(\rbzero.tex_r0[35] ),
    .X(net6734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6208 (.A(net1853),
    .X(net6735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6209 (.A(_04137_),
    .X(net6736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(net6214),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6210 (.A(net1854),
    .X(net6737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6211 (.A(\rbzero.spi_registers.new_leak[5] ),
    .X(net6738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6212 (.A(net2146),
    .X(net6739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6213 (.A(_03371_),
    .X(net6740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6214 (.A(\rbzero.spi_registers.new_mapd[13] ),
    .X(net6741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6215 (.A(net1238),
    .X(net6742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6216 (.A(\rbzero.pov.spi_buffer[47] ),
    .X(net6743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6217 (.A(net1885),
    .X(net6744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6218 (.A(\rbzero.tex_b0[58] ),
    .X(net6745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6219 (.A(net1761),
    .X(net6746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(net6216),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6220 (.A(_04395_),
    .X(net6747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6221 (.A(net1762),
    .X(net6748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6222 (.A(\rbzero.tex_g1[15] ),
    .X(net6749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6223 (.A(net2029),
    .X(net6750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6224 (.A(\rbzero.tex_r1[21] ),
    .X(net6751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6225 (.A(net1912),
    .X(net6752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6226 (.A(\rbzero.tex_r1[22] ),
    .X(net6753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6227 (.A(net1991),
    .X(net6754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6228 (.A(\rbzero.tex_g0[53] ),
    .X(net6755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6229 (.A(net2052),
    .X(net6756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(_01031_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6230 (.A(\rbzero.tex_r1[54] ),
    .X(net6757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6231 (.A(net2131),
    .X(net6758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6232 (.A(_04043_),
    .X(net6759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6233 (.A(net2132),
    .X(net6760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6234 (.A(\rbzero.tex_g0[39] ),
    .X(net6761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6235 (.A(net1900),
    .X(net6762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6236 (.A(\rbzero.tex_b1[45] ),
    .X(net6763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6237 (.A(net2000),
    .X(net6764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6238 (.A(\rbzero.tex_b1[34] ),
    .X(net6765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6239 (.A(net1955),
    .X(net6766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(net3319),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6240 (.A(\rbzero.tex_b0[17] ),
    .X(net6767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6241 (.A(net1952),
    .X(net6768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6242 (.A(_04440_),
    .X(net6769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6243 (.A(net1953),
    .X(net6770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6244 (.A(\rbzero.tex_g1[49] ),
    .X(net6771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6245 (.A(net2008),
    .X(net6772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6246 (.A(\rbzero.tex_g1[16] ),
    .X(net6773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6247 (.A(net2085),
    .X(net6774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6248 (.A(\rbzero.tex_g0[17] ),
    .X(net6775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6249 (.A(net1920),
    .X(net6776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_03560_),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6250 (.A(_04300_),
    .X(net6777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6251 (.A(net1921),
    .X(net6778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6252 (.A(\rbzero.tex_b0[15] ),
    .X(net6779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6253 (.A(net1721),
    .X(net6780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6254 (.A(_04442_),
    .X(net6781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6255 (.A(net1722),
    .X(net6782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6256 (.A(\rbzero.tex_g1[27] ),
    .X(net6783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6257 (.A(net1985),
    .X(net6784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6258 (.A(_04218_),
    .X(net6785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6259 (.A(net1986),
    .X(net6786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_01125_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6260 (.A(\rbzero.tex_b0[45] ),
    .X(net6787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6261 (.A(net1982),
    .X(net6788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6262 (.A(_04409_),
    .X(net6789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6263 (.A(net1983),
    .X(net6790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6264 (.A(\rbzero.spi_registers.sclk_buffer[0] ),
    .X(net6791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6265 (.A(net2055),
    .X(net6792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6266 (.A(_03115_),
    .X(net6793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6267 (.A(net2183),
    .X(net6794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6268 (.A(\rbzero.tex_g1[59] ),
    .X(net6795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6269 (.A(net1994),
    .X(net6796));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold627 (.A(net4611),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6270 (.A(_04180_),
    .X(net6797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6271 (.A(net2050),
    .X(net6798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6272 (.A(\rbzero.spi_registers.new_mapd[1] ),
    .X(net6799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6273 (.A(net1997),
    .X(net6800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6274 (.A(\rbzero.tex_b0[21] ),
    .X(net6801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6275 (.A(net1824),
    .X(net6802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6276 (.A(\rbzero.tex_b0[57] ),
    .X(net6803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6277 (.A(net1819),
    .X(net6804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6278 (.A(_04396_),
    .X(net6805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6279 (.A(net1820),
    .X(net6806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(net4260),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6280 (.A(\rbzero.tex_g1[20] ),
    .X(net6807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6281 (.A(net1961),
    .X(net6808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6282 (.A(_04225_),
    .X(net6809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6283 (.A(net1962),
    .X(net6810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6284 (.A(\rbzero.tex_g1[41] ),
    .X(net6811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6285 (.A(net1935),
    .X(net6812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6286 (.A(_04202_),
    .X(net6813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6287 (.A(net1936),
    .X(net6814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6288 (.A(\rbzero.spi_registers.new_vinf ),
    .X(net6815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6289 (.A(net636),
    .X(net6816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(net5463),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6290 (.A(\rbzero.tex_g1[61] ),
    .X(net6817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6291 (.A(net2226),
    .X(net6818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6292 (.A(_04179_),
    .X(net6819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6293 (.A(net2227),
    .X(net6820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6294 (.A(\rbzero.tex_r0[39] ),
    .X(net6821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6295 (.A(net2101),
    .X(net6822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6296 (.A(_04133_),
    .X(net6823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6297 (.A(net2102),
    .X(net6824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6298 (.A(\rbzero.tex_r0[38] ),
    .X(net6825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6299 (.A(net1517),
    .X(net6826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net5990),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(net5465),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6300 (.A(_04134_),
    .X(net6827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6301 (.A(net1518),
    .X(net6828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6302 (.A(\rbzero.tex_b0[29] ),
    .X(net6829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6303 (.A(net1897),
    .X(net6830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6304 (.A(_04427_),
    .X(net6831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6305 (.A(net1898),
    .X(net6832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6306 (.A(\rbzero.tex_r0[12] ),
    .X(net6833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6307 (.A(net1926),
    .X(net6834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6308 (.A(\rbzero.tex_r1[57] ),
    .X(net6835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6309 (.A(net1976),
    .X(net6836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(net6248),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6310 (.A(_04039_),
    .X(net6837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6311 (.A(net1977),
    .X(net6838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6312 (.A(\rbzero.tex_r0[27] ),
    .X(net6839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6313 (.A(net1845),
    .X(net6840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6314 (.A(_04146_),
    .X(net6841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6315 (.A(net1846),
    .X(net6842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6316 (.A(\rbzero.spi_registers.new_leak[2] ),
    .X(net6843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6317 (.A(net2256),
    .X(net6844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6318 (.A(\rbzero.tex_b1[21] ),
    .X(net6845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6319 (.A(net2107),
    .X(net6846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(net6250),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6320 (.A(_04366_),
    .X(net6847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6321 (.A(net2108),
    .X(net6848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6322 (.A(\rbzero.tex_b0[24] ),
    .X(net6849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6323 (.A(net1758),
    .X(net6850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6324 (.A(_04432_),
    .X(net6851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6325 (.A(net1759),
    .X(net6852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6326 (.A(\rbzero.tex_g0[36] ),
    .X(net6853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6327 (.A(net2563),
    .X(net6854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6328 (.A(_04279_),
    .X(net6855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6329 (.A(net2564),
    .X(net6856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_01329_),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6330 (.A(\rbzero.spi_registers.new_mapd[14] ),
    .X(net6857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6331 (.A(net1133),
    .X(net6858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6332 (.A(\rbzero.tex_r0[28] ),
    .X(net6859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6333 (.A(net2140),
    .X(net6860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6334 (.A(\rbzero.spi_registers.new_texadd[0][17] ),
    .X(net6861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6335 (.A(net2268),
    .X(net6862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6336 (.A(_03449_),
    .X(net6863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6337 (.A(net2269),
    .X(net6864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6338 (.A(\rbzero.tex_b1[30] ),
    .X(net6865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6339 (.A(net1888),
    .X(net6866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(net5471),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6340 (.A(\rbzero.tex_b0[13] ),
    .X(net6867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6341 (.A(net1909),
    .X(net6868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6342 (.A(_04444_),
    .X(net6869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6343 (.A(net1910),
    .X(net6870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6344 (.A(\rbzero.tex_r1[17] ),
    .X(net6871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6345 (.A(net2020),
    .X(net6872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6346 (.A(\rbzero.tex_g0[4] ),
    .X(net6873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6347 (.A(net2116),
    .X(net6874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6348 (.A(_04314_),
    .X(net6875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6349 (.A(net2117),
    .X(net6876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(net5473),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6350 (.A(\rbzero.pov.ready_buffer[39] ),
    .X(net6877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6351 (.A(net1932),
    .X(net6878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6352 (.A(\rbzero.tex_r1[46] ),
    .X(net6879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6353 (.A(net2128),
    .X(net6880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6354 (.A(_04051_),
    .X(net6881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6355 (.A(net2129),
    .X(net6882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6356 (.A(\rbzero.tex_g0[50] ),
    .X(net6883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6357 (.A(net2014),
    .X(net6884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6358 (.A(_04262_),
    .X(net6885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6359 (.A(net2015),
    .X(net6886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(net5467),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6360 (.A(\rbzero.tex_r1[58] ),
    .X(net6887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6361 (.A(net2297),
    .X(net6888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6362 (.A(\rbzero.tex_b1[7] ),
    .X(net6889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6363 (.A(net2536),
    .X(net6890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6364 (.A(_04380_),
    .X(net6891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6365 (.A(net2579),
    .X(net6892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6366 (.A(\rbzero.tex_b1[51] ),
    .X(net6893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6367 (.A(net2063),
    .X(net6894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6368 (.A(_04333_),
    .X(net6895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6369 (.A(net2064),
    .X(net6896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(net5469),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6370 (.A(\rbzero.tex_r1[6] ),
    .X(net6897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6371 (.A(net2336),
    .X(net6898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6372 (.A(_04095_),
    .X(net6899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6373 (.A(net2337),
    .X(net6900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6374 (.A(\rbzero.tex_r1[59] ),
    .X(net6901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6375 (.A(net2348),
    .X(net6902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6376 (.A(\rbzero.tex_b0[63] ),
    .X(net6903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6377 (.A(net1967),
    .X(net6904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6378 (.A(\rbzero.tex_r0[58] ),
    .X(net6905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6379 (.A(net2158),
    .X(net6906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(net6238),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6380 (.A(_04112_),
    .X(net6907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6381 (.A(net2159),
    .X(net6908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6382 (.A(\rbzero.tex_g1[56] ),
    .X(net6909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6383 (.A(net2700),
    .X(net6910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6384 (.A(_04184_),
    .X(net6911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6385 (.A(net2245),
    .X(net6912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6386 (.A(\rbzero.tex_r0[41] ),
    .X(net6913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6387 (.A(net2423),
    .X(net6914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6388 (.A(_04131_),
    .X(net6915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6389 (.A(net2424),
    .X(net6916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(net6240),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6390 (.A(\rbzero.tex_r0[32] ),
    .X(net6917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6391 (.A(net2405),
    .X(net6918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6392 (.A(_04141_),
    .X(net6919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6393 (.A(net2406),
    .X(net6920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6394 (.A(\rbzero.tex_r1[12] ),
    .X(net6921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6395 (.A(net2271),
    .X(net6922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6396 (.A(\rbzero.tex_g0[46] ),
    .X(net6923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6397 (.A(net2035),
    .X(net6924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6398 (.A(_04268_),
    .X(net6925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6399 (.A(net2036),
    .X(net6926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net5992),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_01147_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6400 (.A(\rbzero.tex_r1[3] ),
    .X(net6927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6401 (.A(net1958),
    .X(net6928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6402 (.A(_04099_),
    .X(net6929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6403 (.A(net1959),
    .X(net6930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6404 (.A(\rbzero.tex_b0[9] ),
    .X(net6931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6405 (.A(net2072),
    .X(net6932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6406 (.A(_04449_),
    .X(net6933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6407 (.A(net2073),
    .X(net6934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6408 (.A(\rbzero.tex_g0[20] ),
    .X(net6935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6409 (.A(net2265),
    .X(net6936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(net6230),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6410 (.A(\rbzero.spi_registers.new_leak[0] ),
    .X(net6937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6411 (.A(net2447),
    .X(net6938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6412 (.A(\rbzero.tex_r1[61] ),
    .X(net6939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6413 (.A(net2026),
    .X(net6940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6414 (.A(\rbzero.tex_b0[33] ),
    .X(net6941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6415 (.A(net1773),
    .X(net6942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6416 (.A(_04422_),
    .X(net6943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6417 (.A(net1774),
    .X(net6944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6418 (.A(\rbzero.tex_b0[62] ),
    .X(net6945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6419 (.A(net2082),
    .X(net6946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(net6232),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6420 (.A(\rbzero.tex_b1[23] ),
    .X(net6947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6421 (.A(net2274),
    .X(net6948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6422 (.A(_04363_),
    .X(net6949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6423 (.A(net2275),
    .X(net6950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6424 (.A(\rbzero.tex_r1[51] ),
    .X(net6951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6425 (.A(net2496),
    .X(net6952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6426 (.A(\rbzero.pov.ready_buffer[25] ),
    .X(net6953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6427 (.A(net2485),
    .X(net6954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6428 (.A(\rbzero.tex_b1[5] ),
    .X(net6955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6429 (.A(net2149),
    .X(net6956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(_00660_),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6430 (.A(_04383_),
    .X(net6957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6431 (.A(net2150),
    .X(net6958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6432 (.A(\rbzero.spi_registers.new_vshift[5] ),
    .X(net6959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6433 (.A(net2223),
    .X(net6960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6434 (.A(_03394_),
    .X(net6961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6435 (.A(\rbzero.tex_r0[9] ),
    .X(net6962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6436 (.A(net2122),
    .X(net6963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6437 (.A(_04166_),
    .X(net6964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6438 (.A(net2144),
    .X(net6965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6439 (.A(\rbzero.tex_r1[5] ),
    .X(net6966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(net4590),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6440 (.A(net2324),
    .X(net6967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6441 (.A(\rbzero.tex_b0[5] ),
    .X(net6968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6442 (.A(net1943),
    .X(net6969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6443 (.A(_04453_),
    .X(net6970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6444 (.A(net1944),
    .X(net6971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6445 (.A(\rbzero.tex_b0[59] ),
    .X(net6972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6446 (.A(net2279),
    .X(net6973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6447 (.A(\rbzero.tex_r1[45] ),
    .X(net6974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6448 (.A(net2229),
    .X(net6975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6449 (.A(_04052_),
    .X(net6976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(net4592),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6450 (.A(net2230),
    .X(net6977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6451 (.A(\rbzero.tex_r0[17] ),
    .X(net6978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6452 (.A(net2339),
    .X(net6979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6453 (.A(_04157_),
    .X(net6980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6454 (.A(net2340),
    .X(net6981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6455 (.A(\rbzero.tex_r0[59] ),
    .X(net6982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6456 (.A(net2530),
    .X(net6983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6457 (.A(\rbzero.tex_r1[23] ),
    .X(net6984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6458 (.A(net2173),
    .X(net6985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6459 (.A(\rbzero.tex_b0[31] ),
    .X(net6986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(net6210),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6460 (.A(net2456),
    .X(net6987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6461 (.A(\rbzero.tex_r0[20] ),
    .X(net6988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6462 (.A(net2619),
    .X(net6989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6463 (.A(\rbzero.tex_g1[31] ),
    .X(net6990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6464 (.A(net2566),
    .X(net6991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6465 (.A(_04212_),
    .X(net6992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6466 (.A(net2409),
    .X(net6993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6467 (.A(\rbzero.tex_b0[53] ),
    .X(net6994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6468 (.A(net2167),
    .X(net6995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6469 (.A(_04400_),
    .X(net6996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(net6212),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6470 (.A(net2168),
    .X(net6997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6471 (.A(\rbzero.tex_r1[36] ),
    .X(net6998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6472 (.A(net2560),
    .X(net6999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6473 (.A(\rbzero.tex_g1[30] ),
    .X(net7000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6474 (.A(net2970),
    .X(net7001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6475 (.A(\rbzero.pov.ready_buffer[5] ),
    .X(net7002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6476 (.A(net1970),
    .X(net7003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6477 (.A(\rbzero.tex_g1[10] ),
    .X(net7004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6478 (.A(net2738),
    .X(net7005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6479 (.A(_04235_),
    .X(net7006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_01419_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6480 (.A(net2849),
    .X(net7007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6481 (.A(\rbzero.tex_r0[53] ),
    .X(net7008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6482 (.A(net2247),
    .X(net7009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6483 (.A(_04118_),
    .X(net7010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6484 (.A(net2248),
    .X(net7011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6485 (.A(\rbzero.tex_g0[7] ),
    .X(net7012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6486 (.A(net2354),
    .X(net7013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6487 (.A(\rbzero.tex_g1[47] ),
    .X(net7014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6488 (.A(net2288),
    .X(net7015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6489 (.A(\rbzero.tex_r0[34] ),
    .X(net7016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(net6463),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6490 (.A(net2094),
    .X(net7017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6491 (.A(\rbzero.tex_r0[40] ),
    .X(net7018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6492 (.A(net2043),
    .X(net7019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6493 (.A(\rbzero.pov.ready_buffer[15] ),
    .X(net7020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6494 (.A(net2161),
    .X(net7021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6495 (.A(\rbzero.tex_b0[6] ),
    .X(net7022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6496 (.A(net2315),
    .X(net7023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6497 (.A(\rbzero.tex_b0[39] ),
    .X(net7024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6498 (.A(net1929),
    .X(net7025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6499 (.A(_04416_),
    .X(net7026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_01473_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_03150_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6500 (.A(net1930),
    .X(net7027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6501 (.A(\rbzero.tex_g1[54] ),
    .X(net7028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6502 (.A(net2417),
    .X(net7029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6503 (.A(_04187_),
    .X(net7030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6504 (.A(net2418),
    .X(net7031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6505 (.A(\rbzero.tex_g0[43] ),
    .X(net7032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6506 (.A(net2453),
    .X(net7033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6507 (.A(\rbzero.tex_r0[6] ),
    .X(net7034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6508 (.A(net2761),
    .X(net7035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6509 (.A(_04169_),
    .X(net7036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(net4370),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6510 (.A(net2762),
    .X(net7037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6511 (.A(\rbzero.tex_b1[40] ),
    .X(net7038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6512 (.A(net2509),
    .X(net7039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6513 (.A(_04345_),
    .X(net7040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6514 (.A(net2510),
    .X(net7041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6515 (.A(\rbzero.tex_g1[9] ),
    .X(net7042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6516 (.A(net2965),
    .X(net7043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6517 (.A(\rbzero.pov.ready_buffer[16] ),
    .X(net7044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6518 (.A(net2125),
    .X(net7045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6519 (.A(_03011_),
    .X(net7046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(net6222),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6520 (.A(net2126),
    .X(net7047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6521 (.A(\rbzero.tex_g1[6] ),
    .X(net7048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6522 (.A(net2399),
    .X(net7049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6523 (.A(\rbzero.tex_g0[49] ),
    .X(net7050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6524 (.A(net1964),
    .X(net7051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6525 (.A(_04263_),
    .X(net7052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6526 (.A(net1965),
    .X(net7053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6527 (.A(\rbzero.tex_r1[18] ),
    .X(net7054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6528 (.A(net2641),
    .X(net7055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6529 (.A(\rbzero.tex_g0[44] ),
    .X(net7056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(net6224),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6530 (.A(net2235),
    .X(net7057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6531 (.A(\rbzero.tex_b0[37] ),
    .X(net7058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6532 (.A(net2211),
    .X(net7059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6533 (.A(_04418_),
    .X(net7060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6534 (.A(net2212),
    .X(net7061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6535 (.A(\rbzero.tex_r1[41] ),
    .X(net7062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6536 (.A(net2259),
    .X(net7063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6537 (.A(_04056_),
    .X(net7064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6538 (.A(net2658),
    .X(net7065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6539 (.A(\rbzero.tex_r0[56] ),
    .X(net7066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_01410_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6540 (.A(net2327),
    .X(net7067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6541 (.A(_04114_),
    .X(net7068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6542 (.A(net2328),
    .X(net7069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6543 (.A(\rbzero.tex_g0[25] ),
    .X(net7070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6544 (.A(net2217),
    .X(net7071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6545 (.A(_04291_),
    .X(net7072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6546 (.A(net2218),
    .X(net7073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6547 (.A(\rbzero.tex_b1[11] ),
    .X(net7074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6548 (.A(net2664),
    .X(net7075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6549 (.A(_04377_),
    .X(net7076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(net6246),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6550 (.A(net2665),
    .X(net7077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6551 (.A(\rbzero.tex_g1[45] ),
    .X(net7078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6552 (.A(net2750),
    .X(net7079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6553 (.A(_04198_),
    .X(net7080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6554 (.A(net2751),
    .X(net7081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6555 (.A(\rbzero.pov.ready_buffer[43] ),
    .X(net7082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6556 (.A(net775),
    .X(net7083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6557 (.A(\rbzero.spi_registers.new_mapd[8] ),
    .X(net7084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6558 (.A(net836),
    .X(net7085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6559 (.A(\rbzero.tex_r1[26] ),
    .X(net7086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_03533_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6560 (.A(net2981),
    .X(net7087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6561 (.A(\rbzero.tex_b0[35] ),
    .X(net7088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6562 (.A(net2725),
    .X(net7089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6563 (.A(\rbzero.tex_g1[42] ),
    .X(net7090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6564 (.A(net2432),
    .X(net7091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6565 (.A(\rbzero.pov.ready_buffer[42] ),
    .X(net7092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6566 (.A(net779),
    .X(net7093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6567 (.A(\rbzero.tex_r0[15] ),
    .X(net7094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6568 (.A(net2187),
    .X(net7095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6569 (.A(\rbzero.tex_b1[10] ),
    .X(net7096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_01100_),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6570 (.A(net2601),
    .X(net7097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6571 (.A(\rbzero.tex_b1[37] ),
    .X(net7098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6572 (.A(net2357),
    .X(net7099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6573 (.A(\rbzero.tex_b1[57] ),
    .X(net7100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6574 (.A(net2113),
    .X(net7101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6575 (.A(\rbzero.tex_r0[60] ),
    .X(net7102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6576 (.A(net1842),
    .X(net7103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6577 (.A(\rbzero.tex_g1[39] ),
    .X(net7104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6578 (.A(net2176),
    .X(net7105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6579 (.A(\rbzero.tex_b0[28] ),
    .X(net7106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(net6218),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6580 (.A(net2527),
    .X(net7107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6581 (.A(_04428_),
    .X(net7108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6582 (.A(net2528),
    .X(net7109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6583 (.A(\rbzero.tex_g1[7] ),
    .X(net7110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6584 (.A(net2023),
    .X(net7111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6585 (.A(\rbzero.tex_b0[4] ),
    .X(net7112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6586 (.A(net2164),
    .X(net7113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6587 (.A(_04454_),
    .X(net7114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6588 (.A(net2165),
    .X(net7115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6589 (.A(\rbzero.tex_g1[62] ),
    .X(net7116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(net6220),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6590 (.A(net2747),
    .X(net7117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6591 (.A(\rbzero.tex_b0[14] ),
    .X(net7118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6592 (.A(net2170),
    .X(net7119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6593 (.A(\rbzero.tex_r1[62] ),
    .X(net7120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6594 (.A(net2548),
    .X(net7121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6595 (.A(\rbzero.tex_r1[52] ),
    .X(net7122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6596 (.A(net2688),
    .X(net7123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6597 (.A(\rbzero.tex_b0[19] ),
    .X(net7124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6598 (.A(net2679),
    .X(net7125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6599 (.A(_04438_),
    .X(net7126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net4927),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_01313_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6600 (.A(net2680),
    .X(net7127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6601 (.A(\rbzero.tex_r0[21] ),
    .X(net7128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6602 (.A(net2032),
    .X(net7129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6603 (.A(\rbzero.tex_g0[59] ),
    .X(net7130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6604 (.A(net2420),
    .X(net7131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6605 (.A(_04252_),
    .X(net7132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6606 (.A(net2421),
    .X(net7133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6607 (.A(\rbzero.tex_r0[57] ),
    .X(net7134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6608 (.A(net2201),
    .X(net7135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6609 (.A(\rbzero.tex_g1[43] ),
    .X(net7136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(net6226),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6610 (.A(net2551),
    .X(net7137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6611 (.A(_04199_),
    .X(net7138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6612 (.A(net2377),
    .X(net7139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6613 (.A(\rbzero.tex_r0[55] ),
    .X(net7140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6614 (.A(net2384),
    .X(net7141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6615 (.A(\rbzero.pov.ready_buffer[26] ),
    .X(net7142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6616 (.A(net1915),
    .X(net7143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6617 (.A(\rbzero.tex_g0[60] ),
    .X(net7144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6618 (.A(net2291),
    .X(net7145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6619 (.A(\rbzero.tex_b0[36] ),
    .X(net7146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(net6228),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6620 (.A(net2841),
    .X(net7147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6621 (.A(\rbzero.tex_r0[23] ),
    .X(net7148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6622 (.A(net2294),
    .X(net7149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6623 (.A(_04151_),
    .X(net7150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6624 (.A(net2295),
    .X(net7151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6625 (.A(\rbzero.tex_g1[26] ),
    .X(net7152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6626 (.A(net2515),
    .X(net7153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6627 (.A(\rbzero.pov.ready_buffer[17] ),
    .X(net7154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6628 (.A(net762),
    .X(net7155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6629 (.A(\rbzero.tex_b1[54] ),
    .X(net7156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(_01463_),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6630 (.A(net2208),
    .X(net7157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6631 (.A(_04329_),
    .X(net7158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6632 (.A(net2209),
    .X(net7159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6633 (.A(\rbzero.tex_r1[43] ),
    .X(net7160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6634 (.A(net2011),
    .X(net7161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6635 (.A(_04055_),
    .X(net7162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6636 (.A(net2012),
    .X(net7163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6637 (.A(\rbzero.tex_r1[44] ),
    .X(net7164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6638 (.A(net2499),
    .X(net7165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6639 (.A(\rbzero.tex_g0[41] ),
    .X(net7166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net6242),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6640 (.A(net2282),
    .X(net7167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6641 (.A(_04273_),
    .X(net7168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6642 (.A(net2283),
    .X(net7169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6643 (.A(\rbzero.tex_g1[22] ),
    .X(net7170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6644 (.A(net2402),
    .X(net7171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6645 (.A(_04223_),
    .X(net7172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6646 (.A(net2403),
    .X(net7173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6647 (.A(\rbzero.pov.spi_buffer[65] ),
    .X(net7174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6648 (.A(net2190),
    .X(net7175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6649 (.A(_03590_),
    .X(net7176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(net6244),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6650 (.A(\rbzero.pov.spi_buffer[44] ),
    .X(net7177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6651 (.A(net2069),
    .X(net7178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6652 (.A(\rbzero.tex_g1[36] ),
    .X(net7179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6653 (.A(net2569),
    .X(net7180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6654 (.A(_04208_),
    .X(net7181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6655 (.A(net2570),
    .X(net7182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6656 (.A(\rbzero.tex_r0[50] ),
    .X(net7183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6657 (.A(net2676),
    .X(net7184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6658 (.A(\rbzero.tex_g0[54] ),
    .X(net7185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6659 (.A(net2691),
    .X(net7186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_01451_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6660 (.A(\rbzero.pov.ready_buffer[20] ),
    .X(net7187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6661 (.A(net791),
    .X(net7188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6662 (.A(\rbzero.tex_g0[33] ),
    .X(net7189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6663 (.A(net2616),
    .X(net7190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6664 (.A(\rbzero.tex_r1[24] ),
    .X(net7191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6665 (.A(net2465),
    .X(net7192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6666 (.A(\rbzero.tex_g0[14] ),
    .X(net7193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6667 (.A(net2491),
    .X(net7194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6668 (.A(\rbzero.tex_b1[42] ),
    .X(net7195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6669 (.A(net2554),
    .X(net7196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(net2770),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6670 (.A(_04343_),
    .X(net7197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6671 (.A(net2555),
    .X(net7198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6672 (.A(\rbzero.tex_r0[51] ),
    .X(net7199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6673 (.A(net2444),
    .X(net7200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6674 (.A(\rbzero.tex_b0[26] ),
    .X(net7201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6675 (.A(net2607),
    .X(net7202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6676 (.A(\rbzero.tex_b0[52] ),
    .X(net7203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6677 (.A(net2387),
    .X(net7204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6678 (.A(_04402_),
    .X(net7205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6679 (.A(net2388),
    .X(net7206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_03007_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6680 (.A(\rbzero.tex_r0[18] ),
    .X(net7207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6681 (.A(net2450),
    .X(net7208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6682 (.A(\rbzero.tex_g1[34] ),
    .X(net7209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6683 (.A(net2459),
    .X(net7210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6684 (.A(\rbzero.tex_g0[2] ),
    .X(net7211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6685 (.A(net655),
    .X(net7212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6686 (.A(_04315_),
    .X(net7213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6687 (.A(net2858),
    .X(net7214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6688 (.A(\rbzero.tex_g0[58] ),
    .X(net7215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6689 (.A(net2685),
    .X(net7216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_00659_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6690 (.A(\rbzero.tex_b1[41] ),
    .X(net7217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6691 (.A(net2777),
    .X(net7218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6692 (.A(\rbzero.tex_r0[22] ),
    .X(net7219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6693 (.A(net2635),
    .X(net7220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6694 (.A(\rbzero.tex_r0[26] ),
    .X(net7221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6695 (.A(net2625),
    .X(net7222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6696 (.A(\rbzero.tex_r0[30] ),
    .X(net7223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6697 (.A(net2390),
    .X(net7224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6698 (.A(\rbzero.tex_r1[14] ),
    .X(net7225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6699 (.A(net2342),
    .X(net7226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net4929),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(net6459),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6700 (.A(\rbzero.tex_g0[16] ),
    .X(net7227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6701 (.A(net2017),
    .X(net7228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6702 (.A(_04301_),
    .X(net7229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6703 (.A(net2018),
    .X(net7230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6704 (.A(\rbzero.tex_g0[27] ),
    .X(net7231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6705 (.A(net2722),
    .X(net7232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6706 (.A(\rbzero.tex_g0[34] ),
    .X(net7233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6707 (.A(net2731),
    .X(net7234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6708 (.A(\rbzero.tex_r1[56] ),
    .X(net7235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6709 (.A(net2851),
    .X(net7236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(net6461),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6710 (.A(\rbzero.tex_r0[36] ),
    .X(net7237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6711 (.A(net2755),
    .X(net7238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6712 (.A(\rbzero.tex_b1[55] ),
    .X(net7239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6713 (.A(net2253),
    .X(net7240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6714 (.A(\rbzero.tex_b0[56] ),
    .X(net7241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6715 (.A(net2512),
    .X(net7242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6716 (.A(\rbzero.tex_b0[49] ),
    .X(net7243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6717 (.A(net2572),
    .X(net7244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6718 (.A(_04405_),
    .X(net7245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6719 (.A(net2573),
    .X(net7246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_01067_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6720 (.A(\rbzero.tex_b0[38] ),
    .X(net7247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6721 (.A(net2381),
    .X(net7248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6722 (.A(\rbzero.tex_g1[23] ),
    .X(net7249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6723 (.A(net2651),
    .X(net7250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6724 (.A(\rbzero.tex_r0[5] ),
    .X(net7251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6725 (.A(net2592),
    .X(net7252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6726 (.A(\rbzero.tex_g0[9] ),
    .X(net7253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6727 (.A(net2670),
    .X(net7254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6728 (.A(_04308_),
    .X(net7255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6729 (.A(net2671),
    .X(net7256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(net6256),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6730 (.A(\rbzero.tex_b0[8] ),
    .X(net7257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6731 (.A(net2832),
    .X(net7258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6732 (.A(_04450_),
    .X(net7259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6733 (.A(net2833),
    .X(net7260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6734 (.A(\rbzero.tex_g1[52] ),
    .X(net7261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6735 (.A(net2820),
    .X(net7262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6736 (.A(_04189_),
    .X(net7263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6737 (.A(net2821),
    .X(net7264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6738 (.A(\rbzero.tex_r1[8] ),
    .X(net7265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6739 (.A(net2524),
    .X(net7266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_03828_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6740 (.A(\rbzero.tex_r1[47] ),
    .X(net7267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6741 (.A(net2984),
    .X(net7268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6742 (.A(\rbzero.tex_b0[32] ),
    .X(net7269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6743 (.A(net2744),
    .X(net7270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6744 (.A(\rbzero.pov.sclk_buffer[2] ),
    .X(net7271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6745 (.A(net3305),
    .X(net7272));
 sky130_fd_sc_hd__buf_2 hold6746 (.A(_03486_),
    .X(net7273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6747 (.A(\rbzero.tex_g1[51] ),
    .X(net7274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6748 (.A(net2518),
    .X(net7275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6749 (.A(\rbzero.spi_registers.ss_buffer[0] ),
    .X(net7276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(_01266_),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6750 (.A(net2435),
    .X(net7277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6751 (.A(\rbzero.tex_g0[45] ),
    .X(net7278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6752 (.A(net2589),
    .X(net7279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6753 (.A(\rbzero.tex_b0[12] ),
    .X(net7280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6754 (.A(net2911),
    .X(net7281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6755 (.A(_04446_),
    .X(net7282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6756 (.A(net2912),
    .X(net7283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6757 (.A(\rbzero.tex_r0[8] ),
    .X(net7284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6758 (.A(net2143),
    .X(net7285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6759 (.A(\rbzero.tex_r0[62] ),
    .X(net7286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(net6596),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6760 (.A(net2786),
    .X(net7287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6761 (.A(_04108_),
    .X(net7288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6762 (.A(net2787),
    .X(net7289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6763 (.A(\rbzero.tex_g0[51] ),
    .X(net7290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6764 (.A(net2575),
    .X(net7291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6765 (.A(\rbzero.tex_g1[19] ),
    .X(net7292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6766 (.A(net2638),
    .X(net7293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6767 (.A(\rbzero.tex_r1[34] ),
    .X(net7294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6768 (.A(net2774),
    .X(net7295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6769 (.A(\rbzero.tex_b0[22] ),
    .X(net7296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(_03151_),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6770 (.A(net2479),
    .X(net7297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6771 (.A(\rbzero.tex_r0[31] ),
    .X(net7298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6772 (.A(net2155),
    .X(net7299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6773 (.A(\rbzero.tex_b0[23] ),
    .X(net7300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6774 (.A(net2854),
    .X(net7301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6775 (.A(\rbzero.spi_registers.new_mapd[5] ),
    .X(net7302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6776 (.A(net957),
    .X(net7303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6777 (.A(_03409_),
    .X(net7304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6778 (.A(\rbzero.tex_b1[19] ),
    .X(net7305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6779 (.A(net2694),
    .X(net7306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(net4421),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6780 (.A(_04368_),
    .X(net7307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6781 (.A(net2695),
    .X(net7308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6782 (.A(\rbzero.pov.spi_buffer[6] ),
    .X(net7309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6783 (.A(net1682),
    .X(net7310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6784 (.A(\rbzero.pov.mosi ),
    .X(net7311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6785 (.A(net1814),
    .X(net7312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6786 (.A(\rbzero.tex_g0[8] ),
    .X(net7313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6787 (.A(net2715),
    .X(net7314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6788 (.A(\rbzero.tex_g0[24] ),
    .X(net7315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6789 (.A(net2300),
    .X(net7316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(net6276),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6790 (.A(_04292_),
    .X(net7317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6791 (.A(net2301),
    .X(net7318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6792 (.A(\rbzero.tex_b0[11] ),
    .X(net7319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6793 (.A(net2892),
    .X(net7320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6794 (.A(\rbzero.tex_b1[22] ),
    .X(net7321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6795 (.A(net3092),
    .X(net7322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6796 (.A(\rbzero.tex_r1[9] ),
    .X(net7323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6797 (.A(net2370),
    .X(net7324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6798 (.A(\rbzero.tex_r0[37] ),
    .X(net7325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6799 (.A(net2950),
    .X(net7326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net4931),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(net6278),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6800 (.A(\rbzero.tex_r1[49] ),
    .X(net7327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6801 (.A(net2438),
    .X(net7328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6802 (.A(_04048_),
    .X(net7329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6803 (.A(net2439),
    .X(net7330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6804 (.A(\rbzero.tex_b0[16] ),
    .X(net7331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6805 (.A(net2345),
    .X(net7332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6806 (.A(\rbzero.pov.ready_buffer[40] ),
    .X(net7333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6807 (.A(net816),
    .X(net7334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6808 (.A(\rbzero.tex_g1[21] ),
    .X(net7335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6809 (.A(net2521),
    .X(net7336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(_01498_),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6810 (.A(\rbzero.tex_b1[53] ),
    .X(net7337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6811 (.A(net2545),
    .X(net7338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6812 (.A(\rbzero.tex_g1[17] ),
    .X(net7339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6813 (.A(net2783),
    .X(net7340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6814 (.A(\rbzero.tex_b1[4] ),
    .X(net7341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6815 (.A(net2930),
    .X(net7342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6816 (.A(\rbzero.tex_b1[43] ),
    .X(net7343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6817 (.A(net2937),
    .X(net7344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6818 (.A(\rbzero.tex_b1[38] ),
    .X(net7345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6819 (.A(net2706),
    .X(net7346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(net5483),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6820 (.A(\rbzero.tex_r0[16] ),
    .X(net7347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6821 (.A(net2728),
    .X(net7348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6822 (.A(\rbzero.tex_r1[30] ),
    .X(net7349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6823 (.A(\rbzero.tex_g1[3] ),
    .X(net7350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6824 (.A(net2462),
    .X(net7351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6825 (.A(_04243_),
    .X(net7352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6826 (.A(net2596),
    .X(net7353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6827 (.A(\rbzero.tex_g0[55] ),
    .X(net7354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6828 (.A(net2923),
    .X(net7355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6829 (.A(_04256_),
    .X(net7356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(net5485),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6830 (.A(net2887),
    .X(net7357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6831 (.A(\rbzero.tex_r1[48] ),
    .X(net7358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6832 (.A(net3128),
    .X(net7359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6833 (.A(\rbzero.tex_g0[23] ),
    .X(net7360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6834 (.A(net2482),
    .X(net7361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6835 (.A(\rbzero.tex_b0[51] ),
    .X(net7362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6836 (.A(net2539),
    .X(net7363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6837 (.A(\rbzero.tex_r1[53] ),
    .X(net7364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6838 (.A(net2780),
    .X(net7365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6839 (.A(\rbzero.pov.spi_buffer[51] ),
    .X(net7366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(net6252),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6840 (.A(net2411),
    .X(net7367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6841 (.A(\rbzero.tex_r0[47] ),
    .X(net7368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6842 (.A(net2581),
    .X(net7369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6843 (.A(_04124_),
    .X(net7370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6844 (.A(net2611),
    .X(net7371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6845 (.A(\rbzero.tex_g1[29] ),
    .X(net7372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6846 (.A(net3169),
    .X(net7373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6847 (.A(\rbzero.tex_b0[3] ),
    .X(net7374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6848 (.A(net2895),
    .X(net7375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6849 (.A(\rbzero.tex_b0[48] ),
    .X(net7376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(net6254),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6850 (.A(net2488),
    .X(net7377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6851 (.A(_04406_),
    .X(net7378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6852 (.A(net2489),
    .X(net7379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6853 (.A(\rbzero.tex_g1[40] ),
    .X(net7380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6854 (.A(net2533),
    .X(net7381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6855 (.A(\rbzero.tex_b1[18] ),
    .X(net7382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6856 (.A(net2557),
    .X(net7383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6857 (.A(_04369_),
    .X(net7384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6858 (.A(net2558),
    .X(net7385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6859 (.A(\rbzero.tex_b0[18] ),
    .X(net7386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_00968_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6860 (.A(net2917),
    .X(net7387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6861 (.A(\rbzero.tex_b1[59] ),
    .X(net7388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6862 (.A(net2285),
    .X(net7389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6863 (.A(\rbzero.tex_b0[41] ),
    .X(net7390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6864 (.A(net2673),
    .X(net7391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6865 (.A(\rbzero.tex_b0[42] ),
    .X(net7392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6866 (.A(net2813),
    .X(net7393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6867 (.A(\rbzero.spi_registers.new_mapd[3] ),
    .X(net7394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6868 (.A(net3002),
    .X(net7395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6869 (.A(\rbzero.tex_g0[40] ),
    .X(net7396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net6264),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6870 (.A(net3070),
    .X(net7397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6871 (.A(\rbzero.tex_g1[35] ),
    .X(net7398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6872 (.A(net2471),
    .X(net7399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6873 (.A(\rbzero.tex_b1[39] ),
    .X(net7400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6874 (.A(net2333),
    .X(net7401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6875 (.A(\rbzero.tex_r0[52] ),
    .X(net7402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6876 (.A(net2959),
    .X(net7403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6877 (.A(\rbzero.tex_b0[54] ),
    .X(net7404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6878 (.A(net2987),
    .X(net7405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6879 (.A(\rbzero.tex_b1[17] ),
    .X(net7406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_03823_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6880 (.A(net2367),
    .X(net7407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6881 (.A(\rbzero.pov.ready_buffer[11] ),
    .X(net7408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6882 (.A(net2943),
    .X(net7409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6883 (.A(_03006_),
    .X(net7410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6884 (.A(net2944),
    .X(net7411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6885 (.A(\rbzero.tex_b0[7] ),
    .X(net7412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6886 (.A(net3005),
    .X(net7413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6887 (.A(\rbzero.tex_r0[61] ),
    .X(net7414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6888 (.A(net2914),
    .X(net7415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6889 (.A(\rbzero.tex_b0[43] ),
    .X(net7416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_01262_),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6890 (.A(net2654),
    .X(net7417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6891 (.A(\rbzero.pov.ready_buffer[2] ),
    .X(net7418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6892 (.A(net683),
    .X(net7419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6893 (.A(_02996_),
    .X(net7420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6894 (.A(net2765),
    .X(net7421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6895 (.A(\rbzero.tex_g0[37] ),
    .X(net7422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6896 (.A(net2604),
    .X(net7423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6897 (.A(\rbzero.pov.sclk_buffer[0] ),
    .X(net7424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6898 (.A(net2889),
    .X(net7425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6899 (.A(\rbzero.tex_g1[53] ),
    .X(net7426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net4933),
    .X(net596));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold690 (.A(net5487),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6900 (.A(net2999),
    .X(net7427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6901 (.A(\rbzero.tex_g1[24] ),
    .X(net7428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6902 (.A(net2996),
    .X(net7429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6903 (.A(\rbzero.tex_g0[61] ),
    .X(net7430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6904 (.A(net2826),
    .X(net7431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6905 (.A(\rbzero.tex_g0[29] ),
    .X(net7432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6906 (.A(net3089),
    .X(net7433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6907 (.A(_04286_),
    .X(net7434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6908 (.A(net3090),
    .X(net7435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6909 (.A(\rbzero.tex_g0[35] ),
    .X(net7436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(net5489),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6910 (.A(net3176),
    .X(net7437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6911 (.A(\rbzero.tex_r1[27] ),
    .X(net7438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6912 (.A(net2152),
    .X(net7439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6913 (.A(\rbzero.tex_r0[43] ),
    .X(net7440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6914 (.A(net2993),
    .X(net7441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6915 (.A(\rbzero.pov.spi_buffer[22] ),
    .X(net7442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6916 (.A(net3022),
    .X(net7443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6917 (.A(_03018_),
    .X(net7444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6918 (.A(net3183),
    .X(net7445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6919 (.A(\rbzero.tex_b0[44] ),
    .X(net7446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(net6179),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6920 (.A(net2804),
    .X(net7447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6921 (.A(\rbzero.pov.spi_buffer[62] ),
    .X(net7448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6922 (.A(net2712),
    .X(net7449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6923 (.A(\rbzero.tex_b1[50] ),
    .X(net7450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6924 (.A(net2667),
    .X(net7451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6925 (.A(\rbzero.pov.spi_buffer[46] ),
    .X(net7452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6926 (.A(net3134),
    .X(net7453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6927 (.A(\rbzero.pov.spi_buffer[59] ),
    .X(net7454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6928 (.A(net2903),
    .X(net7455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6929 (.A(\rbzero.tex_r1[31] ),
    .X(net7456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(net6181),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6930 (.A(net2373),
    .X(net7457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6931 (.A(\rbzero.tex_b0[27] ),
    .X(net7458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6932 (.A(net2962),
    .X(net7459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6933 (.A(\rbzero.pov.ready_buffer[41] ),
    .X(net7460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6934 (.A(net3131),
    .X(net7461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6935 (.A(_03039_),
    .X(net7462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6936 (.A(net3132),
    .X(net7463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6937 (.A(\rbzero.pov.ready_buffer[55] ),
    .X(net7464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6938 (.A(net663),
    .X(net7465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6939 (.A(_03054_),
    .X(net7466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_01276_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6940 (.A(net2830),
    .X(net7467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6941 (.A(\rbzero.tex_r0[46] ),
    .X(net7468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6942 (.A(net2610),
    .X(net7469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6943 (.A(\rbzero.pov.ready_buffer[46] ),
    .X(net7470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6944 (.A(net3252),
    .X(net7471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6945 (.A(\rbzero.tex_g0[15] ),
    .X(net7472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6946 (.A(net3029),
    .X(net7473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6947 (.A(\rbzero.spi_registers.new_mapd[7] ),
    .X(net7474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6948 (.A(net2066),
    .X(net7475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6949 (.A(\rbzero.tex_g0[48] ),
    .X(net7476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(net6511),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6950 (.A(net2900),
    .X(net7477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6951 (.A(_04266_),
    .X(net7478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6952 (.A(net2901),
    .X(net7479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6953 (.A(\rbzero.pov.ready_buffer[38] ),
    .X(net7480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6954 (.A(net3690),
    .X(net7481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6955 (.A(_03035_),
    .X(net7482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6956 (.A(\rbzero.tex_g0[28] ),
    .X(net7483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6957 (.A(net3263),
    .X(net7484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6958 (.A(\rbzero.tex_g0[31] ),
    .X(net7485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6959 (.A(net3107),
    .X(net7486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(net6513),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6960 (.A(_04284_),
    .X(net7487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6961 (.A(net3108),
    .X(net7488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6962 (.A(\rbzero.pov.ready_buffer[8] ),
    .X(net7489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6963 (.A(net645),
    .X(net7490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6964 (.A(\rbzero.tex_g1[12] ),
    .X(net7491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6965 (.A(net3152),
    .X(net7492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6966 (.A(_04234_),
    .X(net7493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6967 (.A(net3153),
    .X(net7494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6968 (.A(\rbzero.spi_registers.sclk_buffer[1] ),
    .X(net7495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6969 (.A(net2182),
    .X(net7496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_00670_),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6970 (.A(\rbzero.pov.spi_buffer[18] ),
    .X(net7497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6971 (.A(net3155),
    .X(net7498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6972 (.A(\rbzero.tex_g0[47] ),
    .X(net7499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6973 (.A(net3202),
    .X(net7500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6974 (.A(\rbzero.pov.sclk_buffer[1] ),
    .X(net7501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6975 (.A(net3220),
    .X(net7502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6976 (.A(\rbzero.tex_b0[47] ),
    .X(net7503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6977 (.A(net3117),
    .X(net7504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6978 (.A(\rbzero.pov.ss_buffer[1] ),
    .X(net7505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6979 (.A(net2309),
    .X(net7506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(net6270),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6980 (.A(\rbzero.pov.ready_buffer[9] ),
    .X(net7507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6981 (.A(net676),
    .X(net7508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6982 (.A(\rbzero.pov.spi_buffer[72] ),
    .X(net7509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6983 (.A(net1869),
    .X(net7510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6984 (.A(_03072_),
    .X(net7511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6985 (.A(net3346),
    .X(net7512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6986 (.A(\rbzero.tex_g1[13] ),
    .X(net7513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6987 (.A(net3249),
    .X(net7514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6988 (.A(\rbzero.pov.spi_buffer[31] ),
    .X(net7515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6989 (.A(net3233),
    .X(net7516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(net6272),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6990 (.A(\rbzero.tex_r0[13] ),
    .X(net7517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6991 (.A(net3356),
    .X(net7518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6992 (.A(\rbzero.pov.spi_buffer[61] ),
    .X(net7519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6993 (.A(net3286),
    .X(net7520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6994 (.A(\rbzero.spi_registers.new_mapd[6] ),
    .X(net7521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6995 (.A(net1830),
    .X(net7522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6996 (.A(\rbzero.spi_registers.new_other[9] ),
    .X(net7523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6997 (.A(net889),
    .X(net7524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6998 (.A(_03383_),
    .X(net7525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6999 (.A(net2954),
    .X(net7526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net6392),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_01289_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7000 (.A(\rbzero.pov.spi_buffer[3] ),
    .X(net7527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7001 (.A(\rbzero.pov.spi_buffer[12] ),
    .X(net7528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7002 (.A(\rbzero.tex_b1[20] ),
    .X(net7529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7003 (.A(net3243),
    .X(net7530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7004 (.A(\rbzero.tex_g0[30] ),
    .X(net7531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7005 (.A(net3246),
    .X(net7532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7006 (.A(\rbzero.pov.spi_buffer[41] ),
    .X(net7533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7007 (.A(net3166),
    .X(net7534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7008 (.A(\rbzero.pov.ready_buffer[62] ),
    .X(net7535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7009 (.A(net3269),
    .X(net7536));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold701 (.A(net5479),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7010 (.A(\rbzero.pov.ready_buffer[7] ),
    .X(net7537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7011 (.A(net2468),
    .X(net7538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7012 (.A(\rbzero.pov.spi_buffer[16] ),
    .X(net7539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7013 (.A(net3063),
    .X(net7540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7014 (.A(\rbzero.pov.spi_buffer[11] ),
    .X(net7541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7015 (.A(net2869),
    .X(net7542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7016 (.A(\rbzero.pov.ready_buffer[28] ),
    .X(net7543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7017 (.A(net1055),
    .X(net7544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7018 (.A(_03024_),
    .X(net7545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7019 (.A(net3180),
    .X(net7546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(net5481),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7020 (.A(\rbzero.pov.ready_buffer[24] ),
    .X(net7547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7021 (.A(net3289),
    .X(net7548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7022 (.A(\rbzero.pov.ready_buffer[31] ),
    .X(net7549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7023 (.A(net3276),
    .X(net7550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7024 (.A(\rbzero.pov.ready_buffer[27] ),
    .X(net7551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7025 (.A(net1059),
    .X(net7552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7026 (.A(\rbzero.pov.spi_buffer[2] ),
    .X(net7553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7027 (.A(net2764),
    .X(net7554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7028 (.A(\rbzero.pov.spi_buffer[28] ),
    .X(net7555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7029 (.A(net3179),
    .X(net7556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(net6356),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7030 (.A(\rbzero.spi_registers.new_other[8] ),
    .X(net7557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7031 (.A(net2709),
    .X(net7558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7032 (.A(\rbzero.pov.spi_buffer[55] ),
    .X(net7559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7033 (.A(net2829),
    .X(net7560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7034 (.A(\gpout0.hpos[4] ),
    .X(net7561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7035 (.A(net4057),
    .X(net7562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7036 (.A(_05087_),
    .X(net7563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7037 (.A(\rbzero.pov.ready_buffer[30] ),
    .X(net7564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7038 (.A(net876),
    .X(net7565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7039 (.A(\rbzero.pov.ready_buffer[52] ),
    .X(net7566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_03547_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7040 (.A(net2396),
    .X(net7567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7041 (.A(\rbzero.row_render.vinf ),
    .X(net7568));
 sky130_fd_sc_hd__buf_1 hold7042 (.A(net4450),
    .X(net7569));
 sky130_fd_sc_hd__buf_2 hold7043 (.A(_04907_),
    .X(net7570));
 sky130_fd_sc_hd__clkbuf_4 hold7044 (.A(net4068),
    .X(net7571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7045 (.A(\rbzero.pov.ready_buffer[48] ),
    .X(net7572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7046 (.A(net3414),
    .X(net7573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7047 (.A(\rbzero.wall_tracer.mapY[5] ),
    .X(net7574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7048 (.A(net3447),
    .X(net7575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7049 (.A(_02730_),
    .X(net7576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_01113_),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7050 (.A(net3448),
    .X(net7577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7051 (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .X(net7578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7052 (.A(net3478),
    .X(net7579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7053 (.A(_03101_),
    .X(net7580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7054 (.A(net3482),
    .X(net7581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7055 (.A(\rbzero.pov.ready_buffer[29] ),
    .X(net7582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7056 (.A(net3711),
    .X(net7583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7057 (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .X(net7584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7058 (.A(net1447),
    .X(net7585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7059 (.A(\rbzero.pov.ready_buffer[63] ),
    .X(net7586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(net5491),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7060 (.A(net3543),
    .X(net7587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7061 (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .X(net7588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7062 (.A(net3556),
    .X(net7589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7063 (.A(_03097_),
    .X(net7590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7064 (.A(net3557),
    .X(net7591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7065 (.A(\rbzero.pov.ready_buffer[35] ),
    .X(net7592));
 sky130_fd_sc_hd__buf_1 hold7066 (.A(net1113),
    .X(net7593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7067 (.A(\rbzero.pov.ready_buffer[34] ),
    .X(net7594));
 sky130_fd_sc_hd__buf_1 hold7068 (.A(net2242),
    .X(net7595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7069 (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .X(net7596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(net5493),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7070 (.A(net3481),
    .X(net7597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7071 (.A(_03102_),
    .X(net7598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7072 (.A(net3584),
    .X(net7599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7073 (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .X(net7600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7074 (.A(net3583),
    .X(net7601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7075 (.A(_03103_),
    .X(net7602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7076 (.A(net3632),
    .X(net7603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7077 (.A(\rbzero.pov.ready_buffer[72] ),
    .X(net7604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7078 (.A(net3345),
    .X(net7605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7079 (.A(_03654_),
    .X(net7606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(net6258),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7080 (.A(net3684),
    .X(net7607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7081 (.A(\rbzero.row_render.wall[1] ),
    .X(net7608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7082 (.A(net3648),
    .X(net7609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7083 (.A(_09749_),
    .X(net7610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7084 (.A(net3649),
    .X(net7611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7085 (.A(\rbzero.pov.ready_buffer[32] ),
    .X(net7612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7086 (.A(net3080),
    .X(net7613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7087 (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .X(net7614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7088 (.A(net3674),
    .X(net7615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7089 (.A(_03098_),
    .X(net7616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(net6260),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7090 (.A(net3675),
    .X(net7617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7091 (.A(\gpout0.vpos[4] ),
    .X(net7618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7092 (.A(_03793_),
    .X(net7619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7093 (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .X(net7620));
 sky130_fd_sc_hd__buf_1 hold7094 (.A(net3592),
    .X(net7621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7096 (.A(_03737_),
    .X(net7623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7097 (.A(net3881),
    .X(net7624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7099 (.A(_03733_),
    .X(net7626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_03240_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_01568_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7100 (.A(net3504),
    .X(net7627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7101 (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .X(net7628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7102 (.A(net3866),
    .X(net7629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7103 (.A(\rbzero.wall_tracer.mapX[5] ),
    .X(net7630));
 sky130_fd_sc_hd__buf_1 hold7104 (.A(net3884),
    .X(net7631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7105 (.A(_02750_),
    .X(net7632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7106 (.A(net3885),
    .X(net7633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7107 (.A(\rbzero.debug_overlay.playerY[3] ),
    .X(net7634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7108 (.A(net3473),
    .X(net7635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7109 (.A(_02721_),
    .X(net7636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(net6741),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7110 (.A(_02722_),
    .X(net7637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7112 (.A(_03729_),
    .X(net7639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7113 (.A(net3687),
    .X(net7640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7115 (.A(_03735_),
    .X(net7642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7116 (.A(net3580),
    .X(net7643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7118 (.A(_03741_),
    .X(net7645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7119 (.A(net3712),
    .X(net7646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_03152_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7120 (.A(\rbzero.pov.spi_counter[4] ),
    .X(net7647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7121 (.A(net3921),
    .X(net7648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7122 (.A(_03499_),
    .X(net7649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7123 (.A(_03501_),
    .X(net7650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7125 (.A(_03720_),
    .X(net7652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7126 (.A(net3608),
    .X(net7653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7127 (.A(\rbzero.pov.spi_counter[5] ),
    .X(net7654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7128 (.A(net3823),
    .X(net7655));
 sky130_fd_sc_hd__buf_1 hold7129 (.A(_03502_),
    .X(net7656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(net4432),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7130 (.A(_03504_),
    .X(net7657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7132 (.A(_03716_),
    .X(net7659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7133 (.A(net3436),
    .X(net7660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7135 (.A(_03718_),
    .X(net7662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7136 (.A(net3691),
    .X(net7663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7137 (.A(\rbzero.row_render.wall[0] ),
    .X(net7664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7138 (.A(net3781),
    .X(net7665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7139 (.A(_09748_),
    .X(net7666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(net6298),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7140 (.A(net3782),
    .X(net7667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7141 (.A(\rbzero.map_rom.i_row[4] ),
    .X(net7668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7142 (.A(net3807),
    .X(net7669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7143 (.A(_02726_),
    .X(net7670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7144 (.A(net3808),
    .X(net7671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7145 (.A(\rbzero.pov.spi_counter[3] ),
    .X(net7672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7146 (.A(net3707),
    .X(net7673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7147 (.A(_03496_),
    .X(net7674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7148 (.A(_03498_),
    .X(net7675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7149 (.A(net3709),
    .X(net7676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(_02486_),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7150 (.A(net7743),
    .X(net7677));
 sky130_fd_sc_hd__buf_2 hold7151 (.A(net3954),
    .X(net7678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7152 (.A(_04664_),
    .X(net7679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7153 (.A(\gpout0.vpos[2] ),
    .X(net7680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7154 (.A(net4110),
    .X(net7681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7155 (.A(_01247_),
    .X(net7682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7156 (.A(net3971),
    .X(net7683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7157 (.A(\rbzero.pov.spi_counter[1] ),
    .X(net7684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7158 (.A(net3703),
    .X(net7685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7159 (.A(\rbzero.map_rom.f4 ),
    .X(net7686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_00576_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7160 (.A(net3959),
    .X(net7687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7161 (.A(_02732_),
    .X(net7688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7162 (.A(\rbzero.debug_overlay.playerY[0] ),
    .X(net7689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7163 (.A(net3326),
    .X(net7690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7164 (.A(\rbzero.pov.ready_buffer[73] ),
    .X(net7691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7165 (.A(_03657_),
    .X(net7692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7166 (.A(\rbzero.spi_registers.spi_counter[4] ),
    .X(net7693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7167 (.A(\rbzero.spi_registers.spi_counter[3] ),
    .X(net7694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7168 (.A(_02966_),
    .X(net7695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7169 (.A(\rbzero.spi_registers.spi_counter[2] ),
    .X(net7696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(net6435),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7170 (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .X(net7697));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold7171 (.A(net2953),
    .X(net7698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7172 (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(net7699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7173 (.A(\rbzero.debug_overlay.playerX[3] ),
    .X(net7700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7174 (.A(net3431),
    .X(net7701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7175 (.A(_02742_),
    .X(net7702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7176 (.A(_02743_),
    .X(net7703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7177 (.A(\rbzero.debug_overlay.playerX[4] ),
    .X(net7704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7178 (.A(net3682),
    .X(net7705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7179 (.A(_02745_),
    .X(net7706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(net6437),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7180 (.A(\gpout0.hpos[1] ),
    .X(net7707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7181 (.A(net3857),
    .X(net7708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7182 (.A(\gpout0.hpos[7] ),
    .X(net7709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7183 (.A(net4115),
    .X(net7710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7184 (.A(\rbzero.map_rom.f3 ),
    .X(net7711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7185 (.A(net4033),
    .X(net7712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7186 (.A(_09754_),
    .X(net7713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7187 (.A(_02735_),
    .X(net7714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7188 (.A(\gpout0.vpos[7] ),
    .X(net7715));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold7189 (.A(net4091),
    .X(net7716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(_00680_),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7190 (.A(_01251_),
    .X(net7717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7191 (.A(\rbzero.color_floor[4] ),
    .X(net7718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7192 (.A(net3644),
    .X(net7719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7193 (.A(_05464_),
    .X(net7720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7194 (.A(\rbzero.color_floor[2] ),
    .X(net7721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7195 (.A(net3547),
    .X(net7722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7196 (.A(_05298_),
    .X(net7723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7197 (.A(\rbzero.color_sky[5] ),
    .X(net7724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7198 (.A(net3651),
    .X(net7725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7199 (.A(_05548_),
    .X(net7726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net4199),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(net6262),
    .X(net1247));
 sky130_fd_sc_hd__clkbuf_4 hold7200 (.A(net4173),
    .X(net7727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7201 (.A(\rbzero.spi_registers.got_new_vinf ),
    .X(net7728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7202 (.A(\rbzero.color_floor[0] ),
    .X(net7729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7203 (.A(net3656),
    .X(net7730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7204 (.A(_04908_),
    .X(net7731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7205 (.A(\rbzero.color_sky[3] ),
    .X(net7732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7206 (.A(net3670),
    .X(net7733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7207 (.A(_05381_),
    .X(net7734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7208 (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(net7735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7209 (.A(\rbzero.color_sky[1] ),
    .X(net7736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(_03434_),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7210 (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(net7737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7211 (.A(\gpout0.vpos[6] ),
    .X(net7738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7212 (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(net7739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7214 (.A(_03724_),
    .X(net7741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7215 (.A(\rbzero.spi_registers.got_new_texadd[0] ),
    .X(net7742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7216 (.A(\gpout0.hpos[2] ),
    .X(net7743));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold7217 (.A(net3927),
    .X(net7744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7218 (.A(\rbzero.spi_registers.got_new_vshift ),
    .X(net7745));
 sky130_fd_sc_hd__clkbuf_2 hold7219 (.A(net4002),
    .X(net7746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_00969_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7220 (.A(\rbzero.wall_hot[1] ),
    .X(net7747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7221 (.A(\rbzero.wall_hot[0] ),
    .X(net7748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7222 (.A(\rbzero.trace_state[1] ),
    .X(net7749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7223 (.A(\rbzero.spi_registers.spi_buffer[5] ),
    .X(net7750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7224 (.A(net8315),
    .X(net7751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7225 (.A(net8317),
    .X(net7752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(net5798),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7236 (.A(net8361),
    .X(net7763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7237 (.A(\rbzero.debug_overlay.playerX[-7] ),
    .X(net7764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7238 (.A(net3348),
    .X(net7765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7239 (.A(_09090_),
    .X(net7766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_02987_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7240 (.A(\rbzero.debug_overlay.playerY[-6] ),
    .X(net7767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7241 (.A(net3372),
    .X(net7768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7242 (.A(_09085_),
    .X(net7769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7243 (.A(\rbzero.debug_overlay.playerX[-2] ),
    .X(net7770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7244 (.A(net3461),
    .X(net7771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7245 (.A(_09578_),
    .X(net7772));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold7248 (.A(_06026_),
    .X(net7775));
 sky130_fd_sc_hd__buf_2 hold7249 (.A(_06027_),
    .X(net7776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(net5801),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7250 (.A(_06033_),
    .X(net7777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7251 (.A(_09104_),
    .X(net7778));
 sky130_fd_sc_hd__buf_2 hold7252 (.A(_09105_),
    .X(net7779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7253 (.A(\rbzero.debug_overlay.playerY[-4] ),
    .X(net7780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7254 (.A(net3317),
    .X(net7781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7256 (.A(net8369),
    .X(net7783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7257 (.A(_06547_),
    .X(net7784));
 sky130_fd_sc_hd__buf_2 hold7258 (.A(_07912_),
    .X(net7785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7259 (.A(_06529_),
    .X(net7786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(net5495),
    .X(net1253));
 sky130_fd_sc_hd__clkbuf_2 hold7260 (.A(net530),
    .X(net7787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7261 (.A(\rbzero.wall_tracer.stepDistY[1] ),
    .X(net7788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7262 (.A(net4434),
    .X(net7789));
 sky130_fd_sc_hd__buf_1 hold7266 (.A(_06544_),
    .X(net7793));
 sky130_fd_sc_hd__buf_2 hold7267 (.A(_07989_),
    .X(net7794));
 sky130_fd_sc_hd__clkbuf_2 hold7268 (.A(net8443),
    .X(net7795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7269 (.A(\rbzero.wall_tracer.stepDistY[10] ),
    .X(net7796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(net5497),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7270 (.A(net4412),
    .X(net7797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7271 (.A(net3507),
    .X(net7798));
 sky130_fd_sc_hd__clkbuf_1 hold7272 (.A(net4751),
    .X(net7799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7278 (.A(net550),
    .X(net7805));
 sky130_fd_sc_hd__buf_1 hold7279 (.A(net4703),
    .X(net7806));
 sky130_fd_sc_hd__buf_1 hold728 (.A(net8143),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7280 (.A(net8441),
    .X(net7807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7281 (.A(\rbzero.wall_tracer.stepDistX[7] ),
    .X(net7808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7282 (.A(net4519),
    .X(net7809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7283 (.A(_06493_),
    .X(net7810));
 sky130_fd_sc_hd__buf_2 hold7284 (.A(_06494_),
    .X(net7811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7285 (.A(_06564_),
    .X(net7812));
 sky130_fd_sc_hd__buf_2 hold7286 (.A(_07859_),
    .X(net7813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7287 (.A(\rbzero.wall_tracer.stepDistX[8] ),
    .X(net7814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7288 (.A(net4755),
    .X(net7815));
 sky130_fd_sc_hd__buf_1 hold7289 (.A(net4890),
    .X(net7816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(net5502),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7290 (.A(net8535),
    .X(net7817));
 sky130_fd_sc_hd__clkbuf_4 hold7291 (.A(net4891),
    .X(net7818));
 sky130_fd_sc_hd__buf_1 hold7294 (.A(net4777),
    .X(net7821));
 sky130_fd_sc_hd__buf_1 hold7296 (.A(_06546_),
    .X(net7823));
 sky130_fd_sc_hd__clkbuf_4 hold7297 (.A(_07916_),
    .X(net7824));
 sky130_fd_sc_hd__buf_1 hold7298 (.A(_07957_),
    .X(net7825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7299 (.A(\rbzero.wall_tracer.stepDistY[2] ),
    .X(net7826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net4935),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(net6477),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7300 (.A(net4480),
    .X(net7827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7303 (.A(\rbzero.wall_tracer.stepDistX[2] ),
    .X(net7830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7304 (.A(net4400),
    .X(net7831));
 sky130_fd_sc_hd__clkbuf_1 hold7305 (.A(net4718),
    .X(net7832));
 sky130_fd_sc_hd__buf_2 hold7306 (.A(_06436_),
    .X(net7833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7308 (.A(net8434),
    .X(net7835));
 sky130_fd_sc_hd__buf_2 hold7309 (.A(_08668_),
    .X(net7836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(net6479),
    .X(net1258));
 sky130_fd_sc_hd__clkbuf_4 hold7310 (.A(net7821),
    .X(net7837));
 sky130_fd_sc_hd__clkbuf_2 hold7312 (.A(_06606_),
    .X(net7839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7313 (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .X(net7840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7314 (.A(net3748),
    .X(net7841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7315 (.A(_06551_),
    .X(net7842));
 sky130_fd_sc_hd__buf_2 hold7316 (.A(_07840_),
    .X(net7843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7318 (.A(net563),
    .X(net7845));
 sky130_fd_sc_hd__clkbuf_2 hold7319 (.A(_07924_),
    .X(net7846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_01423_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7320 (.A(\rbzero.wall_tracer.stepDistY[6] ),
    .X(net7847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7321 (.A(net4427),
    .X(net7848));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold7323 (.A(_06557_),
    .X(net7850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7324 (.A(\rbzero.wall_tracer.stepDistY[-5] ),
    .X(net7851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7325 (.A(net4378),
    .X(net7852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7326 (.A(net3450),
    .X(net7853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7327 (.A(\rbzero.traced_texVinit[8] ),
    .X(net7854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7328 (.A(net4228),
    .X(net7855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7329 (.A(net1138),
    .X(net7856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(net6326),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7330 (.A(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(net7857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7331 (.A(net4534),
    .X(net7858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7334 (.A(\rbzero.traced_texVinit[0] ),
    .X(net7861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7335 (.A(net4191),
    .X(net7862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7336 (.A(net647),
    .X(net7863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7339 (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .X(net7866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(net6328),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7340 (.A(net4382),
    .X(net7867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7341 (.A(net3459),
    .X(net7868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7342 (.A(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(net7869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7343 (.A(net4380),
    .X(net7870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7344 (.A(net3460),
    .X(net7871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7345 (.A(\rbzero.wall_tracer.stepDistX[-11] ),
    .X(net7872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7346 (.A(net3821),
    .X(net7873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7347 (.A(\rbzero.wall_tracer.stepDistX[4] ),
    .X(net7874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7348 (.A(net4521),
    .X(net7875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7349 (.A(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(net7876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(_01158_),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7350 (.A(net4350),
    .X(net7877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7351 (.A(net3426),
    .X(net7878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7352 (.A(\rbzero.wall_tracer.stepDistY[4] ),
    .X(net7879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7353 (.A(net4458),
    .X(net7880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7354 (.A(\rbzero.traced_texVinit[10] ),
    .X(net7881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7355 (.A(net4203),
    .X(net7882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7356 (.A(net941),
    .X(net7883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7357 (.A(\rbzero.traced_texVinit[2] ),
    .X(net7884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7358 (.A(net4201),
    .X(net7885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7359 (.A(net950),
    .X(net7886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(net6282),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7360 (.A(\rbzero.traced_texVinit[3] ),
    .X(net7887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7361 (.A(net4210),
    .X(net7888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7362 (.A(net1023),
    .X(net7889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7363 (.A(\rbzero.traced_texVinit[1] ),
    .X(net7890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7364 (.A(net4205),
    .X(net7891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7365 (.A(net1008),
    .X(net7892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7366 (.A(\rbzero.traced_texVinit[5] ),
    .X(net7893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7367 (.A(net4214),
    .X(net7894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7368 (.A(net1086),
    .X(net7895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7369 (.A(\rbzero.traced_texVinit[4] ),
    .X(net7896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(_03821_),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7370 (.A(net4212),
    .X(net7897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7371 (.A(net1075),
    .X(net7898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7372 (.A(\rbzero.traced_texVinit[6] ),
    .X(net7899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7373 (.A(net4218),
    .X(net7900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7374 (.A(net1101),
    .X(net7901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7375 (.A(\rbzero.wall_tracer.stepDistX[3] ),
    .X(net7902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7376 (.A(net4404),
    .X(net7903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7377 (.A(net3492),
    .X(net7904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7378 (.A(\rbzero.row_render.size[1] ),
    .X(net7905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7379 (.A(net4342),
    .X(net7906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_01260_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7380 (.A(net3406),
    .X(net7907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7381 (.A(\rbzero.traced_texVinit[7] ),
    .X(net7908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7382 (.A(net4223),
    .X(net7909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7383 (.A(net1105),
    .X(net7910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7385 (.A(_00500_),
    .X(net7912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7386 (.A(net4243),
    .X(net7913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7387 (.A(net757),
    .X(net7914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7388 (.A(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(net7915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7389 (.A(net4398),
    .X(net7916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(net6320),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7390 (.A(net3475),
    .X(net7917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7391 (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .X(net7918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7392 (.A(net4429),
    .X(net7919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7394 (.A(_00501_),
    .X(net7921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7395 (.A(net4297),
    .X(net7922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7396 (.A(net968),
    .X(net7923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7398 (.A(_00502_),
    .X(net7925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7399 (.A(net4319),
    .X(net7926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net4937),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(net6322),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7400 (.A(net755),
    .X(net7927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7401 (.A(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(net7928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7402 (.A(net4788),
    .X(net7929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7403 (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .X(net7930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7404 (.A(net4505),
    .X(net7931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7406 (.A(_00499_),
    .X(net7933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7407 (.A(net4288),
    .X(net7934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7408 (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(net7935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7409 (.A(net4517),
    .X(net7936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(_00989_),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7410 (.A(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(net7937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7411 (.A(net4352),
    .X(net7938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7412 (.A(net3427),
    .X(net7939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7413 (.A(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(net7940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7414 (.A(net4391),
    .X(net7941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7415 (.A(net3472),
    .X(net7942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7418 (.A(_01209_),
    .X(net7945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7419 (.A(net4410),
    .X(net7946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(net6505),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7420 (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .X(net7947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7421 (.A(net4499),
    .X(net7948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7422 (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .X(net7949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7423 (.A(net4540),
    .X(net7950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7424 (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .X(net7951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7425 (.A(net4564),
    .X(net7952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7426 (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .X(net7953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7427 (.A(net4525),
    .X(net7954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7428 (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(net7955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7429 (.A(net4566),
    .X(net7956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(net6507),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7430 (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .X(net7957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7431 (.A(net4568),
    .X(net7958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7432 (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .X(net7959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7433 (.A(net4574),
    .X(net7960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7434 (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .X(net7961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7435 (.A(net4588),
    .X(net7962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7436 (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .X(net7963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7437 (.A(net4609),
    .X(net7964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7438 (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .X(net7965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7439 (.A(net3789),
    .X(net7966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_01359_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7440 (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .X(net7967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7441 (.A(net3802),
    .X(net7968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7442 (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .X(net7969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7443 (.A(net4650),
    .X(net7970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7444 (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(net7971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7445 (.A(net3846),
    .X(net7972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7446 (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .X(net7973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7447 (.A(net4654),
    .X(net7974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7448 (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .X(net7975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7449 (.A(net4656),
    .X(net7976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(net6499),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7450 (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .X(net7977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7451 (.A(net4668),
    .X(net7978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7452 (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .X(net7979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7453 (.A(net4658),
    .X(net7980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7454 (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .X(net7981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7455 (.A(net4507),
    .X(net7982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7456 (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .X(net7983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7457 (.A(net3750),
    .X(net7984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7458 (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .X(net7985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7459 (.A(net4664),
    .X(net7986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(net6501),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7460 (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .X(net7987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7461 (.A(net4546),
    .X(net7988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7462 (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .X(net7989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7463 (.A(net3810),
    .X(net7990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7464 (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .X(net7991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7465 (.A(net3819),
    .X(net7992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7466 (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .X(net7993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7467 (.A(net3834),
    .X(net7994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7468 (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .X(net7995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7469 (.A(net4580),
    .X(net7996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(_01351_),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7470 (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .X(net7997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7471 (.A(net3925),
    .X(net7998));
 sky130_fd_sc_hd__clkbuf_2 hold7472 (.A(net4690),
    .X(net7999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7473 (.A(_00512_),
    .X(net8000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7474 (.A(net4221),
    .X(net8001));
 sky130_fd_sc_hd__clkbuf_4 hold7475 (.A(net8264),
    .X(net8002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7476 (.A(_00516_),
    .X(net8003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7477 (.A(net4234),
    .X(net8004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7478 (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .X(net8005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7479 (.A(net4722),
    .X(net8006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(net5557),
    .X(net1275));
 sky130_fd_sc_hd__buf_1 hold7480 (.A(net4737),
    .X(net8007));
 sky130_fd_sc_hd__clkbuf_4 hold7481 (.A(_08533_),
    .X(net8008));
 sky130_fd_sc_hd__buf_2 hold7482 (.A(net4757),
    .X(net8009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7483 (.A(_00514_),
    .X(net8010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7484 (.A(net4263),
    .X(net8011));
 sky130_fd_sc_hd__buf_2 hold7485 (.A(net8007),
    .X(net8012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7486 (.A(_00513_),
    .X(net8013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7487 (.A(net4254),
    .X(net8014));
 sky130_fd_sc_hd__clkbuf_4 hold7488 (.A(net8270),
    .X(net8015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7489 (.A(_00515_),
    .X(net8016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(net5559),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7490 (.A(net4248),
    .X(net8017));
 sky130_fd_sc_hd__clkbuf_2 hold7491 (.A(net4550),
    .X(net8018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7492 (.A(_00508_),
    .X(net8019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7493 (.A(net4240),
    .X(net8020));
 sky130_fd_sc_hd__buf_2 hold7494 (.A(net4576),
    .X(net8021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7495 (.A(_00509_),
    .X(net8022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7496 (.A(net4257),
    .X(net8023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7498 (.A(_02800_),
    .X(net8025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7499 (.A(_02802_),
    .X(net8026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net4921),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_01534_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7500 (.A(_02803_),
    .X(net8027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7501 (.A(_00628_),
    .X(net8028));
 sky130_fd_sc_hd__clkbuf_2 hold7502 (.A(net4584),
    .X(net8029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7503 (.A(_00510_),
    .X(net8030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7504 (.A(net4275),
    .X(net8031));
 sky130_fd_sc_hd__clkbuf_2 hold7506 (.A(net8436),
    .X(net8033));
 sky130_fd_sc_hd__clkbuf_4 hold7507 (.A(net7816),
    .X(net8034));
 sky130_fd_sc_hd__buf_2 hold7508 (.A(_06092_),
    .X(net8035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7509 (.A(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(net8036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(net6280),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7510 (.A(net4414),
    .X(net8037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7511 (.A(net3508),
    .X(net8038));
 sky130_fd_sc_hd__buf_1 hold7512 (.A(_02357_),
    .X(net8039));
 sky130_fd_sc_hd__clkbuf_2 hold7514 (.A(_08445_),
    .X(net8041));
 sky130_fd_sc_hd__clkbuf_2 hold7515 (.A(_08446_),
    .X(net8042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7517 (.A(_08313_),
    .X(net8044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7518 (.A(_08314_),
    .X(net8045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_03439_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7520 (.A(_02562_),
    .X(net8047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7521 (.A(_02563_),
    .X(net8048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7522 (.A(_02564_),
    .X(net8049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7523 (.A(_00600_),
    .X(net8050));
 sky130_fd_sc_hd__clkbuf_4 hold7524 (.A(net4811),
    .X(net8051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7525 (.A(_00001_),
    .X(net8052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7526 (.A(net4812),
    .X(net8053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7528 (.A(_08274_),
    .X(net8055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7529 (.A(\rbzero.wall_tracer.stepDistY[-3] ),
    .X(net8056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(_00974_),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7530 (.A(net4389),
    .X(net8057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7531 (.A(net3468),
    .X(net8058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7533 (.A(_02879_),
    .X(net8060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7534 (.A(_02881_),
    .X(net8061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7535 (.A(_02885_),
    .X(net8062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7536 (.A(_00634_),
    .X(net8063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7538 (.A(net8420),
    .X(net8065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7539 (.A(\rbzero.traced_texa[9] ),
    .X(net8066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(net6290),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7540 (.A(net1028),
    .X(net8067));
 sky130_fd_sc_hd__clkbuf_4 hold7541 (.A(net8467),
    .X(net8068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7542 (.A(_00517_),
    .X(net8069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7543 (.A(net4226),
    .X(net8070));
 sky130_fd_sc_hd__buf_1 hold7544 (.A(net7999),
    .X(net8071));
 sky130_fd_sc_hd__buf_1 hold7545 (.A(_08140_),
    .X(net8072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7547 (.A(_02582_),
    .X(net8074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7548 (.A(_02585_),
    .X(net8075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7549 (.A(_02586_),
    .X(net8076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_02484_),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7550 (.A(_00602_),
    .X(net8077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7551 (.A(\rbzero.traced_texa[10] ),
    .X(net8078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7552 (.A(net850),
    .X(net8079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7553 (.A(_00520_),
    .X(net8080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7554 (.A(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(net8081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7555 (.A(net4538),
    .X(net8082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7557 (.A(_02640_),
    .X(net8084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7558 (.A(_02642_),
    .X(net8085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7559 (.A(_02646_),
    .X(net8086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_00575_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7560 (.A(_00606_),
    .X(net8087));
 sky130_fd_sc_hd__buf_2 hold7561 (.A(net4912),
    .X(net8088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7562 (.A(_00518_),
    .X(net8089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7563 (.A(net4291),
    .X(net8090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7565 (.A(_02821_),
    .X(net8092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7566 (.A(_02824_),
    .X(net8093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7567 (.A(_02825_),
    .X(net8094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7568 (.A(_00630_),
    .X(net8095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7569 (.A(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(net8096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(net5521),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7570 (.A(net652),
    .X(net8097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7571 (.A(_01651_),
    .X(net8098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7572 (.A(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(net8099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7573 (.A(net681),
    .X(net8100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7574 (.A(_01652_),
    .X(net8101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7575 (.A(\rbzero.pov.ready_buffer[13] ),
    .X(net8102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7576 (.A(net638),
    .X(net8103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7577 (.A(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(net8104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7578 (.A(net693),
    .X(net8105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7579 (.A(_01648_),
    .X(net8106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(net5523),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7581 (.A(_02606_),
    .X(net8108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7582 (.A(net1609),
    .X(net8109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7583 (.A(_00604_),
    .X(net8110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7585 (.A(_02845_),
    .X(net8112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7586 (.A(net1675),
    .X(net8113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7587 (.A(_00632_),
    .X(net8114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7588 (.A(\rbzero.spi_registers.texadd2[19] ),
    .X(net8115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7589 (.A(net4195),
    .X(net8116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(net6354),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7590 (.A(\rbzero.spi_registers.texadd2[1] ),
    .X(net8117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7591 (.A(net4198),
    .X(net8118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7592 (.A(\rbzero.traced_texa[1] ),
    .X(net8119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7593 (.A(net948),
    .X(net8120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7594 (.A(_00511_),
    .X(net8121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7595 (.A(\rbzero.traced_texa[-3] ),
    .X(net8122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7596 (.A(net896),
    .X(net8123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7597 (.A(_00507_),
    .X(net8124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7598 (.A(\rbzero.traced_texa[-7] ),
    .X(net8125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7599 (.A(net960),
    .X(net8126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net4923),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_02478_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7600 (.A(_00503_),
    .X(net8127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7601 (.A(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(net8128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7602 (.A(net1002),
    .X(net8129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7603 (.A(_00624_),
    .X(net8130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7604 (.A(\rbzero.traced_texa[-6] ),
    .X(net8131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7605 (.A(net1048),
    .X(net8132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7606 (.A(_00504_),
    .X(net8133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7607 (.A(\rbzero.spi_registers.texadd1[14] ),
    .X(net8134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7608 (.A(net4207),
    .X(net8135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7609 (.A(_00821_),
    .X(net8136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(_00572_),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7610 (.A(\rbzero.traced_texa[-5] ),
    .X(net8137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7611 (.A(net1120),
    .X(net8138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7612 (.A(_00505_),
    .X(net8139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7613 (.A(\rbzero.traced_texa[-4] ),
    .X(net8140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7614 (.A(net1106),
    .X(net8141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7615 (.A(_00506_),
    .X(net8142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7616 (.A(\rbzero.floor_leak[3] ),
    .X(net8143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7617 (.A(\rbzero.spi_registers.vshift[3] ),
    .X(net8144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7618 (.A(\rbzero.row_render.texu[1] ),
    .X(net8145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7619 (.A(\rbzero.row_render.texu[3] ),
    .X(net8146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(net6481),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7620 (.A(\rbzero.spi_registers.vshift[2] ),
    .X(net8147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7621 (.A(\rbzero.row_render.texu[0] ),
    .X(net8148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7622 (.A(_00494_),
    .X(net8149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7623 (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .X(net8150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7624 (.A(\rbzero.traced_texa[-11] ),
    .X(net8151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7625 (.A(\rbzero.map_overlay.i_othery[4] ),
    .X(net8152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7626 (.A(\rbzero.row_render.texu[2] ),
    .X(net8153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7627 (.A(_00496_),
    .X(net8154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7628 (.A(\rbzero.spi_registers.vshift[1] ),
    .X(net8155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7629 (.A(\rbzero.map_overlay.i_othery[3] ),
    .X(net8156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(_03148_),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7630 (.A(\rbzero.map_overlay.i_otherx[4] ),
    .X(net8157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7631 (.A(\rbzero.map_overlay.i_otherx[2] ),
    .X(net8158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7632 (.A(\rbzero.spi_registers.vshift[0] ),
    .X(net8159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7633 (.A(\rbzero.map_overlay.i_otherx[1] ),
    .X(net8160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7634 (.A(\rbzero.map_overlay.i_othery[1] ),
    .X(net8161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7635 (.A(\rbzero.map_overlay.i_othery[0] ),
    .X(net8162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7636 (.A(\rbzero.map_overlay.i_othery[2] ),
    .X(net8163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7637 (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .X(net8164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7638 (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .X(net8165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7639 (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .X(net8166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(net4355),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7640 (.A(\rbzero.map_overlay.i_mapdy[1] ),
    .X(net8167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7641 (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .X(net8168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7642 (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .X(net8169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7643 (.A(\rbzero.map_overlay.i_otherx[3] ),
    .X(net8170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7644 (.A(\rbzero.pov.ready_buffer[33] ),
    .X(net8171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7645 (.A(_01197_),
    .X(net8172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7646 (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .X(net8173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7647 (.A(\rbzero.spi_registers.got_new_texadd[3] ),
    .X(net8174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7648 (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .X(net8175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(net6286),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7650 (.A(_03739_),
    .X(net8177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7652 (.A(_03714_),
    .X(net8179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7653 (.A(\rbzero.traced_texa[0] ),
    .X(net8180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7654 (.A(_03933_),
    .X(net8181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7655 (.A(_01611_),
    .X(net8182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7657 (.A(_03713_),
    .X(net8184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7659 (.A(_03740_),
    .X(net8186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(net6288),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7661 (.A(_08041_),
    .X(net8188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7663 (.A(_08039_),
    .X(net8190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7664 (.A(\rbzero.traced_texa[-10] ),
    .X(net8191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7665 (.A(\rbzero.debug_overlay.playerX[-1] ),
    .X(net8192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7666 (.A(net2898),
    .X(net8193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7667 (.A(\rbzero.spi_registers.got_new_texadd[1] ),
    .X(net8194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7668 (.A(\rbzero.traced_texa[2] ),
    .X(net8195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7669 (.A(\rbzero.traced_texa[-1] ),
    .X(net8196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(_00954_),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7670 (.A(_03929_),
    .X(net8197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7671 (.A(_01610_),
    .X(net8198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7672 (.A(\rbzero.traced_texa[8] ),
    .X(net8199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7673 (.A(_03982_),
    .X(net8200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7675 (.A(_08040_),
    .X(net8202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7676 (.A(\rbzero.traced_texa[-2] ),
    .X(net8203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7678 (.A(_08042_),
    .X(net8205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7679 (.A(\rbzero.debug_overlay.playerY[-3] ),
    .X(net8206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(net6296),
    .X(net1295));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold7680 (.A(net3433),
    .X(net8207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7681 (.A(\rbzero.traced_texa[4] ),
    .X(net8208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7682 (.A(_03958_),
    .X(net8209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7683 (.A(_01615_),
    .X(net8210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7685 (.A(_03722_),
    .X(net8212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7686 (.A(net8519),
    .X(net8213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7687 (.A(net3457),
    .X(net8214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7688 (.A(\rbzero.debug_overlay.playerY[-5] ),
    .X(net8215));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold7689 (.A(net4344),
    .X(net8216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(_03437_),
    .X(net1296));
 sky130_fd_sc_hd__clkbuf_4 hold7690 (.A(net5779),
    .X(net8217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7691 (.A(_00000_),
    .X(net8218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7692 (.A(net8541),
    .X(net8219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7693 (.A(net3489),
    .X(net8220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7694 (.A(\rbzero.traced_texa[7] ),
    .X(net8221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7695 (.A(_03974_),
    .X(net8222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7696 (.A(\rbzero.traced_texa[3] ),
    .X(net8223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7697 (.A(\rbzero.debug_overlay.playerY[-2] ),
    .X(net8224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7698 (.A(net3445),
    .X(net8225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7699 (.A(\rbzero.debug_overlay.playerX[-8] ),
    .X(net8226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net4939),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_00972_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7700 (.A(net3536),
    .X(net8227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7701 (.A(\rbzero.traced_texa[6] ),
    .X(net8228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7702 (.A(_03968_),
    .X(net8229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7703 (.A(_01617_),
    .X(net8230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7704 (.A(\rbzero.traced_texa[-8] ),
    .X(net8231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7705 (.A(_03893_),
    .X(net8232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7706 (.A(\rbzero.traced_texa[5] ),
    .X(net8233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7707 (.A(\rbzero.traced_texa[-9] ),
    .X(net8234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7708 (.A(\rbzero.debug_overlay.playerY[2] ),
    .X(net8235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7709 (.A(\rbzero.debug_overlay.playerX[0] ),
    .X(net8236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(net6344),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7711 (.A(_08045_),
    .X(net8238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7713 (.A(_08046_),
    .X(net8240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7714 (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(net8241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7715 (.A(_02904_),
    .X(net8242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7716 (.A(_02910_),
    .X(net8243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7717 (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(net8244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7718 (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(net8245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7719 (.A(_02938_),
    .X(net8246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_04321_),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7720 (.A(_02939_),
    .X(net8247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7721 (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(net8248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7722 (.A(_04013_),
    .X(net8249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7723 (.A(\rbzero.debug_overlay.playerX[-9] ),
    .X(net8250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7724 (.A(net4167),
    .X(net8251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7725 (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(net8252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7726 (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(net8253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7727 (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(net8254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7728 (.A(_02523_),
    .X(net8255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(_01339_),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7730 (.A(_02666_),
    .X(net8257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7731 (.A(_02672_),
    .X(net8258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7732 (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(net8259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7733 (.A(_02700_),
    .X(net8260));
 sky130_fd_sc_hd__clkbuf_2 hold7734 (.A(net8071),
    .X(net8261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7735 (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(net8262));
 sky130_fd_sc_hd__clkbuf_2 hold7736 (.A(net8018),
    .X(net8263));
 sky130_fd_sc_hd__clkbuf_2 hold7737 (.A(net7832),
    .X(net8264));
 sky130_fd_sc_hd__clkbuf_2 hold7738 (.A(net8009),
    .X(net8265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7739 (.A(_08058_),
    .X(net8266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(net6304),
    .X(net1301));
 sky130_fd_sc_hd__clkbuf_2 hold7740 (.A(net8012),
    .X(net8267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7741 (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(net8268));
 sky130_fd_sc_hd__clkbuf_2 hold7742 (.A(net8029),
    .X(net8269));
 sky130_fd_sc_hd__clkbuf_2 hold7743 (.A(net7799),
    .X(net8270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7745 (.A(\rbzero.map_rom.a6 ),
    .X(net8272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7746 (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .X(net8273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7747 (.A(net4761),
    .X(net8274));
 sky130_fd_sc_hd__clkbuf_2 hold7748 (.A(net8088),
    .X(net8275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7749 (.A(\rbzero.spi_registers.new_texadd[0][22] ),
    .X(net8276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(_03431_),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_00966_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7769 (.A(\rbzero.row_render.size[10] ),
    .X(net8296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(net6408),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7770 (.A(net4193),
    .X(net8297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7771 (.A(net654),
    .X(net8298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7774 (.A(\rbzero.traced_texVinit[9] ),
    .X(net8301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7775 (.A(net4216),
    .X(net8302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7776 (.A(net1079),
    .X(net8303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7779 (.A(\rbzero.row_render.size[0] ),
    .X(net8306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_03818_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7780 (.A(net4245),
    .X(net8307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7781 (.A(net1361),
    .X(net8308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7782 (.A(\rbzero.row_render.size[3] ),
    .X(net8309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7783 (.A(net4302),
    .X(net8310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7784 (.A(net2910),
    .X(net8311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7785 (.A(\rbzero.row_render.size[9] ),
    .X(net8312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7786 (.A(net4340),
    .X(net8313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7787 (.A(net3388),
    .X(net8314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7788 (.A(\rbzero.texu_hot[5] ),
    .X(net8315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7789 (.A(net7751),
    .X(net8316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(_01257_),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7790 (.A(net3391),
    .X(net8317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7791 (.A(\rbzero.row_render.size[4] ),
    .X(net8318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7792 (.A(net4406),
    .X(net8319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7793 (.A(\rbzero.wall_tracer.stepDistX[9] ),
    .X(net8320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7794 (.A(net4387),
    .X(net8321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7795 (.A(net3466),
    .X(net8322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7796 (.A(\rbzero.wall_tracer.stepDistY[-7] ),
    .X(net8323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7797 (.A(net4402),
    .X(net8324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7798 (.A(net3491),
    .X(net8325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7799 (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(net8326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net4941),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(net6473),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7800 (.A(net4484),
    .X(net8327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7801 (.A(\rbzero.wall_tracer.stepDistX[1] ),
    .X(net8328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7802 (.A(net4482),
    .X(net8329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7803 (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .X(net8330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7804 (.A(net4497),
    .X(net8331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7805 (.A(\rbzero.wall_tracer.stepDistY[7] ),
    .X(net8332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7806 (.A(net4536),
    .X(net8333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7807 (.A(\rbzero.wall_tracer.stepDistY[8] ),
    .X(net8334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7808 (.A(net4523),
    .X(net8335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7809 (.A(\rbzero.wall_tracer.stepDistX[10] ),
    .X(net8336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(_03458_),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7810 (.A(net4621),
    .X(net8337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7811 (.A(\rbzero.wall_tracer.stepDistX[6] ),
    .X(net8338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7812 (.A(net4623),
    .X(net8339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7813 (.A(\rbzero.texu_hot[0] ),
    .X(net8340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7814 (.A(net4558),
    .X(net8341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7815 (.A(\rbzero.wall_tracer.stepDistY[9] ),
    .X(net8342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7816 (.A(net4607),
    .X(net8343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7817 (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .X(net8344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7818 (.A(net4666),
    .X(net8345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7819 (.A(\rbzero.texu_hot[2] ),
    .X(net8346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_00990_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7820 (.A(net4639),
    .X(net8347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7821 (.A(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(net8348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7822 (.A(net4460),
    .X(net8349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7823 (.A(\rbzero.wall_tracer.stepDistX[-7] ),
    .X(net8350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7824 (.A(net4629),
    .X(net8351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7825 (.A(\rbzero.texu_hot[4] ),
    .X(net8352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7826 (.A(net4768),
    .X(net8353));
 sky130_fd_sc_hd__buf_2 hold7827 (.A(_06676_),
    .X(net8354));
 sky130_fd_sc_hd__buf_2 hold7828 (.A(_07104_),
    .X(net8355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7829 (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .X(net8356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(net6312),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7830 (.A(net4741),
    .X(net8357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7831 (.A(\rbzero.texu_hot[3] ),
    .X(net8358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7832 (.A(net3501),
    .X(net8359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7834 (.A(_06632_),
    .X(net8361));
 sky130_fd_sc_hd__clkbuf_2 hold7835 (.A(net7763),
    .X(net8362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7837 (.A(_08134_),
    .X(net8364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7838 (.A(net4893),
    .X(net8365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7839 (.A(\rbzero.wall_tracer.stepDistY[-1] ),
    .X(net8366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_03459_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7840 (.A(net3776),
    .X(net8367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7842 (.A(_06687_),
    .X(net8369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7843 (.A(net7783),
    .X(net8370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7845 (.A(_08163_),
    .X(net8372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7846 (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .X(net8373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7847 (.A(net4372),
    .X(net8374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7848 (.A(_09885_),
    .X(net8375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(_00991_),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7850 (.A(_06016_),
    .X(net8377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7851 (.A(_08182_),
    .X(net8378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7852 (.A(\rbzero.wall_tracer.stepDistY[5] ),
    .X(net8379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7853 (.A(net4439),
    .X(net8380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7854 (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(net8381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7855 (.A(net4396),
    .X(net8382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7856 (.A(_09886_),
    .X(net8383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(net6455),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7863 (.A(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(net8390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7864 (.A(net4470),
    .X(net8391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7866 (.A(_08222_),
    .X(net8393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7867 (.A(\rbzero.wall_tracer.stepDistY[0] ),
    .X(net8394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7868 (.A(net4495),
    .X(net8395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(net6457),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7870 (.A(_08201_),
    .X(net8397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7872 (.A(_08431_),
    .X(net8399));
 sky130_fd_sc_hd__buf_1 hold7873 (.A(_08432_),
    .X(net8400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7875 (.A(_08120_),
    .X(net8402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7876 (.A(net4895),
    .X(net8403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7877 (.A(\rbzero.wall_tracer.stepDistX[5] ),
    .X(net8404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7878 (.A(net4652),
    .X(net8405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_01438_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7882 (.A(_08151_),
    .X(net8409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7883 (.A(_08152_),
    .X(net8410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7884 (.A(_08153_),
    .X(net8411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7885 (.A(_08154_),
    .X(net8412));
 sky130_fd_sc_hd__buf_1 hold7886 (.A(_08156_),
    .X(net8413));
 sky130_fd_sc_hd__clkbuf_4 hold7887 (.A(_08209_),
    .X(net8414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7888 (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(net8415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7889 (.A(net4582),
    .X(net8416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(net6412),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7891 (.A(_08249_),
    .X(net8418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7893 (.A(_08435_),
    .X(net8420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7895 (.A(_08174_),
    .X(net8422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7896 (.A(_08180_),
    .X(net8423));
 sky130_fd_sc_hd__buf_1 hold7898 (.A(_08193_),
    .X(net8425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net4951),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(net6414),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7907 (.A(_08149_),
    .X(net8434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7909 (.A(_08455_),
    .X(net8436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(_01091_),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7914 (.A(_06571_),
    .X(net8441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7915 (.A(net7807),
    .X(net8442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7916 (.A(_06553_),
    .X(net8443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7917 (.A(net7795),
    .X(net8444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7919 (.A(\rbzero.wall_tracer.stepDistX[-3] ),
    .X(net8446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(net6394),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7920 (.A(net4775),
    .X(net8447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(net6396),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7930 (.A(\rbzero.texu_hot[1] ),
    .X(net8457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_00947_),
    .X(net1321));
 sky130_fd_sc_hd__clkbuf_2 hold7940 (.A(net4907),
    .X(net8467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(net6308),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(net6310),
    .X(net1323));
 sky130_fd_sc_hd__clkbuf_2 hold7964 (.A(net5902),
    .X(net8491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(_01263_),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7970 (.A(_05999_),
    .X(net8497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7971 (.A(_08370_),
    .X(net8498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7973 (.A(_05995_),
    .X(net8500));
 sky130_fd_sc_hd__buf_1 hold7974 (.A(_08407_),
    .X(net8501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(net6346),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(net6348),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7992 (.A(\rbzero.debug_overlay.playerX[-3] ),
    .X(net8519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7993 (.A(_09451_),
    .X(net8520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net4953),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_01006_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8008 (.A(_09594_),
    .X(net8535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(net6300),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8014 (.A(\rbzero.debug_overlay.playerY[-8] ),
    .X(net8541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8015 (.A(_09092_),
    .X(net8542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(net6302),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(_00982_),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(net6400),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(net6402),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_00986_),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(net3737),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_03473_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(_01004_),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net4947),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(net6340),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(net6342),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_00992_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(net6274),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_03815_),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(_01254_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(net6190),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(net6192),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_00592_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(net6439),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net4949),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_03462_),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(_00994_),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(net6324),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(_03470_),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_01001_),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(net6441),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(net6443),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(_01321_),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(net6371),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(_03830_),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net5044),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_01268_),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(net3272),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_03555_),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(_01120_),
    .X(net1360));
 sky130_fd_sc_hd__buf_1 hold834 (.A(net8307),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(net6316),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(net6318),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(_01272_),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(net2097),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_03340_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net5046),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(net4231),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(net6373),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(net6375),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(_01256_),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(net6383),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(net6385),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_00588_),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(net6366),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(net6368),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(_00971_),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net4955),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(net6284),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(_03432_),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_00967_),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(net6338),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_02498_),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(_00586_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(net6553),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(net6555),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_01537_),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(net6175),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net4957),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(net6177),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_01277_),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(net6330),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(net6332),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_00595_),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(net3744),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_03415_),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(_00956_),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(net4027),
    .X(net1395));
 sky130_fd_sc_hd__buf_4 hold869 (.A(net4029),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net4943),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_02480_),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(_00573_),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(net6135),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(net6137),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_01274_),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(net5561),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_03391_),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(_00938_),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(net6387),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(_03445_),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net4945),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_00979_),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(net6523),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(net6525),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(_01312_),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(net6266),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(net6268),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_01278_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(net5508),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(net5510),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(net6418),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net6686),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(net6420),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(_00995_),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(net6389),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(net6391),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_00577_),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(net6334),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(net6336),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(_00574_),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(net4073),
    .X(net1425));
 sky130_fd_sc_hd__buf_4 hold899 (.A(net4075),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_03686_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_03378_),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(_00928_),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(net6410),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(_03404_),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_00945_),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(net6429),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(net6431),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(_00988_),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(net6306),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(_02494_),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net4749),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_00582_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(net5705),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(net5707),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(_01518_),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(net6377),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(_03822_),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_01261_),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(net6379),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(net6381),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(_00587_),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net4959),
    .X(net619));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold920 (.A(net7584),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(net6427),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_00591_),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(net6465),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(net6467),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(_01455_),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(net6369),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(_03471_),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_01002_),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(net6406),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net4961),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_02496_),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(_00584_),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(net6509),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(_03819_),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_01258_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(net6483),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_03472_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(_01003_),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(net6449),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(net6451),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net4963),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_01259_),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(net6314),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_03442_),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(_00976_),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(net3158),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(_03063_),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_00710_),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(net6445),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_03826_),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(_01264_),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net4965),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(net3837),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(_03414_),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_00955_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(net6018),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_03355_),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(_00911_),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(net6433),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(_03444_),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_00978_),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(net6614),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net6025),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(net6616),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(_01460_),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(net6416),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(_03469_),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_01000_),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(net6475),
    .X(net1492));
 sky130_fd_sc_hd__buf_4 hold966 (.A(_02481_),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(_03377_),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_00927_),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(net6421),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net6027),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(net6423),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(_01005_),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(net6533),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(net6535),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_01076_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(net6469),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_03829_),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(_01267_),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(net6147),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(net6149),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_01081_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_00593_),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(net6404),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_02491_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(_00580_),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(net6350),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(net6352),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_00999_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(net6362),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(net6364),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(_00581_),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net5585),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(net6825),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(net6827),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_01507_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(net6487),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(net6489),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(_01488_),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(net6206),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(net6208),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_01013_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(net6547),
    .X(net1526));
 sky130_fd_sc_hd__buf_2 input1 (.A(i_debug_map_overlay),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(i_gpout1_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(i_gpout1_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(i_gpout1_sel[2]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(i_gpout1_sel[3]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(i_gpout1_sel[4]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(i_gpout1_sel[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(i_gpout2_sel[0]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(i_gpout2_sel[1]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(i_gpout2_sel[2]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(i_gpout2_sel[3]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(i_debug_trace_overlay),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(i_gpout2_sel[4]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(i_gpout2_sel[5]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(i_gpout3_sel[0]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(i_gpout3_sel[1]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(i_gpout3_sel[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(i_gpout3_sel[3]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_gpout3_sel[4]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(i_gpout3_sel[5]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(i_gpout4_sel[0]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(i_gpout4_sel[1]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(i_debug_vec_overlay),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(i_gpout4_sel[2]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(i_gpout4_sel[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(i_gpout4_sel[4]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(i_gpout4_sel[5]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(i_gpout5_sel[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(i_gpout5_sel[1]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(i_gpout5_sel[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(i_gpout5_sel[3]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(i_gpout5_sel[4]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(i_gpout5_sel[5]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(i_gpout0_sel[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input40 (.A(i_mode[0]),
    .X(net40));
 sky130_fd_sc_hd__buf_8 input41 (.A(i_mode[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input42 (.A(i_mode[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_6 input43 (.A(i_reg_csb),
    .X(net43));
 sky130_fd_sc_hd__buf_6 input44 (.A(i_reg_mosi),
    .X(net44));
 sky130_fd_sc_hd__buf_6 input45 (.A(i_reg_outs_enb),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input46 (.A(i_reg_sclk),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(i_reset_lock_a),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_reset_lock_b),
    .X(net48));
 sky130_fd_sc_hd__buf_8 input49 (.A(i_tex_in[0]),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input5 (.A(i_gpout0_sel[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_8 input50 (.A(i_tex_in[1]),
    .X(net50));
 sky130_fd_sc_hd__buf_8 input51 (.A(i_tex_in[2]),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(i_tex_in[3]),
    .X(net52));
 sky130_fd_sc_hd__buf_6 input53 (.A(i_vec_csb),
    .X(net53));
 sky130_fd_sc_hd__buf_6 input54 (.A(i_vec_mosi),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 input55 (.A(i_vec_sclk),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(i_gpout0_sel[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(i_gpout0_sel[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(i_gpout0_sel[4]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(i_gpout0_sel[5]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_06465_),
    .X(net1608));
 sky130_fd_sc_hd__buf_6 max_cap75 (.A(_09172_),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 max_cap76 (.A(_07692_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 max_cap77 (.A(_06722_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 max_cap78 (.A(_06722_),
    .X(net78));
 sky130_fd_sc_hd__buf_6 max_cap79 (.A(_06643_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 max_cap81 (.A(_06539_),
    .X(net81));
 sky130_fd_sc_hd__buf_6 max_cap82 (.A(_06464_),
    .X(net82));
 sky130_fd_sc_hd__buf_2 max_cap85 (.A(_04851_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 max_cap86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_2 max_cap87 (.A(_04850_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 max_cap88 (.A(_04846_),
    .X(net88));
 sky130_fd_sc_hd__buf_2 max_cap89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 max_cap91 (.A(_09787_),
    .X(net91));
 sky130_fd_sc_hd__buf_4 max_cap92 (.A(_04028_),
    .X(net92));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_leaf_67_i_clk),
    .Y(net144));
 sky130_fd_sc_hd__buf_1 output56 (.A(net56),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__buf_1 output57 (.A(net57),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__buf_1 output58 (.A(net58),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__buf_1 output59 (.A(net59),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__buf_1 output60 (.A(net60),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__buf_1 output61 (.A(net61),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(o_hsync));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(o_reset));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(o_tex_csb));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(o_tex_out0));
 sky130_fd_sc_hd__buf_1 output73 (.A(net143),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(o_vsync));
 sky130_fd_sc_hd__buf_1 rebuffer1 (.A(_06536_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(_06987_),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_1 rebuffer11 (.A(_06944_),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_1 rebuffer12 (.A(_06898_),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_2 rebuffer13 (.A(_06808_),
    .X(net540));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer14 (.A(net540),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(net541),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 rebuffer16 (.A(net542),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 rebuffer17 (.A(net540),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 rebuffer18 (.A(net557),
    .X(net545));
 sky130_fd_sc_hd__buf_1 rebuffer19 (.A(_06663_),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_2 rebuffer2 (.A(_07028_),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 rebuffer20 (.A(net546),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_1 rebuffer21 (.A(_06978_),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_1 rebuffer22 (.A(_06945_),
    .X(net549));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer23 (.A(_06951_),
    .X(net1674));
 sky130_fd_sc_hd__clkbuf_1 rebuffer24 (.A(_06878_),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_1 rebuffer25 (.A(_06952_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer26 (.A(_08439_),
    .X(net553));
 sky130_fd_sc_hd__buf_1 rebuffer27 (.A(_06502_),
    .X(net554));
 sky130_fd_sc_hd__buf_1 rebuffer28 (.A(_06681_),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_1 rebuffer29 (.A(net555),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(net7786),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_1 rebuffer30 (.A(_06900_),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_1 rebuffer31 (.A(net3463),
    .X(net558));
 sky130_fd_sc_hd__buf_2 rebuffer32 (.A(_06902_),
    .X(net3463));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer33 (.A(_07091_),
    .X(net3498));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer34 (.A(_06996_),
    .X(net3503));
 sky130_fd_sc_hd__buf_1 rebuffer35 (.A(_06526_),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 rebuffer36 (.A(net562),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 rebuffer37 (.A(_07832_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer38 (.A(_08439_),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_2 rebuffer39 (.A(_06988_),
    .X(net566));
 sky130_fd_sc_hd__buf_1 rebuffer4 (.A(net7787),
    .X(net531));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer40 (.A(_06618_),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 rebuffer41 (.A(net567),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_1 rebuffer42 (.A(_06913_),
    .X(net3513));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer43 (.A(_06395_),
    .X(net570));
 sky130_fd_sc_hd__buf_6 rebuffer44 (.A(_06815_),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 rebuffer45 (.A(net571),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_1 rebuffer46 (.A(net571),
    .X(net573));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer47 (.A(_06953_),
    .X(net3523));
 sky130_fd_sc_hd__clkbuf_1 rebuffer48 (.A(_06643_),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_2 rebuffer49 (.A(_06643_),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(net7787),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_1 rebuffer50 (.A(net3523),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_2 rebuffer51 (.A(_06980_),
    .X(net578));
 sky130_fd_sc_hd__buf_1 rebuffer52 (.A(_06694_),
    .X(net579));
 sky130_fd_sc_hd__buf_1 rebuffer53 (.A(net579),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_1 rebuffer54 (.A(_06694_),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 rebuffer55 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_1 rebuffer56 (.A(_06744_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(_06960_),
    .X(net3526));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(_06734_),
    .X(net3533));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(net3533),
    .X(net3579));
 sky130_fd_sc_hd__clkbuf_1 rebuffer6 (.A(net1674),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(_06734_),
    .X(net3607));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer61 (.A(net3607),
    .X(net3634));
 sky130_fd_sc_hd__clkbuf_2 rebuffer7 (.A(_06981_),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_2 rebuffer8 (.A(_07071_),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_1 rebuffer9 (.A(_07026_),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_1 split23 (.A(_06503_),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_2 split32 (.A(_06435_),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_2 split33 (.A(_06533_),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_2 split34 (.A(_06531_),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_2 split42 (.A(_07304_),
    .X(net569));
 sky130_fd_sc_hd__buf_1 split47 (.A(_06433_),
    .X(net574));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_127 (.HI(net127));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_128 (.HI(net128));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_129 (.HI(net129));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_130 (.HI(net130));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_131 (.HI(net131));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_132 (.HI(net132));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_133 (.HI(net133));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_134 (.HI(net134));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_135 (.HI(net135));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_136 (.HI(net136));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_137 (.HI(net137));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_138 (.HI(net138));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_139 (.HI(net139));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_140 (.HI(net140));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_141 (.HI(net141));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_142 (.HI(net142));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__buf_6 wire80 (.A(_06655_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 wire83 (.A(net1608),
    .X(net83));
 sky130_fd_sc_hd__buf_2 wire84 (.A(_04851_),
    .X(net84));
 sky130_fd_sc_hd__buf_2 wire90 (.A(_09787_),
    .X(net90));
 assign o_rgb[0] = net93;
 assign o_rgb[10] = net101;
 assign o_rgb[11] = net102;
 assign o_rgb[12] = net103;
 assign o_rgb[13] = net104;
 assign o_rgb[16] = net105;
 assign o_rgb[17] = net106;
 assign o_rgb[18] = net107;
 assign o_rgb[19] = net108;
 assign o_rgb[1] = net94;
 assign o_rgb[20] = net109;
 assign o_rgb[21] = net110;
 assign o_rgb[2] = net95;
 assign o_rgb[3] = net96;
 assign o_rgb[4] = net97;
 assign o_rgb[5] = net98;
 assign o_rgb[8] = net99;
 assign o_rgb[9] = net100;
 assign ones[0] = net127;
 assign ones[10] = net137;
 assign ones[11] = net138;
 assign ones[12] = net139;
 assign ones[13] = net140;
 assign ones[14] = net141;
 assign ones[15] = net142;
 assign ones[1] = net128;
 assign ones[2] = net129;
 assign ones[3] = net130;
 assign ones[4] = net131;
 assign ones[5] = net132;
 assign ones[6] = net133;
 assign ones[7] = net134;
 assign ones[8] = net135;
 assign ones[9] = net136;
 assign zeros[0] = net111;
 assign zeros[10] = net121;
 assign zeros[11] = net122;
 assign zeros[12] = net123;
 assign zeros[13] = net124;
 assign zeros[14] = net125;
 assign zeros[15] = net126;
 assign zeros[1] = net112;
 assign zeros[2] = net113;
 assign zeros[3] = net114;
 assign zeros[4] = net115;
 assign zeros[5] = net116;
 assign zeros[6] = net117;
 assign zeros[7] = net118;
 assign zeros[8] = net119;
 assign zeros[9] = net120;
endmodule

